module bright_gauss_blur_1_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 113;
    end
  end

endmodule


module bright_gauss_blur_1_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1231 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f314
  logic [0:0] f314_wen;
  logic [31:0] f314_wdata;
  logic [0:0] f314_clk;
  logic [0:0] f314_rst;
  logic [31:0] f314_rdata;
  sr_buffer_32_1 f314(.wen(f314_wen), .wdata(f314_wdata), .clk(f314_clk), .rst(f314_rst), .rdata(f314_rdata));
  assign f314_clk = clk;
  assign f314_rst = rst;
  // Bindings to f314

  // f316
  logic [0:0] f316_wen;
  logic [31:0] f316_wdata;
  logic [0:0] f316_clk;
  logic [0:0] f316_rst;
  logic [31:0] f316_rdata;
  sr_buffer_32_1 f316(.wen(f316_wen), .wdata(f316_wdata), .clk(f316_clk), .rst(f316_rst), .rdata(f316_rdata));
  assign f316_clk = clk;
  assign f316_rst = rst;
  // Bindings to f316

  // f318
  logic [0:0] f318_wen;
  logic [31:0] f318_wdata;
  logic [0:0] f318_clk;
  logic [0:0] f318_rst;
  logic [31:0] f318_rdata;
  sr_buffer_32_1 f318(.wen(f318_wen), .wdata(f318_wdata), .clk(f318_clk), .rst(f318_rst), .rdata(f318_rdata));
  assign f318_clk = clk;
  assign f318_rst = rst;
  // Bindings to f318

  // f320
  logic [0:0] f320_wen;
  logic [31:0] f320_wdata;
  logic [0:0] f320_clk;
  logic [0:0] f320_rst;
  logic [31:0] f320_rdata;
  sr_buffer_32_1 f320(.wen(f320_wen), .wdata(f320_wdata), .clk(f320_clk), .rst(f320_rst), .rdata(f320_rdata));
  assign f320_clk = clk;
  assign f320_rst = rst;
  // Bindings to f320

  // f322
  logic [0:0] f322_wen;
  logic [31:0] f322_wdata;
  logic [0:0] f322_clk;
  logic [0:0] f322_rst;
  logic [31:0] f322_rdata;
  sr_buffer_32_1 f322(.wen(f322_wen), .wdata(f322_wdata), .clk(f322_clk), .rst(f322_rst), .rdata(f322_rdata));
  assign f322_clk = clk;
  assign f322_rst = rst;
  // Bindings to f322

  // f324
  logic [0:0] f324_wen;
  logic [31:0] f324_wdata;
  logic [0:0] f324_clk;
  logic [0:0] f324_rst;
  logic [31:0] f324_rdata;
  sr_buffer_32_1 f324(.wen(f324_wen), .wdata(f324_wdata), .clk(f324_clk), .rst(f324_rst), .rdata(f324_rdata));
  assign f324_clk = clk;
  assign f324_rst = rst;
  // Bindings to f324

  // f326
  logic [0:0] f326_wen;
  logic [31:0] f326_wdata;
  logic [0:0] f326_clk;
  logic [0:0] f326_rst;
  logic [31:0] f326_rdata;
  sr_buffer_32_1 f326(.wen(f326_wen), .wdata(f326_wdata), .clk(f326_clk), .rst(f326_rst), .rdata(f326_rdata));
  assign f326_clk = clk;
  assign f326_rst = rst;
  // Bindings to f326

  // f328
  logic [0:0] f328_wen;
  logic [31:0] f328_wdata;
  logic [0:0] f328_clk;
  logic [0:0] f328_rst;
  logic [31:0] f328_rdata;
  sr_buffer_32_1 f328(.wen(f328_wen), .wdata(f328_wdata), .clk(f328_clk), .rst(f328_rst), .rdata(f328_rdata));
  assign f328_clk = clk;
  assign f328_rst = rst;
  // Bindings to f328

  // f330
  logic [0:0] f330_wen;
  logic [31:0] f330_wdata;
  logic [0:0] f330_clk;
  logic [0:0] f330_rst;
  logic [31:0] f330_rdata;
  sr_buffer_32_1 f330(.wen(f330_wen), .wdata(f330_wdata), .clk(f330_clk), .rst(f330_rst), .rdata(f330_rdata));
  assign f330_clk = clk;
  assign f330_rst = rst;
  // Bindings to f330

  // f332
  logic [0:0] f332_wen;
  logic [31:0] f332_wdata;
  logic [0:0] f332_clk;
  logic [0:0] f332_rst;
  logic [31:0] f332_rdata;
  sr_buffer_32_1 f332(.wen(f332_wen), .wdata(f332_wdata), .clk(f332_clk), .rst(f332_rst), .rdata(f332_rdata));
  assign f332_clk = clk;
  assign f332_rst = rst;
  // Bindings to f332

  // f334
  logic [0:0] f334_wen;
  logic [31:0] f334_wdata;
  logic [0:0] f334_clk;
  logic [0:0] f334_rst;
  logic [31:0] f334_rdata;
  sr_buffer_32_1 f334(.wen(f334_wen), .wdata(f334_wdata), .clk(f334_clk), .rst(f334_rst), .rdata(f334_rdata));
  assign f334_clk = clk;
  assign f334_rst = rst;
  // Bindings to f334

  // f336
  logic [0:0] f336_wen;
  logic [31:0] f336_wdata;
  logic [0:0] f336_clk;
  logic [0:0] f336_rst;
  logic [31:0] f336_rdata;
  sr_buffer_32_1 f336(.wen(f336_wen), .wdata(f336_wdata), .clk(f336_clk), .rst(f336_rst), .rdata(f336_rdata));
  assign f336_clk = clk;
  assign f336_rst = rst;
  // Bindings to f336

  // f338
  logic [0:0] f338_wen;
  logic [31:0] f338_wdata;
  logic [0:0] f338_clk;
  logic [0:0] f338_rst;
  logic [31:0] f338_rdata;
  sr_buffer_32_1 f338(.wen(f338_wen), .wdata(f338_wdata), .clk(f338_clk), .rst(f338_rst), .rdata(f338_rdata));
  assign f338_clk = clk;
  assign f338_rst = rst;
  // Bindings to f338

  // f340
  logic [0:0] f340_wen;
  logic [31:0] f340_wdata;
  logic [0:0] f340_clk;
  logic [0:0] f340_rst;
  logic [31:0] f340_rdata;
  sr_buffer_32_1 f340(.wen(f340_wen), .wdata(f340_wdata), .clk(f340_clk), .rst(f340_rst), .rdata(f340_rdata));
  assign f340_clk = clk;
  assign f340_rst = rst;
  // Bindings to f340

  // f342
  logic [0:0] f342_wen;
  logic [31:0] f342_wdata;
  logic [0:0] f342_clk;
  logic [0:0] f342_rst;
  logic [31:0] f342_rdata;
  sr_buffer_32_1 f342(.wen(f342_wen), .wdata(f342_wdata), .clk(f342_clk), .rst(f342_rst), .rdata(f342_rdata));
  assign f342_clk = clk;
  assign f342_rst = rst;
  // Bindings to f342

  // f344
  logic [0:0] f344_wen;
  logic [31:0] f344_wdata;
  logic [0:0] f344_clk;
  logic [0:0] f344_rst;
  logic [31:0] f344_rdata;
  sr_buffer_32_1 f344(.wen(f344_wen), .wdata(f344_wdata), .clk(f344_clk), .rst(f344_rst), .rdata(f344_rdata));
  assign f344_clk = clk;
  assign f344_rst = rst;
  // Bindings to f344

  // f346
  logic [0:0] f346_wen;
  logic [31:0] f346_wdata;
  logic [0:0] f346_clk;
  logic [0:0] f346_rst;
  logic [31:0] f346_rdata;
  sr_buffer_32_1 f346(.wen(f346_wen), .wdata(f346_wdata), .clk(f346_clk), .rst(f346_rst), .rdata(f346_rdata));
  assign f346_clk = clk;
  assign f346_rst = rst;
  // Bindings to f346

  // f348
  logic [0:0] f348_wen;
  logic [31:0] f348_wdata;
  logic [0:0] f348_clk;
  logic [0:0] f348_rst;
  logic [31:0] f348_rdata;
  sr_buffer_32_1 f348(.wen(f348_wen), .wdata(f348_wdata), .clk(f348_clk), .rst(f348_rst), .rdata(f348_rdata));
  assign f348_clk = clk;
  assign f348_rst = rst;
  // Bindings to f348

  // f350
  logic [0:0] f350_wen;
  logic [31:0] f350_wdata;
  logic [0:0] f350_clk;
  logic [0:0] f350_rst;
  logic [31:0] f350_rdata;
  sr_buffer_32_1 f350(.wen(f350_wen), .wdata(f350_wdata), .clk(f350_clk), .rst(f350_rst), .rdata(f350_rdata));
  assign f350_clk = clk;
  assign f350_rst = rst;
  // Bindings to f350

  // f352
  logic [0:0] f352_wen;
  logic [31:0] f352_wdata;
  logic [0:0] f352_clk;
  logic [0:0] f352_rst;
  logic [31:0] f352_rdata;
  sr_buffer_32_1 f352(.wen(f352_wen), .wdata(f352_wdata), .clk(f352_clk), .rst(f352_rst), .rdata(f352_rdata));
  assign f352_clk = clk;
  assign f352_rst = rst;
  // Bindings to f352

  // f354
  logic [0:0] f354_wen;
  logic [31:0] f354_wdata;
  logic [0:0] f354_clk;
  logic [0:0] f354_rst;
  logic [31:0] f354_rdata;
  sr_buffer_32_1 f354(.wen(f354_wen), .wdata(f354_wdata), .clk(f354_clk), .rst(f354_rst), .rdata(f354_rdata));
  assign f354_clk = clk;
  assign f354_rst = rst;
  // Bindings to f354

  // f356
  logic [0:0] f356_wen;
  logic [31:0] f356_wdata;
  logic [0:0] f356_clk;
  logic [0:0] f356_rst;
  logic [31:0] f356_rdata;
  sr_buffer_32_1 f356(.wen(f356_wen), .wdata(f356_wdata), .clk(f356_clk), .rst(f356_rst), .rdata(f356_rdata));
  assign f356_clk = clk;
  assign f356_rst = rst;
  // Bindings to f356

  // f358
  logic [0:0] f358_wen;
  logic [31:0] f358_wdata;
  logic [0:0] f358_clk;
  logic [0:0] f358_rst;
  logic [31:0] f358_rdata;
  sr_buffer_32_1 f358(.wen(f358_wen), .wdata(f358_wdata), .clk(f358_clk), .rst(f358_rst), .rdata(f358_rdata));
  assign f358_clk = clk;
  assign f358_rst = rst;
  // Bindings to f358

  // f360
  logic [0:0] f360_wen;
  logic [31:0] f360_wdata;
  logic [0:0] f360_clk;
  logic [0:0] f360_rst;
  logic [31:0] f360_rdata;
  sr_buffer_32_1 f360(.wen(f360_wen), .wdata(f360_wdata), .clk(f360_clk), .rst(f360_rst), .rdata(f360_rdata));
  assign f360_clk = clk;
  assign f360_rst = rst;
  // Bindings to f360

  // f362
  logic [0:0] f362_wen;
  logic [31:0] f362_wdata;
  logic [0:0] f362_clk;
  logic [0:0] f362_rst;
  logic [31:0] f362_rdata;
  sr_buffer_32_1 f362(.wen(f362_wen), .wdata(f362_wdata), .clk(f362_clk), .rst(f362_rst), .rdata(f362_rdata));
  assign f362_clk = clk;
  assign f362_rst = rst;
  // Bindings to f362

  // f364
  logic [0:0] f364_wen;
  logic [31:0] f364_wdata;
  logic [0:0] f364_clk;
  logic [0:0] f364_rst;
  logic [31:0] f364_rdata;
  sr_buffer_32_1 f364(.wen(f364_wen), .wdata(f364_wdata), .clk(f364_clk), .rst(f364_rst), .rdata(f364_rdata));
  assign f364_clk = clk;
  assign f364_rst = rst;
  // Bindings to f364

  // f366
  logic [0:0] f366_wen;
  logic [31:0] f366_wdata;
  logic [0:0] f366_clk;
  logic [0:0] f366_rst;
  logic [31:0] f366_rdata;
  sr_buffer_32_1 f366(.wen(f366_wen), .wdata(f366_wdata), .clk(f366_clk), .rst(f366_rst), .rdata(f366_rdata));
  assign f366_clk = clk;
  assign f366_rst = rst;
  // Bindings to f366

  // f368
  logic [0:0] f368_wen;
  logic [31:0] f368_wdata;
  logic [0:0] f368_clk;
  logic [0:0] f368_rst;
  logic [31:0] f368_rdata;
  sr_buffer_32_1 f368(.wen(f368_wen), .wdata(f368_wdata), .clk(f368_clk), .rst(f368_rst), .rdata(f368_rdata));
  assign f368_clk = clk;
  assign f368_rst = rst;
  // Bindings to f368

  // f370
  logic [0:0] f370_wen;
  logic [31:0] f370_wdata;
  logic [0:0] f370_clk;
  logic [0:0] f370_rst;
  logic [31:0] f370_rdata;
  sr_buffer_32_1 f370(.wen(f370_wen), .wdata(f370_wdata), .clk(f370_clk), .rst(f370_rst), .rdata(f370_rdata));
  assign f370_clk = clk;
  assign f370_rst = rst;
  // Bindings to f370

  // f372
  logic [0:0] f372_wen;
  logic [31:0] f372_wdata;
  logic [0:0] f372_clk;
  logic [0:0] f372_rst;
  logic [31:0] f372_rdata;
  sr_buffer_32_1 f372(.wen(f372_wen), .wdata(f372_wdata), .clk(f372_clk), .rst(f372_rst), .rdata(f372_rdata));
  assign f372_clk = clk;
  assign f372_rst = rst;
  // Bindings to f372

  // f374
  logic [0:0] f374_wen;
  logic [31:0] f374_wdata;
  logic [0:0] f374_clk;
  logic [0:0] f374_rst;
  logic [31:0] f374_rdata;
  sr_buffer_32_1 f374(.wen(f374_wen), .wdata(f374_wdata), .clk(f374_clk), .rst(f374_rst), .rdata(f374_rdata));
  assign f374_clk = clk;
  assign f374_rst = rst;
  // Bindings to f374

  // f376
  logic [0:0] f376_wen;
  logic [31:0] f376_wdata;
  logic [0:0] f376_clk;
  logic [0:0] f376_rst;
  logic [31:0] f376_rdata;
  sr_buffer_32_1 f376(.wen(f376_wen), .wdata(f376_wdata), .clk(f376_clk), .rst(f376_rst), .rdata(f376_rdata));
  assign f376_clk = clk;
  assign f376_rst = rst;
  // Bindings to f376

  // f378
  logic [0:0] f378_wen;
  logic [31:0] f378_wdata;
  logic [0:0] f378_clk;
  logic [0:0] f378_rst;
  logic [31:0] f378_rdata;
  sr_buffer_32_1 f378(.wen(f378_wen), .wdata(f378_wdata), .clk(f378_clk), .rst(f378_rst), .rdata(f378_rdata));
  assign f378_clk = clk;
  assign f378_rst = rst;
  // Bindings to f378

  // f380
  logic [0:0] f380_wen;
  logic [31:0] f380_wdata;
  logic [0:0] f380_clk;
  logic [0:0] f380_rst;
  logic [31:0] f380_rdata;
  sr_buffer_32_1 f380(.wen(f380_wen), .wdata(f380_wdata), .clk(f380_clk), .rst(f380_rst), .rdata(f380_rdata));
  assign f380_clk = clk;
  assign f380_rst = rst;
  // Bindings to f380

  // f382
  logic [0:0] f382_wen;
  logic [31:0] f382_wdata;
  logic [0:0] f382_clk;
  logic [0:0] f382_rst;
  logic [31:0] f382_rdata;
  sr_buffer_32_1 f382(.wen(f382_wen), .wdata(f382_wdata), .clk(f382_clk), .rst(f382_rst), .rdata(f382_rdata));
  assign f382_clk = clk;
  assign f382_rst = rst;
  // Bindings to f382

  // f384
  logic [0:0] f384_wen;
  logic [31:0] f384_wdata;
  logic [0:0] f384_clk;
  logic [0:0] f384_rst;
  logic [31:0] f384_rdata;
  sr_buffer_32_1 f384(.wen(f384_wen), .wdata(f384_wdata), .clk(f384_clk), .rst(f384_rst), .rdata(f384_rdata));
  assign f384_clk = clk;
  assign f384_rst = rst;
  // Bindings to f384

  // f386
  logic [0:0] f386_wen;
  logic [31:0] f386_wdata;
  logic [0:0] f386_clk;
  logic [0:0] f386_rst;
  logic [31:0] f386_rdata;
  sr_buffer_32_1 f386(.wen(f386_wen), .wdata(f386_wdata), .clk(f386_clk), .rst(f386_rst), .rdata(f386_rdata));
  assign f386_clk = clk;
  assign f386_rst = rst;
  // Bindings to f386

  // f388
  logic [0:0] f388_wen;
  logic [31:0] f388_wdata;
  logic [0:0] f388_clk;
  logic [0:0] f388_rst;
  logic [31:0] f388_rdata;
  sr_buffer_32_1 f388(.wen(f388_wen), .wdata(f388_wdata), .clk(f388_clk), .rst(f388_rst), .rdata(f388_rdata));
  assign f388_clk = clk;
  assign f388_rst = rst;
  // Bindings to f388

  // f390
  logic [0:0] f390_wen;
  logic [31:0] f390_wdata;
  logic [0:0] f390_clk;
  logic [0:0] f390_rst;
  logic [31:0] f390_rdata;
  sr_buffer_32_1 f390(.wen(f390_wen), .wdata(f390_wdata), .clk(f390_clk), .rst(f390_rst), .rdata(f390_rdata));
  assign f390_clk = clk;
  assign f390_rst = rst;
  // Bindings to f390

  // f392
  logic [0:0] f392_wen;
  logic [31:0] f392_wdata;
  logic [0:0] f392_clk;
  logic [0:0] f392_rst;
  logic [31:0] f392_rdata;
  sr_buffer_32_1 f392(.wen(f392_wen), .wdata(f392_wdata), .clk(f392_clk), .rst(f392_rst), .rdata(f392_rdata));
  assign f392_clk = clk;
  assign f392_rst = rst;
  // Bindings to f392

  // f394
  logic [0:0] f394_wen;
  logic [31:0] f394_wdata;
  logic [0:0] f394_clk;
  logic [0:0] f394_rst;
  logic [31:0] f394_rdata;
  sr_buffer_32_1 f394(.wen(f394_wen), .wdata(f394_wdata), .clk(f394_clk), .rst(f394_rst), .rdata(f394_rdata));
  assign f394_clk = clk;
  assign f394_rst = rst;
  // Bindings to f394

  // f396
  logic [0:0] f396_wen;
  logic [31:0] f396_wdata;
  logic [0:0] f396_clk;
  logic [0:0] f396_rst;
  logic [31:0] f396_rdata;
  sr_buffer_32_1 f396(.wen(f396_wen), .wdata(f396_wdata), .clk(f396_clk), .rst(f396_rst), .rdata(f396_rdata));
  assign f396_clk = clk;
  assign f396_rst = rst;
  // Bindings to f396

  // f398
  logic [0:0] f398_wen;
  logic [31:0] f398_wdata;
  logic [0:0] f398_clk;
  logic [0:0] f398_rst;
  logic [31:0] f398_rdata;
  sr_buffer_32_1 f398(.wen(f398_wen), .wdata(f398_wdata), .clk(f398_clk), .rst(f398_rst), .rdata(f398_rdata));
  assign f398_clk = clk;
  assign f398_rst = rst;
  // Bindings to f398

  // f400
  logic [0:0] f400_wen;
  logic [31:0] f400_wdata;
  logic [0:0] f400_clk;
  logic [0:0] f400_rst;
  logic [31:0] f400_rdata;
  sr_buffer_32_1 f400(.wen(f400_wen), .wdata(f400_wdata), .clk(f400_clk), .rst(f400_rst), .rdata(f400_rdata));
  assign f400_clk = clk;
  assign f400_rst = rst;
  // Bindings to f400

  // f402
  logic [0:0] f402_wen;
  logic [31:0] f402_wdata;
  logic [0:0] f402_clk;
  logic [0:0] f402_rst;
  logic [31:0] f402_rdata;
  sr_buffer_32_1 f402(.wen(f402_wen), .wdata(f402_wdata), .clk(f402_clk), .rst(f402_rst), .rdata(f402_rdata));
  assign f402_clk = clk;
  assign f402_rst = rst;
  // Bindings to f402

  // f404
  logic [0:0] f404_wen;
  logic [31:0] f404_wdata;
  logic [0:0] f404_clk;
  logic [0:0] f404_rst;
  logic [31:0] f404_rdata;
  sr_buffer_32_1 f404(.wen(f404_wen), .wdata(f404_wdata), .clk(f404_clk), .rst(f404_rst), .rdata(f404_rdata));
  assign f404_clk = clk;
  assign f404_rst = rst;
  // Bindings to f404

  // f406
  logic [0:0] f406_wen;
  logic [31:0] f406_wdata;
  logic [0:0] f406_clk;
  logic [0:0] f406_rst;
  logic [31:0] f406_rdata;
  sr_buffer_32_1 f406(.wen(f406_wen), .wdata(f406_wdata), .clk(f406_clk), .rst(f406_rst), .rdata(f406_rdata));
  assign f406_clk = clk;
  assign f406_rst = rst;
  // Bindings to f406

  // f408
  logic [0:0] f408_wen;
  logic [31:0] f408_wdata;
  logic [0:0] f408_clk;
  logic [0:0] f408_rst;
  logic [31:0] f408_rdata;
  sr_buffer_32_1 f408(.wen(f408_wen), .wdata(f408_wdata), .clk(f408_clk), .rst(f408_rst), .rdata(f408_rdata));
  assign f408_clk = clk;
  assign f408_rst = rst;
  // Bindings to f408

  // f410
  logic [0:0] f410_wen;
  logic [31:0] f410_wdata;
  logic [0:0] f410_clk;
  logic [0:0] f410_rst;
  logic [31:0] f410_rdata;
  sr_buffer_32_1 f410(.wen(f410_wen), .wdata(f410_wdata), .clk(f410_clk), .rst(f410_rst), .rdata(f410_rdata));
  assign f410_clk = clk;
  assign f410_rst = rst;
  // Bindings to f410

  // f412
  logic [0:0] f412_wen;
  logic [31:0] f412_wdata;
  logic [0:0] f412_clk;
  logic [0:0] f412_rst;
  logic [31:0] f412_rdata;
  sr_buffer_32_1 f412(.wen(f412_wen), .wdata(f412_wdata), .clk(f412_clk), .rst(f412_rst), .rdata(f412_rdata));
  assign f412_clk = clk;
  assign f412_rst = rst;
  // Bindings to f412

  // f414
  logic [0:0] f414_wen;
  logic [31:0] f414_wdata;
  logic [0:0] f414_clk;
  logic [0:0] f414_rst;
  logic [31:0] f414_rdata;
  sr_buffer_32_1 f414(.wen(f414_wen), .wdata(f414_wdata), .clk(f414_clk), .rst(f414_rst), .rdata(f414_rdata));
  assign f414_clk = clk;
  assign f414_rst = rst;
  // Bindings to f414

  // f416
  logic [0:0] f416_wen;
  logic [31:0] f416_wdata;
  logic [0:0] f416_clk;
  logic [0:0] f416_rst;
  logic [31:0] f416_rdata;
  sr_buffer_32_1 f416(.wen(f416_wen), .wdata(f416_wdata), .clk(f416_clk), .rst(f416_rst), .rdata(f416_rdata));
  assign f416_clk = clk;
  assign f416_rst = rst;
  // Bindings to f416

  // f418
  logic [0:0] f418_wen;
  logic [31:0] f418_wdata;
  logic [0:0] f418_clk;
  logic [0:0] f418_rst;
  logic [31:0] f418_rdata;
  sr_buffer_32_1 f418(.wen(f418_wen), .wdata(f418_wdata), .clk(f418_clk), .rst(f418_rst), .rdata(f418_rdata));
  assign f418_clk = clk;
  assign f418_rst = rst;
  // Bindings to f418

  // f420
  logic [0:0] f420_wen;
  logic [31:0] f420_wdata;
  logic [0:0] f420_clk;
  logic [0:0] f420_rst;
  logic [31:0] f420_rdata;
  sr_buffer_32_1 f420(.wen(f420_wen), .wdata(f420_wdata), .clk(f420_clk), .rst(f420_rst), .rdata(f420_rdata));
  assign f420_clk = clk;
  assign f420_rst = rst;
  // Bindings to f420

  // f422
  logic [0:0] f422_wen;
  logic [31:0] f422_wdata;
  logic [0:0] f422_clk;
  logic [0:0] f422_rst;
  logic [31:0] f422_rdata;
  sr_buffer_32_1 f422(.wen(f422_wen), .wdata(f422_wdata), .clk(f422_clk), .rst(f422_rst), .rdata(f422_rdata));
  assign f422_clk = clk;
  assign f422_rst = rst;
  // Bindings to f422

  // f424
  logic [0:0] f424_wen;
  logic [31:0] f424_wdata;
  logic [0:0] f424_clk;
  logic [0:0] f424_rst;
  logic [31:0] f424_rdata;
  sr_buffer_32_1 f424(.wen(f424_wen), .wdata(f424_wdata), .clk(f424_clk), .rst(f424_rst), .rdata(f424_rdata));
  assign f424_clk = clk;
  assign f424_rst = rst;
  // Bindings to f424

  // f426
  logic [0:0] f426_wen;
  logic [31:0] f426_wdata;
  logic [0:0] f426_clk;
  logic [0:0] f426_rst;
  logic [31:0] f426_rdata;
  sr_buffer_32_1 f426(.wen(f426_wen), .wdata(f426_wdata), .clk(f426_clk), .rst(f426_rst), .rdata(f426_rdata));
  assign f426_clk = clk;
  assign f426_rst = rst;
  // Bindings to f426

  // f428
  logic [0:0] f428_wen;
  logic [31:0] f428_wdata;
  logic [0:0] f428_clk;
  logic [0:0] f428_rst;
  logic [31:0] f428_rdata;
  sr_buffer_32_1 f428(.wen(f428_wen), .wdata(f428_wdata), .clk(f428_clk), .rst(f428_rst), .rdata(f428_rdata));
  assign f428_clk = clk;
  assign f428_rst = rst;
  // Bindings to f428

  // f430
  logic [0:0] f430_wen;
  logic [31:0] f430_wdata;
  logic [0:0] f430_clk;
  logic [0:0] f430_rst;
  logic [31:0] f430_rdata;
  sr_buffer_32_1 f430(.wen(f430_wen), .wdata(f430_wdata), .clk(f430_clk), .rst(f430_rst), .rdata(f430_rdata));
  assign f430_clk = clk;
  assign f430_rst = rst;
  // Bindings to f430

  // f432
  logic [0:0] f432_wen;
  logic [31:0] f432_wdata;
  logic [0:0] f432_clk;
  logic [0:0] f432_rst;
  logic [31:0] f432_rdata;
  sr_buffer_32_1 f432(.wen(f432_wen), .wdata(f432_wdata), .clk(f432_clk), .rst(f432_rst), .rdata(f432_rdata));
  assign f432_clk = clk;
  assign f432_rst = rst;
  // Bindings to f432

  // f434
  logic [0:0] f434_wen;
  logic [31:0] f434_wdata;
  logic [0:0] f434_clk;
  logic [0:0] f434_rst;
  logic [31:0] f434_rdata;
  sr_buffer_32_1 f434(.wen(f434_wen), .wdata(f434_wdata), .clk(f434_clk), .rst(f434_rst), .rdata(f434_rdata));
  assign f434_clk = clk;
  assign f434_rst = rst;
  // Bindings to f434

  // f436
  logic [0:0] f436_wen;
  logic [31:0] f436_wdata;
  logic [0:0] f436_clk;
  logic [0:0] f436_rst;
  logic [31:0] f436_rdata;
  sr_buffer_32_1 f436(.wen(f436_wen), .wdata(f436_wdata), .clk(f436_clk), .rst(f436_rst), .rdata(f436_rdata));
  assign f436_clk = clk;
  assign f436_rst = rst;
  // Bindings to f436

  // f438
  logic [0:0] f438_wen;
  logic [31:0] f438_wdata;
  logic [0:0] f438_clk;
  logic [0:0] f438_rst;
  logic [31:0] f438_rdata;
  sr_buffer_32_1 f438(.wen(f438_wen), .wdata(f438_wdata), .clk(f438_clk), .rst(f438_rst), .rdata(f438_rdata));
  assign f438_clk = clk;
  assign f438_rst = rst;
  // Bindings to f438

  // f440
  logic [0:0] f440_wen;
  logic [31:0] f440_wdata;
  logic [0:0] f440_clk;
  logic [0:0] f440_rst;
  logic [31:0] f440_rdata;
  sr_buffer_32_1 f440(.wen(f440_wen), .wdata(f440_wdata), .clk(f440_clk), .rst(f440_rst), .rdata(f440_rdata));
  assign f440_clk = clk;
  assign f440_rst = rst;
  // Bindings to f440

  // f442
  logic [0:0] f442_wen;
  logic [31:0] f442_wdata;
  logic [0:0] f442_clk;
  logic [0:0] f442_rst;
  logic [31:0] f442_rdata;
  sr_buffer_32_1 f442(.wen(f442_wen), .wdata(f442_wdata), .clk(f442_clk), .rst(f442_rst), .rdata(f442_rdata));
  assign f442_clk = clk;
  assign f442_rst = rst;
  // Bindings to f442

  // f444
  logic [0:0] f444_wen;
  logic [31:0] f444_wdata;
  logic [0:0] f444_clk;
  logic [0:0] f444_rst;
  logic [31:0] f444_rdata;
  sr_buffer_32_1 f444(.wen(f444_wen), .wdata(f444_wdata), .clk(f444_clk), .rst(f444_rst), .rdata(f444_rdata));
  assign f444_clk = clk;
  assign f444_rst = rst;
  // Bindings to f444

  // f446
  logic [0:0] f446_wen;
  logic [31:0] f446_wdata;
  logic [0:0] f446_clk;
  logic [0:0] f446_rst;
  logic [31:0] f446_rdata;
  sr_buffer_32_1 f446(.wen(f446_wen), .wdata(f446_wdata), .clk(f446_clk), .rst(f446_rst), .rdata(f446_rdata));
  assign f446_clk = clk;
  assign f446_rst = rst;
  // Bindings to f446

  // f448
  logic [0:0] f448_wen;
  logic [31:0] f448_wdata;
  logic [0:0] f448_clk;
  logic [0:0] f448_rst;
  logic [31:0] f448_rdata;
  sr_buffer_32_1 f448(.wen(f448_wen), .wdata(f448_wdata), .clk(f448_clk), .rst(f448_rst), .rdata(f448_rdata));
  assign f448_clk = clk;
  assign f448_rst = rst;
  // Bindings to f448

  // f450
  logic [0:0] f450_wen;
  logic [31:0] f450_wdata;
  logic [0:0] f450_clk;
  logic [0:0] f450_rst;
  logic [31:0] f450_rdata;
  sr_buffer_32_1 f450(.wen(f450_wen), .wdata(f450_wdata), .clk(f450_clk), .rst(f450_rst), .rdata(f450_rdata));
  assign f450_clk = clk;
  assign f450_rst = rst;
  // Bindings to f450

  // f452
  logic [0:0] f452_wen;
  logic [31:0] f452_wdata;
  logic [0:0] f452_clk;
  logic [0:0] f452_rst;
  logic [31:0] f452_rdata;
  sr_buffer_32_1 f452(.wen(f452_wen), .wdata(f452_wdata), .clk(f452_clk), .rst(f452_rst), .rdata(f452_rdata));
  assign f452_clk = clk;
  assign f452_rst = rst;
  // Bindings to f452

  // f454
  logic [0:0] f454_wen;
  logic [31:0] f454_wdata;
  logic [0:0] f454_clk;
  logic [0:0] f454_rst;
  logic [31:0] f454_rdata;
  sr_buffer_32_1 f454(.wen(f454_wen), .wdata(f454_wdata), .clk(f454_clk), .rst(f454_rst), .rdata(f454_rdata));
  assign f454_clk = clk;
  assign f454_rst = rst;
  // Bindings to f454

  // f456
  logic [0:0] f456_wen;
  logic [31:0] f456_wdata;
  logic [0:0] f456_clk;
  logic [0:0] f456_rst;
  logic [31:0] f456_rdata;
  sr_buffer_32_1 f456(.wen(f456_wen), .wdata(f456_wdata), .clk(f456_clk), .rst(f456_rst), .rdata(f456_rdata));
  assign f456_clk = clk;
  assign f456_rst = rst;
  // Bindings to f456

  // f458
  logic [0:0] f458_wen;
  logic [31:0] f458_wdata;
  logic [0:0] f458_clk;
  logic [0:0] f458_rst;
  logic [31:0] f458_rdata;
  sr_buffer_32_1 f458(.wen(f458_wen), .wdata(f458_wdata), .clk(f458_clk), .rst(f458_rst), .rdata(f458_rdata));
  assign f458_clk = clk;
  assign f458_rst = rst;
  // Bindings to f458

  // f460
  logic [0:0] f460_wen;
  logic [31:0] f460_wdata;
  logic [0:0] f460_clk;
  logic [0:0] f460_rst;
  logic [31:0] f460_rdata;
  sr_buffer_32_1 f460(.wen(f460_wen), .wdata(f460_wdata), .clk(f460_clk), .rst(f460_rst), .rdata(f460_rdata));
  assign f460_clk = clk;
  assign f460_rst = rst;
  // Bindings to f460

  // f462
  logic [0:0] f462_wen;
  logic [31:0] f462_wdata;
  logic [0:0] f462_clk;
  logic [0:0] f462_rst;
  logic [31:0] f462_rdata;
  sr_buffer_32_1 f462(.wen(f462_wen), .wdata(f462_wdata), .clk(f462_clk), .rst(f462_rst), .rdata(f462_rdata));
  assign f462_clk = clk;
  assign f462_rst = rst;
  // Bindings to f462

  // f464
  logic [0:0] f464_wen;
  logic [31:0] f464_wdata;
  logic [0:0] f464_clk;
  logic [0:0] f464_rst;
  logic [31:0] f464_rdata;
  sr_buffer_32_1 f464(.wen(f464_wen), .wdata(f464_wdata), .clk(f464_clk), .rst(f464_rst), .rdata(f464_rdata));
  assign f464_clk = clk;
  assign f464_rst = rst;
  // Bindings to f464

  // f466
  logic [0:0] f466_wen;
  logic [31:0] f466_wdata;
  logic [0:0] f466_clk;
  logic [0:0] f466_rst;
  logic [31:0] f466_rdata;
  sr_buffer_32_1 f466(.wen(f466_wen), .wdata(f466_wdata), .clk(f466_clk), .rst(f466_rst), .rdata(f466_rdata));
  assign f466_clk = clk;
  assign f466_rst = rst;
  // Bindings to f466

  // f468
  logic [0:0] f468_wen;
  logic [31:0] f468_wdata;
  logic [0:0] f468_clk;
  logic [0:0] f468_rst;
  logic [31:0] f468_rdata;
  sr_buffer_32_1 f468(.wen(f468_wen), .wdata(f468_wdata), .clk(f468_clk), .rst(f468_rst), .rdata(f468_rdata));
  assign f468_clk = clk;
  assign f468_rst = rst;
  // Bindings to f468

  // f470
  logic [0:0] f470_wen;
  logic [31:0] f470_wdata;
  logic [0:0] f470_clk;
  logic [0:0] f470_rst;
  logic [31:0] f470_rdata;
  sr_buffer_32_1 f470(.wen(f470_wen), .wdata(f470_wdata), .clk(f470_clk), .rst(f470_rst), .rdata(f470_rdata));
  assign f470_clk = clk;
  assign f470_rst = rst;
  // Bindings to f470

  // f472
  logic [0:0] f472_wen;
  logic [31:0] f472_wdata;
  logic [0:0] f472_clk;
  logic [0:0] f472_rst;
  logic [31:0] f472_rdata;
  sr_buffer_32_1 f472(.wen(f472_wen), .wdata(f472_wdata), .clk(f472_clk), .rst(f472_rst), .rdata(f472_rdata));
  assign f472_clk = clk;
  assign f472_rst = rst;
  // Bindings to f472

  // f474
  logic [0:0] f474_wen;
  logic [31:0] f474_wdata;
  logic [0:0] f474_clk;
  logic [0:0] f474_rst;
  logic [31:0] f474_rdata;
  sr_buffer_32_1 f474(.wen(f474_wen), .wdata(f474_wdata), .clk(f474_clk), .rst(f474_rst), .rdata(f474_rdata));
  assign f474_clk = clk;
  assign f474_rst = rst;
  // Bindings to f474

  // f476
  logic [0:0] f476_wen;
  logic [31:0] f476_wdata;
  logic [0:0] f476_clk;
  logic [0:0] f476_rst;
  logic [31:0] f476_rdata;
  sr_buffer_32_1 f476(.wen(f476_wen), .wdata(f476_wdata), .clk(f476_clk), .rst(f476_rst), .rdata(f476_rdata));
  assign f476_clk = clk;
  assign f476_rst = rst;
  // Bindings to f476

  // f478
  logic [0:0] f478_wen;
  logic [31:0] f478_wdata;
  logic [0:0] f478_clk;
  logic [0:0] f478_rst;
  logic [31:0] f478_rdata;
  sr_buffer_32_1 f478(.wen(f478_wen), .wdata(f478_wdata), .clk(f478_clk), .rst(f478_rst), .rdata(f478_rdata));
  assign f478_clk = clk;
  assign f478_rst = rst;
  // Bindings to f478

  // f480
  logic [0:0] f480_wen;
  logic [31:0] f480_wdata;
  logic [0:0] f480_clk;
  logic [0:0] f480_rst;
  logic [31:0] f480_rdata;
  sr_buffer_32_1 f480(.wen(f480_wen), .wdata(f480_wdata), .clk(f480_clk), .rst(f480_rst), .rdata(f480_rdata));
  assign f480_clk = clk;
  assign f480_rst = rst;
  // Bindings to f480

  // f482
  logic [0:0] f482_wen;
  logic [31:0] f482_wdata;
  logic [0:0] f482_clk;
  logic [0:0] f482_rst;
  logic [31:0] f482_rdata;
  sr_buffer_32_1 f482(.wen(f482_wen), .wdata(f482_wdata), .clk(f482_clk), .rst(f482_rst), .rdata(f482_rdata));
  assign f482_clk = clk;
  assign f482_rst = rst;
  // Bindings to f482

  // f484
  logic [0:0] f484_wen;
  logic [31:0] f484_wdata;
  logic [0:0] f484_clk;
  logic [0:0] f484_rst;
  logic [31:0] f484_rdata;
  sr_buffer_32_1 f484(.wen(f484_wen), .wdata(f484_wdata), .clk(f484_clk), .rst(f484_rst), .rdata(f484_rdata));
  assign f484_clk = clk;
  assign f484_rst = rst;
  // Bindings to f484

  // f486
  logic [0:0] f486_wen;
  logic [31:0] f486_wdata;
  logic [0:0] f486_clk;
  logic [0:0] f486_rst;
  logic [31:0] f486_rdata;
  sr_buffer_32_1 f486(.wen(f486_wen), .wdata(f486_wdata), .clk(f486_clk), .rst(f486_rst), .rdata(f486_rdata));
  assign f486_clk = clk;
  assign f486_rst = rst;
  // Bindings to f486

  // f488
  logic [0:0] f488_wen;
  logic [31:0] f488_wdata;
  logic [0:0] f488_clk;
  logic [0:0] f488_rst;
  logic [31:0] f488_rdata;
  sr_buffer_32_1 f488(.wen(f488_wen), .wdata(f488_wdata), .clk(f488_clk), .rst(f488_rst), .rdata(f488_rdata));
  assign f488_clk = clk;
  assign f488_rst = rst;
  // Bindings to f488

  // f490
  logic [0:0] f490_wen;
  logic [31:0] f490_wdata;
  logic [0:0] f490_clk;
  logic [0:0] f490_rst;
  logic [31:0] f490_rdata;
  sr_buffer_32_1 f490(.wen(f490_wen), .wdata(f490_wdata), .clk(f490_clk), .rst(f490_rst), .rdata(f490_rdata));
  assign f490_clk = clk;
  assign f490_rst = rst;
  // Bindings to f490

  // f492
  logic [0:0] f492_wen;
  logic [31:0] f492_wdata;
  logic [0:0] f492_clk;
  logic [0:0] f492_rst;
  logic [31:0] f492_rdata;
  sr_buffer_32_1 f492(.wen(f492_wen), .wdata(f492_wdata), .clk(f492_clk), .rst(f492_rst), .rdata(f492_rdata));
  assign f492_clk = clk;
  assign f492_rst = rst;
  // Bindings to f492

  // f494
  logic [0:0] f494_wen;
  logic [31:0] f494_wdata;
  logic [0:0] f494_clk;
  logic [0:0] f494_rst;
  logic [31:0] f494_rdata;
  sr_buffer_32_1 f494(.wen(f494_wen), .wdata(f494_wdata), .clk(f494_clk), .rst(f494_rst), .rdata(f494_rdata));
  assign f494_clk = clk;
  assign f494_rst = rst;
  // Bindings to f494

  // f496
  logic [0:0] f496_wen;
  logic [31:0] f496_wdata;
  logic [0:0] f496_clk;
  logic [0:0] f496_rst;
  logic [31:0] f496_rdata;
  sr_buffer_32_1 f496(.wen(f496_wen), .wdata(f496_wdata), .clk(f496_clk), .rst(f496_rst), .rdata(f496_rdata));
  assign f496_clk = clk;
  assign f496_rst = rst;
  // Bindings to f496

  // f498
  logic [0:0] f498_wen;
  logic [31:0] f498_wdata;
  logic [0:0] f498_clk;
  logic [0:0] f498_rst;
  logic [31:0] f498_rdata;
  sr_buffer_32_1 f498(.wen(f498_wen), .wdata(f498_wdata), .clk(f498_clk), .rst(f498_rst), .rdata(f498_rdata));
  assign f498_clk = clk;
  assign f498_rst = rst;
  // Bindings to f498

  // f500
  logic [0:0] f500_wen;
  logic [31:0] f500_wdata;
  logic [0:0] f500_clk;
  logic [0:0] f500_rst;
  logic [31:0] f500_rdata;
  sr_buffer_32_1 f500(.wen(f500_wen), .wdata(f500_wdata), .clk(f500_clk), .rst(f500_rst), .rdata(f500_rdata));
  assign f500_clk = clk;
  assign f500_rst = rst;
  // Bindings to f500

  // f502
  logic [0:0] f502_wen;
  logic [31:0] f502_wdata;
  logic [0:0] f502_clk;
  logic [0:0] f502_rst;
  logic [31:0] f502_rdata;
  sr_buffer_32_1 f502(.wen(f502_wen), .wdata(f502_wdata), .clk(f502_clk), .rst(f502_rst), .rdata(f502_rdata));
  assign f502_clk = clk;
  assign f502_rst = rst;
  // Bindings to f502

  // f504
  logic [0:0] f504_wen;
  logic [31:0] f504_wdata;
  logic [0:0] f504_clk;
  logic [0:0] f504_rst;
  logic [31:0] f504_rdata;
  sr_buffer_32_1 f504(.wen(f504_wen), .wdata(f504_wdata), .clk(f504_clk), .rst(f504_rst), .rdata(f504_rdata));
  assign f504_clk = clk;
  assign f504_rst = rst;
  // Bindings to f504

  // f506
  logic [0:0] f506_wen;
  logic [31:0] f506_wdata;
  logic [0:0] f506_clk;
  logic [0:0] f506_rst;
  logic [31:0] f506_rdata;
  sr_buffer_32_1 f506(.wen(f506_wen), .wdata(f506_wdata), .clk(f506_clk), .rst(f506_rst), .rdata(f506_rdata));
  assign f506_clk = clk;
  assign f506_rst = rst;
  // Bindings to f506

  // f508
  logic [0:0] f508_wen;
  logic [31:0] f508_wdata;
  logic [0:0] f508_clk;
  logic [0:0] f508_rst;
  logic [31:0] f508_rdata;
  sr_buffer_32_1 f508(.wen(f508_wen), .wdata(f508_wdata), .clk(f508_clk), .rst(f508_rst), .rdata(f508_rdata));
  assign f508_clk = clk;
  assign f508_rst = rst;
  // Bindings to f508

  // f510
  logic [0:0] f510_wen;
  logic [31:0] f510_wdata;
  logic [0:0] f510_clk;
  logic [0:0] f510_rst;
  logic [31:0] f510_rdata;
  sr_buffer_32_1 f510(.wen(f510_wen), .wdata(f510_wdata), .clk(f510_clk), .rst(f510_rst), .rdata(f510_rdata));
  assign f510_clk = clk;
  assign f510_rst = rst;
  // Bindings to f510

  // f512
  logic [0:0] f512_wen;
  logic [31:0] f512_wdata;
  logic [0:0] f512_clk;
  logic [0:0] f512_rst;
  logic [31:0] f512_rdata;
  sr_buffer_32_1 f512(.wen(f512_wen), .wdata(f512_wdata), .clk(f512_clk), .rst(f512_rst), .rdata(f512_rdata));
  assign f512_clk = clk;
  assign f512_rst = rst;
  // Bindings to f512

  // f514
  logic [0:0] f514_wen;
  logic [31:0] f514_wdata;
  logic [0:0] f514_clk;
  logic [0:0] f514_rst;
  logic [31:0] f514_rdata;
  sr_buffer_32_1 f514(.wen(f514_wen), .wdata(f514_wdata), .clk(f514_clk), .rst(f514_rst), .rdata(f514_rdata));
  assign f514_clk = clk;
  assign f514_rst = rst;
  // Bindings to f514

  // f516
  logic [0:0] f516_wen;
  logic [31:0] f516_wdata;
  logic [0:0] f516_clk;
  logic [0:0] f516_rst;
  logic [31:0] f516_rdata;
  sr_buffer_32_1 f516(.wen(f516_wen), .wdata(f516_wdata), .clk(f516_clk), .rst(f516_rst), .rdata(f516_rdata));
  assign f516_clk = clk;
  assign f516_rst = rst;
  // Bindings to f516

  // f518
  logic [0:0] f518_wen;
  logic [31:0] f518_wdata;
  logic [0:0] f518_clk;
  logic [0:0] f518_rst;
  logic [31:0] f518_rdata;
  sr_buffer_32_1 f518(.wen(f518_wen), .wdata(f518_wdata), .clk(f518_clk), .rst(f518_rst), .rdata(f518_rdata));
  assign f518_clk = clk;
  assign f518_rst = rst;
  // Bindings to f518

  // f520
  logic [0:0] f520_wen;
  logic [31:0] f520_wdata;
  logic [0:0] f520_clk;
  logic [0:0] f520_rst;
  logic [31:0] f520_rdata;
  sr_buffer_32_1 f520(.wen(f520_wen), .wdata(f520_wdata), .clk(f520_clk), .rst(f520_rst), .rdata(f520_rdata));
  assign f520_clk = clk;
  assign f520_rst = rst;
  // Bindings to f520

  // f522
  logic [0:0] f522_wen;
  logic [31:0] f522_wdata;
  logic [0:0] f522_clk;
  logic [0:0] f522_rst;
  logic [31:0] f522_rdata;
  sr_buffer_32_1 f522(.wen(f522_wen), .wdata(f522_wdata), .clk(f522_clk), .rst(f522_rst), .rdata(f522_rdata));
  assign f522_clk = clk;
  assign f522_rst = rst;
  // Bindings to f522

  // f524
  logic [0:0] f524_wen;
  logic [31:0] f524_wdata;
  logic [0:0] f524_clk;
  logic [0:0] f524_rst;
  logic [31:0] f524_rdata;
  sr_buffer_32_1 f524(.wen(f524_wen), .wdata(f524_wdata), .clk(f524_clk), .rst(f524_rst), .rdata(f524_rdata));
  assign f524_clk = clk;
  assign f524_rst = rst;
  // Bindings to f524

  // f526
  logic [0:0] f526_wen;
  logic [31:0] f526_wdata;
  logic [0:0] f526_clk;
  logic [0:0] f526_rst;
  logic [31:0] f526_rdata;
  sr_buffer_32_1 f526(.wen(f526_wen), .wdata(f526_wdata), .clk(f526_clk), .rst(f526_rst), .rdata(f526_rdata));
  assign f526_clk = clk;
  assign f526_rst = rst;
  // Bindings to f526

  // f528
  logic [0:0] f528_wen;
  logic [31:0] f528_wdata;
  logic [0:0] f528_clk;
  logic [0:0] f528_rst;
  logic [31:0] f528_rdata;
  sr_buffer_32_1 f528(.wen(f528_wen), .wdata(f528_wdata), .clk(f528_clk), .rst(f528_rst), .rdata(f528_rdata));
  assign f528_clk = clk;
  assign f528_rst = rst;
  // Bindings to f528

  // f530
  logic [0:0] f530_wen;
  logic [31:0] f530_wdata;
  logic [0:0] f530_clk;
  logic [0:0] f530_rst;
  logic [31:0] f530_rdata;
  sr_buffer_32_1 f530(.wen(f530_wen), .wdata(f530_wdata), .clk(f530_clk), .rst(f530_rst), .rdata(f530_rdata));
  assign f530_clk = clk;
  assign f530_rst = rst;
  // Bindings to f530

  // f532
  logic [0:0] f532_wen;
  logic [31:0] f532_wdata;
  logic [0:0] f532_clk;
  logic [0:0] f532_rst;
  logic [31:0] f532_rdata;
  sr_buffer_32_1 f532(.wen(f532_wen), .wdata(f532_wdata), .clk(f532_clk), .rst(f532_rst), .rdata(f532_rdata));
  assign f532_clk = clk;
  assign f532_rst = rst;
  // Bindings to f532

  // f534
  logic [0:0] f534_wen;
  logic [31:0] f534_wdata;
  logic [0:0] f534_clk;
  logic [0:0] f534_rst;
  logic [31:0] f534_rdata;
  sr_buffer_32_1 f534(.wen(f534_wen), .wdata(f534_wdata), .clk(f534_clk), .rst(f534_rst), .rdata(f534_rdata));
  assign f534_clk = clk;
  assign f534_rst = rst;
  // Bindings to f534

  // f536
  logic [0:0] f536_wen;
  logic [31:0] f536_wdata;
  logic [0:0] f536_clk;
  logic [0:0] f536_rst;
  logic [31:0] f536_rdata;
  sr_buffer_32_1 f536(.wen(f536_wen), .wdata(f536_wdata), .clk(f536_clk), .rst(f536_rst), .rdata(f536_rdata));
  assign f536_clk = clk;
  assign f536_rst = rst;
  // Bindings to f536

  // f538
  logic [0:0] f538_wen;
  logic [31:0] f538_wdata;
  logic [0:0] f538_clk;
  logic [0:0] f538_rst;
  logic [31:0] f538_rdata;
  sr_buffer_32_1 f538(.wen(f538_wen), .wdata(f538_wdata), .clk(f538_clk), .rst(f538_rst), .rdata(f538_rdata));
  assign f538_clk = clk;
  assign f538_rst = rst;
  // Bindings to f538

  // f540
  logic [0:0] f540_wen;
  logic [31:0] f540_wdata;
  logic [0:0] f540_clk;
  logic [0:0] f540_rst;
  logic [31:0] f540_rdata;
  sr_buffer_32_1 f540(.wen(f540_wen), .wdata(f540_wdata), .clk(f540_clk), .rst(f540_rst), .rdata(f540_rdata));
  assign f540_clk = clk;
  assign f540_rst = rst;
  // Bindings to f540

  // f542
  logic [0:0] f542_wen;
  logic [31:0] f542_wdata;
  logic [0:0] f542_clk;
  logic [0:0] f542_rst;
  logic [31:0] f542_rdata;
  sr_buffer_32_1 f542(.wen(f542_wen), .wdata(f542_wdata), .clk(f542_clk), .rst(f542_rst), .rdata(f542_rdata));
  assign f542_clk = clk;
  assign f542_rst = rst;
  // Bindings to f542

  // f544
  logic [0:0] f544_wen;
  logic [31:0] f544_wdata;
  logic [0:0] f544_clk;
  logic [0:0] f544_rst;
  logic [31:0] f544_rdata;
  sr_buffer_32_1 f544(.wen(f544_wen), .wdata(f544_wdata), .clk(f544_clk), .rst(f544_rst), .rdata(f544_rdata));
  assign f544_clk = clk;
  assign f544_rst = rst;
  // Bindings to f544

  // f546
  logic [0:0] f546_wen;
  logic [31:0] f546_wdata;
  logic [0:0] f546_clk;
  logic [0:0] f546_rst;
  logic [31:0] f546_rdata;
  sr_buffer_32_1 f546(.wen(f546_wen), .wdata(f546_wdata), .clk(f546_clk), .rst(f546_rst), .rdata(f546_rdata));
  assign f546_clk = clk;
  assign f546_rst = rst;
  // Bindings to f546

  // f548
  logic [0:0] f548_wen;
  logic [31:0] f548_wdata;
  logic [0:0] f548_clk;
  logic [0:0] f548_rst;
  logic [31:0] f548_rdata;
  sr_buffer_32_1 f548(.wen(f548_wen), .wdata(f548_wdata), .clk(f548_clk), .rst(f548_rst), .rdata(f548_rdata));
  assign f548_clk = clk;
  assign f548_rst = rst;
  // Bindings to f548

  // f550
  logic [0:0] f550_wen;
  logic [31:0] f550_wdata;
  logic [0:0] f550_clk;
  logic [0:0] f550_rst;
  logic [31:0] f550_rdata;
  sr_buffer_32_1 f550(.wen(f550_wen), .wdata(f550_wdata), .clk(f550_clk), .rst(f550_rst), .rdata(f550_rdata));
  assign f550_clk = clk;
  assign f550_rst = rst;
  // Bindings to f550

  // f552
  logic [0:0] f552_wen;
  logic [31:0] f552_wdata;
  logic [0:0] f552_clk;
  logic [0:0] f552_rst;
  logic [31:0] f552_rdata;
  sr_buffer_32_1 f552(.wen(f552_wen), .wdata(f552_wdata), .clk(f552_clk), .rst(f552_rst), .rdata(f552_rdata));
  assign f552_clk = clk;
  assign f552_rst = rst;
  // Bindings to f552

  // f554
  logic [0:0] f554_wen;
  logic [31:0] f554_wdata;
  logic [0:0] f554_clk;
  logic [0:0] f554_rst;
  logic [31:0] f554_rdata;
  sr_buffer_32_1 f554(.wen(f554_wen), .wdata(f554_wdata), .clk(f554_clk), .rst(f554_rst), .rdata(f554_rdata));
  assign f554_clk = clk;
  assign f554_rst = rst;
  // Bindings to f554

  // f556
  logic [0:0] f556_wen;
  logic [31:0] f556_wdata;
  logic [0:0] f556_clk;
  logic [0:0] f556_rst;
  logic [31:0] f556_rdata;
  sr_buffer_32_1 f556(.wen(f556_wen), .wdata(f556_wdata), .clk(f556_clk), .rst(f556_rst), .rdata(f556_rdata));
  assign f556_clk = clk;
  assign f556_rst = rst;
  // Bindings to f556

  // f558
  logic [0:0] f558_wen;
  logic [31:0] f558_wdata;
  logic [0:0] f558_clk;
  logic [0:0] f558_rst;
  logic [31:0] f558_rdata;
  sr_buffer_32_1 f558(.wen(f558_wen), .wdata(f558_wdata), .clk(f558_clk), .rst(f558_rst), .rdata(f558_rdata));
  assign f558_clk = clk;
  assign f558_rst = rst;
  // Bindings to f558

  // f560
  logic [0:0] f560_wen;
  logic [31:0] f560_wdata;
  logic [0:0] f560_clk;
  logic [0:0] f560_rst;
  logic [31:0] f560_rdata;
  sr_buffer_32_1 f560(.wen(f560_wen), .wdata(f560_wdata), .clk(f560_clk), .rst(f560_rst), .rdata(f560_rdata));
  assign f560_clk = clk;
  assign f560_rst = rst;
  // Bindings to f560

  // f562
  logic [0:0] f562_wen;
  logic [31:0] f562_wdata;
  logic [0:0] f562_clk;
  logic [0:0] f562_rst;
  logic [31:0] f562_rdata;
  sr_buffer_32_1 f562(.wen(f562_wen), .wdata(f562_wdata), .clk(f562_clk), .rst(f562_rst), .rdata(f562_rdata));
  assign f562_clk = clk;
  assign f562_rst = rst;
  // Bindings to f562

  // f564
  logic [0:0] f564_wen;
  logic [31:0] f564_wdata;
  logic [0:0] f564_clk;
  logic [0:0] f564_rst;
  logic [31:0] f564_rdata;
  sr_buffer_32_1 f564(.wen(f564_wen), .wdata(f564_wdata), .clk(f564_clk), .rst(f564_rst), .rdata(f564_rdata));
  assign f564_clk = clk;
  assign f564_rst = rst;
  // Bindings to f564

  // f566
  logic [0:0] f566_wen;
  logic [31:0] f566_wdata;
  logic [0:0] f566_clk;
  logic [0:0] f566_rst;
  logic [31:0] f566_rdata;
  sr_buffer_32_1 f566(.wen(f566_wen), .wdata(f566_wdata), .clk(f566_clk), .rst(f566_rst), .rdata(f566_rdata));
  assign f566_clk = clk;
  assign f566_rst = rst;
  // Bindings to f566

  // f568
  logic [0:0] f568_wen;
  logic [31:0] f568_wdata;
  logic [0:0] f568_clk;
  logic [0:0] f568_rst;
  logic [31:0] f568_rdata;
  sr_buffer_32_1 f568(.wen(f568_wen), .wdata(f568_wdata), .clk(f568_clk), .rst(f568_rst), .rdata(f568_rdata));
  assign f568_clk = clk;
  assign f568_rst = rst;
  // Bindings to f568

  // f570
  logic [0:0] f570_wen;
  logic [31:0] f570_wdata;
  logic [0:0] f570_clk;
  logic [0:0] f570_rst;
  logic [31:0] f570_rdata;
  sr_buffer_32_1 f570(.wen(f570_wen), .wdata(f570_wdata), .clk(f570_clk), .rst(f570_rst), .rdata(f570_rdata));
  assign f570_clk = clk;
  assign f570_rst = rst;
  // Bindings to f570

  // f572
  logic [0:0] f572_wen;
  logic [31:0] f572_wdata;
  logic [0:0] f572_clk;
  logic [0:0] f572_rst;
  logic [31:0] f572_rdata;
  sr_buffer_32_1 f572(.wen(f572_wen), .wdata(f572_wdata), .clk(f572_clk), .rst(f572_rst), .rdata(f572_rdata));
  assign f572_clk = clk;
  assign f572_rst = rst;
  // Bindings to f572

  // f574
  logic [0:0] f574_wen;
  logic [31:0] f574_wdata;
  logic [0:0] f574_clk;
  logic [0:0] f574_rst;
  logic [31:0] f574_rdata;
  sr_buffer_32_1 f574(.wen(f574_wen), .wdata(f574_wdata), .clk(f574_clk), .rst(f574_rst), .rdata(f574_rdata));
  assign f574_clk = clk;
  assign f574_rst = rst;
  // Bindings to f574

  // f576
  logic [0:0] f576_wen;
  logic [31:0] f576_wdata;
  logic [0:0] f576_clk;
  logic [0:0] f576_rst;
  logic [31:0] f576_rdata;
  sr_buffer_32_1 f576(.wen(f576_wen), .wdata(f576_wdata), .clk(f576_clk), .rst(f576_rst), .rdata(f576_rdata));
  assign f576_clk = clk;
  assign f576_rst = rst;
  // Bindings to f576

  // f578
  logic [0:0] f578_wen;
  logic [31:0] f578_wdata;
  logic [0:0] f578_clk;
  logic [0:0] f578_rst;
  logic [31:0] f578_rdata;
  sr_buffer_32_1 f578(.wen(f578_wen), .wdata(f578_wdata), .clk(f578_clk), .rst(f578_rst), .rdata(f578_rdata));
  assign f578_clk = clk;
  assign f578_rst = rst;
  // Bindings to f578

  // f580
  logic [0:0] f580_wen;
  logic [31:0] f580_wdata;
  logic [0:0] f580_clk;
  logic [0:0] f580_rst;
  logic [31:0] f580_rdata;
  sr_buffer_32_1 f580(.wen(f580_wen), .wdata(f580_wdata), .clk(f580_clk), .rst(f580_rst), .rdata(f580_rdata));
  assign f580_clk = clk;
  assign f580_rst = rst;
  // Bindings to f580

  // f582
  logic [0:0] f582_wen;
  logic [31:0] f582_wdata;
  logic [0:0] f582_clk;
  logic [0:0] f582_rst;
  logic [31:0] f582_rdata;
  sr_buffer_32_1 f582(.wen(f582_wen), .wdata(f582_wdata), .clk(f582_clk), .rst(f582_rst), .rdata(f582_rdata));
  assign f582_clk = clk;
  assign f582_rst = rst;
  // Bindings to f582

  // f584
  logic [0:0] f584_wen;
  logic [31:0] f584_wdata;
  logic [0:0] f584_clk;
  logic [0:0] f584_rst;
  logic [31:0] f584_rdata;
  sr_buffer_32_1 f584(.wen(f584_wen), .wdata(f584_wdata), .clk(f584_clk), .rst(f584_rst), .rdata(f584_rdata));
  assign f584_clk = clk;
  assign f584_rst = rst;
  // Bindings to f584

  // f586
  logic [0:0] f586_wen;
  logic [31:0] f586_wdata;
  logic [0:0] f586_clk;
  logic [0:0] f586_rst;
  logic [31:0] f586_rdata;
  sr_buffer_32_1 f586(.wen(f586_wen), .wdata(f586_wdata), .clk(f586_clk), .rst(f586_rst), .rdata(f586_rdata));
  assign f586_clk = clk;
  assign f586_rst = rst;
  // Bindings to f586

  // f588
  logic [0:0] f588_wen;
  logic [31:0] f588_wdata;
  logic [0:0] f588_clk;
  logic [0:0] f588_rst;
  logic [31:0] f588_rdata;
  sr_buffer_32_1 f588(.wen(f588_wen), .wdata(f588_wdata), .clk(f588_clk), .rst(f588_rst), .rdata(f588_rdata));
  assign f588_clk = clk;
  assign f588_rst = rst;
  // Bindings to f588

  // f590
  logic [0:0] f590_wen;
  logic [31:0] f590_wdata;
  logic [0:0] f590_clk;
  logic [0:0] f590_rst;
  logic [31:0] f590_rdata;
  sr_buffer_32_1 f590(.wen(f590_wen), .wdata(f590_wdata), .clk(f590_clk), .rst(f590_rst), .rdata(f590_rdata));
  assign f590_clk = clk;
  assign f590_rst = rst;
  // Bindings to f590

  // f592
  logic [0:0] f592_wen;
  logic [31:0] f592_wdata;
  logic [0:0] f592_clk;
  logic [0:0] f592_rst;
  logic [31:0] f592_rdata;
  sr_buffer_32_1 f592(.wen(f592_wen), .wdata(f592_wdata), .clk(f592_clk), .rst(f592_rst), .rdata(f592_rdata));
  assign f592_clk = clk;
  assign f592_rst = rst;
  // Bindings to f592

  // f594
  logic [0:0] f594_wen;
  logic [31:0] f594_wdata;
  logic [0:0] f594_clk;
  logic [0:0] f594_rst;
  logic [31:0] f594_rdata;
  sr_buffer_32_1 f594(.wen(f594_wen), .wdata(f594_wdata), .clk(f594_clk), .rst(f594_rst), .rdata(f594_rdata));
  assign f594_clk = clk;
  assign f594_rst = rst;
  // Bindings to f594

  // f596
  logic [0:0] f596_wen;
  logic [31:0] f596_wdata;
  logic [0:0] f596_clk;
  logic [0:0] f596_rst;
  logic [31:0] f596_rdata;
  sr_buffer_32_1 f596(.wen(f596_wen), .wdata(f596_wdata), .clk(f596_clk), .rst(f596_rst), .rdata(f596_rdata));
  assign f596_clk = clk;
  assign f596_rst = rst;
  // Bindings to f596

  // f598
  logic [0:0] f598_wen;
  logic [31:0] f598_wdata;
  logic [0:0] f598_clk;
  logic [0:0] f598_rst;
  logic [31:0] f598_rdata;
  sr_buffer_32_1 f598(.wen(f598_wen), .wdata(f598_wdata), .clk(f598_clk), .rst(f598_rst), .rdata(f598_rdata));
  assign f598_clk = clk;
  assign f598_rst = rst;
  // Bindings to f598

  // f600
  logic [0:0] f600_wen;
  logic [31:0] f600_wdata;
  logic [0:0] f600_clk;
  logic [0:0] f600_rst;
  logic [31:0] f600_rdata;
  sr_buffer_32_1 f600(.wen(f600_wen), .wdata(f600_wdata), .clk(f600_clk), .rst(f600_rst), .rdata(f600_rdata));
  assign f600_clk = clk;
  assign f600_rst = rst;
  // Bindings to f600

  // f602
  logic [0:0] f602_wen;
  logic [31:0] f602_wdata;
  logic [0:0] f602_clk;
  logic [0:0] f602_rst;
  logic [31:0] f602_rdata;
  sr_buffer_32_1 f602(.wen(f602_wen), .wdata(f602_wdata), .clk(f602_clk), .rst(f602_rst), .rdata(f602_rdata));
  assign f602_clk = clk;
  assign f602_rst = rst;
  // Bindings to f602

  // f604
  logic [0:0] f604_wen;
  logic [31:0] f604_wdata;
  logic [0:0] f604_clk;
  logic [0:0] f604_rst;
  logic [31:0] f604_rdata;
  sr_buffer_32_1 f604(.wen(f604_wen), .wdata(f604_wdata), .clk(f604_clk), .rst(f604_rst), .rdata(f604_rdata));
  assign f604_clk = clk;
  assign f604_rst = rst;
  // Bindings to f604

  // f606
  logic [0:0] f606_wen;
  logic [31:0] f606_wdata;
  logic [0:0] f606_clk;
  logic [0:0] f606_rst;
  logic [31:0] f606_rdata;
  sr_buffer_32_1 f606(.wen(f606_wen), .wdata(f606_wdata), .clk(f606_clk), .rst(f606_rst), .rdata(f606_rdata));
  assign f606_clk = clk;
  assign f606_rst = rst;
  // Bindings to f606

  // f608
  logic [0:0] f608_wen;
  logic [31:0] f608_wdata;
  logic [0:0] f608_clk;
  logic [0:0] f608_rst;
  logic [31:0] f608_rdata;
  sr_buffer_32_1 f608(.wen(f608_wen), .wdata(f608_wdata), .clk(f608_clk), .rst(f608_rst), .rdata(f608_rdata));
  assign f608_clk = clk;
  assign f608_rst = rst;
  // Bindings to f608

  // f610
  logic [0:0] f610_wen;
  logic [31:0] f610_wdata;
  logic [0:0] f610_clk;
  logic [0:0] f610_rst;
  logic [31:0] f610_rdata;
  sr_buffer_32_1 f610(.wen(f610_wen), .wdata(f610_wdata), .clk(f610_clk), .rst(f610_rst), .rdata(f610_rdata));
  assign f610_clk = clk;
  assign f610_rst = rst;
  // Bindings to f610

  // f612
  logic [0:0] f612_wen;
  logic [31:0] f612_wdata;
  logic [0:0] f612_clk;
  logic [0:0] f612_rst;
  logic [31:0] f612_rdata;
  sr_buffer_32_1 f612(.wen(f612_wen), .wdata(f612_wdata), .clk(f612_clk), .rst(f612_rst), .rdata(f612_rdata));
  assign f612_clk = clk;
  assign f612_rst = rst;
  // Bindings to f612

  // f614
  logic [0:0] f614_wen;
  logic [31:0] f614_wdata;
  logic [0:0] f614_clk;
  logic [0:0] f614_rst;
  logic [31:0] f614_rdata;
  sr_buffer_32_1 f614(.wen(f614_wen), .wdata(f614_wdata), .clk(f614_clk), .rst(f614_rst), .rdata(f614_rdata));
  assign f614_clk = clk;
  assign f614_rst = rst;
  // Bindings to f614

  // f616
  logic [0:0] f616_wen;
  logic [31:0] f616_wdata;
  logic [0:0] f616_clk;
  logic [0:0] f616_rst;
  logic [31:0] f616_rdata;
  sr_buffer_32_1 f616(.wen(f616_wen), .wdata(f616_wdata), .clk(f616_clk), .rst(f616_rst), .rdata(f616_rdata));
  assign f616_clk = clk;
  assign f616_rst = rst;
  // Bindings to f616

  // f618
  logic [0:0] f618_wen;
  logic [31:0] f618_wdata;
  logic [0:0] f618_clk;
  logic [0:0] f618_rst;
  logic [31:0] f618_rdata;
  sr_buffer_32_1 f618(.wen(f618_wen), .wdata(f618_wdata), .clk(f618_clk), .rst(f618_rst), .rdata(f618_rdata));
  assign f618_clk = clk;
  assign f618_rst = rst;
  // Bindings to f618

  // f620
  logic [0:0] f620_wen;
  logic [31:0] f620_wdata;
  logic [0:0] f620_clk;
  logic [0:0] f620_rst;
  logic [31:0] f620_rdata;
  sr_buffer_32_1 f620(.wen(f620_wen), .wdata(f620_wdata), .clk(f620_clk), .rst(f620_rst), .rdata(f620_rdata));
  assign f620_clk = clk;
  assign f620_rst = rst;
  // Bindings to f620

  // f622
  logic [0:0] f622_wen;
  logic [31:0] f622_wdata;
  logic [0:0] f622_clk;
  logic [0:0] f622_rst;
  logic [31:0] f622_rdata;
  sr_buffer_32_1 f622(.wen(f622_wen), .wdata(f622_wdata), .clk(f622_clk), .rst(f622_rst), .rdata(f622_rdata));
  assign f622_clk = clk;
  assign f622_rst = rst;
  // Bindings to f622

  // f624
  logic [0:0] f624_wen;
  logic [31:0] f624_wdata;
  logic [0:0] f624_clk;
  logic [0:0] f624_rst;
  logic [31:0] f624_rdata;
  sr_buffer_32_1 f624(.wen(f624_wen), .wdata(f624_wdata), .clk(f624_clk), .rst(f624_rst), .rdata(f624_rdata));
  assign f624_clk = clk;
  assign f624_rst = rst;
  // Bindings to f624

  // f626
  logic [0:0] f626_wen;
  logic [31:0] f626_wdata;
  logic [0:0] f626_clk;
  logic [0:0] f626_rst;
  logic [31:0] f626_rdata;
  sr_buffer_32_1 f626(.wen(f626_wen), .wdata(f626_wdata), .clk(f626_clk), .rst(f626_rst), .rdata(f626_rdata));
  assign f626_clk = clk;
  assign f626_rst = rst;
  // Bindings to f626

  // f628
  logic [0:0] f628_wen;
  logic [31:0] f628_wdata;
  logic [0:0] f628_clk;
  logic [0:0] f628_rst;
  logic [31:0] f628_rdata;
  sr_buffer_32_1 f628(.wen(f628_wen), .wdata(f628_wdata), .clk(f628_clk), .rst(f628_rst), .rdata(f628_rdata));
  assign f628_clk = clk;
  assign f628_rst = rst;
  // Bindings to f628

  // f630
  logic [0:0] f630_wen;
  logic [31:0] f630_wdata;
  logic [0:0] f630_clk;
  logic [0:0] f630_rst;
  logic [31:0] f630_rdata;
  sr_buffer_32_1 f630(.wen(f630_wen), .wdata(f630_wdata), .clk(f630_clk), .rst(f630_rst), .rdata(f630_rdata));
  assign f630_clk = clk;
  assign f630_rst = rst;
  // Bindings to f630

  // f632
  logic [0:0] f632_wen;
  logic [31:0] f632_wdata;
  logic [0:0] f632_clk;
  logic [0:0] f632_rst;
  logic [31:0] f632_rdata;
  sr_buffer_32_1 f632(.wen(f632_wen), .wdata(f632_wdata), .clk(f632_clk), .rst(f632_rst), .rdata(f632_rdata));
  assign f632_clk = clk;
  assign f632_rst = rst;
  // Bindings to f632

  // f634
  logic [0:0] f634_wen;
  logic [31:0] f634_wdata;
  logic [0:0] f634_clk;
  logic [0:0] f634_rst;
  logic [31:0] f634_rdata;
  sr_buffer_32_1 f634(.wen(f634_wen), .wdata(f634_wdata), .clk(f634_clk), .rst(f634_rst), .rdata(f634_rdata));
  assign f634_clk = clk;
  assign f634_rst = rst;
  // Bindings to f634

  // f636
  logic [0:0] f636_wen;
  logic [31:0] f636_wdata;
  logic [0:0] f636_clk;
  logic [0:0] f636_rst;
  logic [31:0] f636_rdata;
  sr_buffer_32_1 f636(.wen(f636_wen), .wdata(f636_wdata), .clk(f636_clk), .rst(f636_rst), .rdata(f636_rdata));
  assign f636_clk = clk;
  assign f636_rst = rst;
  // Bindings to f636

  // f638
  logic [0:0] f638_wen;
  logic [31:0] f638_wdata;
  logic [0:0] f638_clk;
  logic [0:0] f638_rst;
  logic [31:0] f638_rdata;
  sr_buffer_32_1 f638(.wen(f638_wen), .wdata(f638_wdata), .clk(f638_clk), .rst(f638_rst), .rdata(f638_rdata));
  assign f638_clk = clk;
  assign f638_rst = rst;
  // Bindings to f638

  // f640
  logic [0:0] f640_wen;
  logic [31:0] f640_wdata;
  logic [0:0] f640_clk;
  logic [0:0] f640_rst;
  logic [31:0] f640_rdata;
  sr_buffer_32_1 f640(.wen(f640_wen), .wdata(f640_wdata), .clk(f640_clk), .rst(f640_rst), .rdata(f640_rdata));
  assign f640_clk = clk;
  assign f640_rst = rst;
  // Bindings to f640

  // f642
  logic [0:0] f642_wen;
  logic [31:0] f642_wdata;
  logic [0:0] f642_clk;
  logic [0:0] f642_rst;
  logic [31:0] f642_rdata;
  sr_buffer_32_1 f642(.wen(f642_wen), .wdata(f642_wdata), .clk(f642_clk), .rst(f642_rst), .rdata(f642_rdata));
  assign f642_clk = clk;
  assign f642_rst = rst;
  // Bindings to f642

  // f644
  logic [0:0] f644_wen;
  logic [31:0] f644_wdata;
  logic [0:0] f644_clk;
  logic [0:0] f644_rst;
  logic [31:0] f644_rdata;
  sr_buffer_32_1 f644(.wen(f644_wen), .wdata(f644_wdata), .clk(f644_clk), .rst(f644_rst), .rdata(f644_rdata));
  assign f644_clk = clk;
  assign f644_rst = rst;
  // Bindings to f644

  // f646
  logic [0:0] f646_wen;
  logic [31:0] f646_wdata;
  logic [0:0] f646_clk;
  logic [0:0] f646_rst;
  logic [31:0] f646_rdata;
  sr_buffer_32_1 f646(.wen(f646_wen), .wdata(f646_wdata), .clk(f646_clk), .rst(f646_rst), .rdata(f646_rdata));
  assign f646_clk = clk;
  assign f646_rst = rst;
  // Bindings to f646

  // f648
  logic [0:0] f648_wen;
  logic [31:0] f648_wdata;
  logic [0:0] f648_clk;
  logic [0:0] f648_rst;
  logic [31:0] f648_rdata;
  sr_buffer_32_1 f648(.wen(f648_wen), .wdata(f648_wdata), .clk(f648_clk), .rst(f648_rst), .rdata(f648_rdata));
  assign f648_clk = clk;
  assign f648_rst = rst;
  // Bindings to f648

  // f650
  logic [0:0] f650_wen;
  logic [31:0] f650_wdata;
  logic [0:0] f650_clk;
  logic [0:0] f650_rst;
  logic [31:0] f650_rdata;
  sr_buffer_32_1 f650(.wen(f650_wen), .wdata(f650_wdata), .clk(f650_clk), .rst(f650_rst), .rdata(f650_rdata));
  assign f650_clk = clk;
  assign f650_rst = rst;
  // Bindings to f650

  // f652
  logic [0:0] f652_wen;
  logic [31:0] f652_wdata;
  logic [0:0] f652_clk;
  logic [0:0] f652_rst;
  logic [31:0] f652_rdata;
  sr_buffer_32_1 f652(.wen(f652_wen), .wdata(f652_wdata), .clk(f652_clk), .rst(f652_rst), .rdata(f652_rdata));
  assign f652_clk = clk;
  assign f652_rst = rst;
  // Bindings to f652

  // f654
  logic [0:0] f654_wen;
  logic [31:0] f654_wdata;
  logic [0:0] f654_clk;
  logic [0:0] f654_rst;
  logic [31:0] f654_rdata;
  sr_buffer_32_1 f654(.wen(f654_wen), .wdata(f654_wdata), .clk(f654_clk), .rst(f654_rst), .rdata(f654_rdata));
  assign f654_clk = clk;
  assign f654_rst = rst;
  // Bindings to f654

  // f656
  logic [0:0] f656_wen;
  logic [31:0] f656_wdata;
  logic [0:0] f656_clk;
  logic [0:0] f656_rst;
  logic [31:0] f656_rdata;
  sr_buffer_32_1 f656(.wen(f656_wen), .wdata(f656_wdata), .clk(f656_clk), .rst(f656_rst), .rdata(f656_rdata));
  assign f656_clk = clk;
  assign f656_rst = rst;
  // Bindings to f656

  // f658
  logic [0:0] f658_wen;
  logic [31:0] f658_wdata;
  logic [0:0] f658_clk;
  logic [0:0] f658_rst;
  logic [31:0] f658_rdata;
  sr_buffer_32_1 f658(.wen(f658_wen), .wdata(f658_wdata), .clk(f658_clk), .rst(f658_rst), .rdata(f658_rdata));
  assign f658_clk = clk;
  assign f658_rst = rst;
  // Bindings to f658

  // f660
  logic [0:0] f660_wen;
  logic [31:0] f660_wdata;
  logic [0:0] f660_clk;
  logic [0:0] f660_rst;
  logic [31:0] f660_rdata;
  sr_buffer_32_1 f660(.wen(f660_wen), .wdata(f660_wdata), .clk(f660_clk), .rst(f660_rst), .rdata(f660_rdata));
  assign f660_clk = clk;
  assign f660_rst = rst;
  // Bindings to f660

  // f662
  logic [0:0] f662_wen;
  logic [31:0] f662_wdata;
  logic [0:0] f662_clk;
  logic [0:0] f662_rst;
  logic [31:0] f662_rdata;
  sr_buffer_32_1 f662(.wen(f662_wen), .wdata(f662_wdata), .clk(f662_clk), .rst(f662_rst), .rdata(f662_rdata));
  assign f662_clk = clk;
  assign f662_rst = rst;
  // Bindings to f662

  // f664
  logic [0:0] f664_wen;
  logic [31:0] f664_wdata;
  logic [0:0] f664_clk;
  logic [0:0] f664_rst;
  logic [31:0] f664_rdata;
  sr_buffer_32_1 f664(.wen(f664_wen), .wdata(f664_wdata), .clk(f664_clk), .rst(f664_rst), .rdata(f664_rdata));
  assign f664_clk = clk;
  assign f664_rst = rst;
  // Bindings to f664

  // f666
  logic [0:0] f666_wen;
  logic [31:0] f666_wdata;
  logic [0:0] f666_clk;
  logic [0:0] f666_rst;
  logic [31:0] f666_rdata;
  sr_buffer_32_1 f666(.wen(f666_wen), .wdata(f666_wdata), .clk(f666_clk), .rst(f666_rst), .rdata(f666_rdata));
  assign f666_clk = clk;
  assign f666_rst = rst;
  // Bindings to f666

  // f668
  logic [0:0] f668_wen;
  logic [31:0] f668_wdata;
  logic [0:0] f668_clk;
  logic [0:0] f668_rst;
  logic [31:0] f668_rdata;
  sr_buffer_32_1 f668(.wen(f668_wen), .wdata(f668_wdata), .clk(f668_clk), .rst(f668_rst), .rdata(f668_rdata));
  assign f668_clk = clk;
  assign f668_rst = rst;
  // Bindings to f668

  // f670
  logic [0:0] f670_wen;
  logic [31:0] f670_wdata;
  logic [0:0] f670_clk;
  logic [0:0] f670_rst;
  logic [31:0] f670_rdata;
  sr_buffer_32_1 f670(.wen(f670_wen), .wdata(f670_wdata), .clk(f670_clk), .rst(f670_rst), .rdata(f670_rdata));
  assign f670_clk = clk;
  assign f670_rst = rst;
  // Bindings to f670

  // f672
  logic [0:0] f672_wen;
  logic [31:0] f672_wdata;
  logic [0:0] f672_clk;
  logic [0:0] f672_rst;
  logic [31:0] f672_rdata;
  sr_buffer_32_1 f672(.wen(f672_wen), .wdata(f672_wdata), .clk(f672_clk), .rst(f672_rst), .rdata(f672_rdata));
  assign f672_clk = clk;
  assign f672_rst = rst;
  // Bindings to f672

  // f674
  logic [0:0] f674_wen;
  logic [31:0] f674_wdata;
  logic [0:0] f674_clk;
  logic [0:0] f674_rst;
  logic [31:0] f674_rdata;
  sr_buffer_32_1 f674(.wen(f674_wen), .wdata(f674_wdata), .clk(f674_clk), .rst(f674_rst), .rdata(f674_rdata));
  assign f674_clk = clk;
  assign f674_rst = rst;
  // Bindings to f674



endmodule


module bright_gauss_blur_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 224;
    end
  end

endmodule


module bright_gauss_blur_1_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 112;
    end
  end

endmodule


module bright_gauss_blur_1_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 223;
    end
  end

endmodule


module bright_gauss_blur_1_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module bright_gauss_blur_1_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_update_0_write_wen(output [0:0] bright_update_0_write_wen);

endmodule


module bright_weights_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module bright_gauss_blur_1_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (107 - d0 >= 0) ? (222) : (-108 + d0 == 0) ? (222) : 0;
    end
  end

endmodule


module bright_gauss_blur_1_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (107 - d0 >= 0) ? (111) : (-108 + d0 == 0) ? (111) : 0;
    end
  end

endmodule


module in_wire_bright_update_0_write_wdata(output [31:0] bright_update_0_write_wdata);

endmodule


module bright_gauss_blur_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_gauss_blur_1_update_0_write_wen, input [31:0] bright_gauss_blur_1_update_0_write_wdata, input [31:0] bright_gauss_ds_1_update_0_read_dummy, output [31:0] bright_gauss_ds_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to bright_gauss_blur_1_update_0_write_wen
    // rd_0
  assign rd_0 = bright_gauss_blur_1_update_0_write_wen;

  // selector_bright_gauss_ds_1_rd0_select
  logic [0:0] selector_bright_gauss_ds_1_rd0_select_clk;
  logic [0:0] selector_bright_gauss_ds_1_rd0_select_rst;
  logic [31:0] selector_bright_gauss_ds_1_rd0_select_d0;
  logic [31:0] selector_bright_gauss_ds_1_rd0_select_d1;
  logic [31:0] selector_bright_gauss_ds_1_rd0_select_out;
  bright_gauss_ds_1_rd0_select selector_bright_gauss_ds_1_rd0_select(.clk(selector_bright_gauss_ds_1_rd0_select_clk), .rst(selector_bright_gauss_ds_1_rd0_select_rst), .d0(selector_bright_gauss_ds_1_rd0_select_d0), .d1(selector_bright_gauss_ds_1_rd0_select_d1), .out(selector_bright_gauss_ds_1_rd0_select_out));
  assign selector_bright_gauss_ds_1_rd0_select_clk = clk;
  assign selector_bright_gauss_ds_1_rd0_select_rst = rst;
  // Bindings to selector_bright_gauss_ds_1_rd0_select

  // bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1
  logic [0:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_done;
  bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1 bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1(.clk(bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_clk), .rst(bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_rst), .start(bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_start), .done(bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_done));
  assign bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_clk = clk;
  assign bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1

  // Bindings to bright_gauss_blur_1_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_gauss_blur_1_update_0_write_wdata;

  // Bindings to bright_gauss_ds_1_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_gauss_ds_1_update_0_read_dummy;

  // Bindings to bright_gauss_ds_1_update_0_read_rdata
    // wr_3
  assign bright_gauss_ds_1_update_0_read_rdata = rd_2;



endmodule


module in_wire_bright_gauss_blur_1_update_0_read_dummy(output [287:0] bright_gauss_blur_1_update_0_read_dummy);

endmodule


module out_wire_bright_gauss_blur_1_update_0_read_rdata(input [287:0] bright_gauss_blur_1_update_0_read_rdata);

endmodule


module in_wire_bright_laplace_diff_0_update_0_read_dummy(output [31:0] bright_laplace_diff_0_update_0_read_dummy);

endmodule


module out_wire_bright_laplace_diff_0_update_0_read_rdata(input [31:0] bright_laplace_diff_0_update_0_read_rdata);

endmodule


module in_wire_bright_weights_update_0_read_dummy(output [31:0] bright_weights_update_0_read_dummy);

endmodule


module out_wire_bright_weights_update_0_read_rdata(input [31:0] bright_weights_update_0_read_rdata);

endmodule


module in_wire_bright_gauss_blur_2_update_0_write_wen(output [0:0] bright_gauss_blur_2_update_0_write_wen);

endmodule


module bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module bright_gauss_ds_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_gauss_blur_2_update_0_write_wdata(output [31:0] bright_gauss_blur_2_update_0_write_wdata);

endmodule


module in_wire_bright_gauss_ds_2_update_0_read_dummy(output [31:0] bright_gauss_ds_2_update_0_read_dummy);

endmodule


module out_wire_bright_gauss_ds_2_update_0_read_rdata(input [31:0] bright_gauss_ds_2_update_0_read_rdata);

endmodule


module bright_gauss_blur_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_gauss_blur_2_update_0_write_wen, input [31:0] bright_gauss_blur_2_update_0_write_wdata, input [31:0] bright_gauss_ds_2_update_0_read_dummy, output [31:0] bright_gauss_ds_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1
  logic [0:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_done;
  bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1 bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1(.clk(bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_clk), .rst(bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_rst), .start(bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_start), .done(bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_done));
  assign bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_clk = clk;
  assign bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1

  // Bindings to bright_gauss_blur_2_update_0_write_wen
    // rd_0
  assign rd_0 = bright_gauss_blur_2_update_0_write_wen;

  // selector_bright_gauss_ds_2_rd0_select
  logic [0:0] selector_bright_gauss_ds_2_rd0_select_clk;
  logic [0:0] selector_bright_gauss_ds_2_rd0_select_rst;
  logic [31:0] selector_bright_gauss_ds_2_rd0_select_d0;
  logic [31:0] selector_bright_gauss_ds_2_rd0_select_d1;
  logic [31:0] selector_bright_gauss_ds_2_rd0_select_out;
  bright_gauss_ds_2_rd0_select selector_bright_gauss_ds_2_rd0_select(.clk(selector_bright_gauss_ds_2_rd0_select_clk), .rst(selector_bright_gauss_ds_2_rd0_select_rst), .d0(selector_bright_gauss_ds_2_rd0_select_d0), .d1(selector_bright_gauss_ds_2_rd0_select_d1), .out(selector_bright_gauss_ds_2_rd0_select_out));
  assign selector_bright_gauss_ds_2_rd0_select_clk = clk;
  assign selector_bright_gauss_ds_2_rd0_select_rst = rst;
  // Bindings to selector_bright_gauss_ds_2_rd0_select

  // Bindings to bright_gauss_blur_2_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_gauss_blur_2_update_0_write_wdata;

  // Bindings to bright_gauss_ds_2_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_gauss_ds_2_update_0_read_dummy;

  // Bindings to bright_gauss_ds_2_update_0_read_rdata
    // wr_3
  assign bright_gauss_ds_2_update_0_read_rdata = rd_2;



endmodule


module bright_gauss_ds_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_gauss_blur_3_update_0_write_wen(output [0:0] bright_gauss_blur_3_update_0_write_wen);

endmodule


module bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_278 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_gauss_blur_3_update_0_write_wdata(output [31:0] bright_gauss_blur_3_update_0_write_wdata);

endmodule


module in_wire_bright_gauss_ds_3_update_0_read_dummy(output [31:0] bright_gauss_ds_3_update_0_read_dummy);

endmodule


module out_wire_bright_gauss_ds_3_update_0_read_rdata(input [31:0] bright_gauss_ds_3_update_0_read_rdata);

endmodule


module bright_gauss_blur_2_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 56;
    end
  end

endmodule


module bright_gauss_blur_2_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module bright_gauss_blur_2_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 57;
    end
  end

endmodule


module bright_gauss_blur_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 112;
    end
  end

endmodule


module bright_gauss_blur_2_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module bright_gauss_blur_2_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 111;
    end
  end

endmodule


module bright_gauss_blur_2_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_gauss_ds_1_update_0_write_wen(output [0:0] bright_gauss_ds_1_update_0_write_wen);

endmodule


module bright_gauss_blur_2_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (51 - d0 >= 0) ? (110) : (-52 + d0 == 0) ? (110) : 0;
    end
  end

endmodule


module bright_gauss_blur_2_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (51 - d0 >= 0) ? (55) : (-52 + d0 == 0) ? (55) : 0;
    end
  end

endmodule


module in_wire_bright_gauss_ds_1_update_0_write_wdata(output [31:0] bright_gauss_ds_1_update_0_write_wdata);

endmodule


module bright_laplace_us_0_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (d1 == 0 && -98 + d0 >= 0) ? (335) : (-98 + d1 >= 0) ? ((329 - floord(d0, 2))) : (-1 + d1 == 0) ? ((384 - floord(d0, 2))) : (d1 == 0 && 97 - d0 >= 0) ? (336) : ((-d1) % 2 == 0 && -98 + d0 >= 0 && -2 + d1 >= 0 && 96 - d1 >= 0) ? (335) : ((-1 - d1) % 2 == 0 && -3 + d1 >= 0 && 97 - d1 >= 0) ? ((384 - floord(d0, 2))) : ((-d1) % 2 == 0 && 97 - d0 >= 0 && -2 + d1 >= 0 && 96 - d1 >= 0) ? (336) : 0;
    end
  end

endmodule


module in_wire_bright_gauss_blur_2_update_0_read_dummy(output [287:0] bright_gauss_blur_2_update_0_read_dummy);

endmodule


module out_wire_bright_gauss_blur_2_update_0_read_rdata(input [287:0] bright_gauss_blur_2_update_0_read_rdata);

endmodule


module in_wire_bright_laplace_diff_1_update_0_read_dummy(output [31:0] bright_laplace_diff_1_update_0_read_dummy);

endmodule


module out_wire_bright_laplace_diff_1_update_0_read_rdata(input [31:0] bright_laplace_diff_1_update_0_read_rdata);

endmodule


module in_wire_bright_laplace_us_0_update_0_read_dummy(output [31:0] bright_laplace_us_0_update_0_read_dummy);

endmodule


module out_wire_bright_laplace_us_0_update_0_read_rdata(input [31:0] bright_laplace_us_0_update_0_read_rdata);

endmodule


module in_wire_bright_laplace_diff_0_update_0_write_wen(output [0:0] bright_laplace_diff_0_update_0_write_wen);

endmodule


module in_wire_bright_laplace_diff_0_update_0_write_wdata(output [31:0] bright_laplace_diff_0_update_0_write_wdata);

endmodule


module in_wire_fused_level_0_update_0_read_dummy(output [31:0] fused_level_0_update_0_read_dummy);

endmodule


module out_wire_fused_level_0_update_0_read_rdata(input [31:0] fused_level_0_update_0_read_rdata);

endmodule


module bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_laplace_diff_1_update_0_write_wen(output [0:0] bright_laplace_diff_1_update_0_write_wen);

endmodule


module bright_laplace_diff_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_laplace_diff_0_update_0_write_wen, input [31:0] fused_level_0_update_0_read_dummy, input [31:0] bright_laplace_diff_0_update_0_write_wdata, output [31:0] fused_level_0_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to bright_laplace_diff_0_update_0_write_wen
    // rd_0
  assign rd_0 = bright_laplace_diff_0_update_0_write_wen;

  // Bindings to fused_level_0_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_0_update_0_read_dummy;

  // Bindings to bright_laplace_diff_0_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_laplace_diff_0_update_0_write_wdata;

  // Bindings to fused_level_0_update_0_read_rdata
    // wr_3
  assign fused_level_0_update_0_read_rdata = rd_2;

  // bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1
  logic [0:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_done;
  bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1 bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1(.clk(bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_clk), .rst(bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_rst), .start(bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_start), .done(bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_done));
  assign bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_clk = clk;
  assign bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1

  // selector_fused_level_0_rd0_select
  logic [0:0] selector_fused_level_0_rd0_select_clk;
  logic [0:0] selector_fused_level_0_rd0_select_rst;
  logic [31:0] selector_fused_level_0_rd0_select_d0;
  logic [31:0] selector_fused_level_0_rd0_select_d1;
  logic [31:0] selector_fused_level_0_rd0_select_out;
  fused_level_0_rd0_select selector_fused_level_0_rd0_select(.clk(selector_fused_level_0_rd0_select_clk), .rst(selector_fused_level_0_rd0_select_rst), .d0(selector_fused_level_0_rd0_select_d0), .d1(selector_fused_level_0_rd0_select_d1), .out(selector_fused_level_0_rd0_select_out));
  assign selector_fused_level_0_rd0_select_clk = clk;
  assign selector_fused_level_0_rd0_select_rst = rst;
  // Bindings to selector_fused_level_0_rd0_select



endmodule


module in_wire_bright_laplace_diff_1_update_0_write_wdata(output [31:0] bright_laplace_diff_1_update_0_write_wdata);

endmodule


module in_wire_fused_level_1_update_0_read_dummy(output [31:0] fused_level_1_update_0_read_dummy);

endmodule


module out_wire_fused_level_1_update_0_read_rdata(input [31:0] fused_level_1_update_0_read_rdata);

endmodule


module bright_weights_normed_gauss_ds_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [287:0] bright_weights_normed_gauss_blur_2_update_0_read_dummy, input [0:0] bright_weights_normed_gauss_ds_1_update_0_write_wen, input [31:0] bright_weights_normed_gauss_ds_1_update_0_write_wdata, output [287:0] bright_weights_normed_gauss_blur_2_update_0_read_rdata, input [31:0] fused_level_1_update_0_read_dummy, output [31:0] fused_level_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9
  logic [0:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_clk;
  logic [0:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_rst;
  logic [0:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_start;
  logic [0:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_done;
  bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9 bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9(.clk(bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_clk), .rst(bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_rst), .start(bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_start), .done(bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_done));
  assign bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_clk = clk;
  assign bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_rst = rst;
  // Bindings to bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9

  // bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0
  logic [0:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_clk;
  logic [0:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_rst;
  logic [0:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_start;
  logic [0:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_done;
  bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0 bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0(.clk(bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_clk), .rst(bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_rst), .start(bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_start), .done(bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_done));
  assign bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_clk = clk;
  assign bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_rst = rst;
  // Bindings to bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0

  // Bindings to bright_weights_normed_gauss_blur_2_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_gauss_blur_2_update_0_read_dummy;

  // selector_bright_weights_normed_gauss_blur_2_rd0_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd0_select_out;
  bright_weights_normed_gauss_blur_2_rd0_select selector_bright_weights_normed_gauss_blur_2_rd0_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd0_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd0_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd0_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd0_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd0_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd0_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd0_select

  // selector_bright_weights_normed_gauss_blur_2_rd1_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd1_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd1_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd1_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd1_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd1_select_out;
  bright_weights_normed_gauss_blur_2_rd1_select selector_bright_weights_normed_gauss_blur_2_rd1_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd1_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd1_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd1_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd1_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd1_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd1_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd1_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd1_select

  // selector_bright_weights_normed_gauss_blur_2_rd2_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd2_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd2_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd2_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd2_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd2_select_out;
  bright_weights_normed_gauss_blur_2_rd2_select selector_bright_weights_normed_gauss_blur_2_rd2_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd2_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd2_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd2_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd2_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd2_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd2_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd2_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd2_select

  // selector_fused_level_1_rd0_select
  logic [0:0] selector_fused_level_1_rd0_select_clk;
  logic [0:0] selector_fused_level_1_rd0_select_rst;
  logic [31:0] selector_fused_level_1_rd0_select_d0;
  logic [31:0] selector_fused_level_1_rd0_select_d1;
  logic [31:0] selector_fused_level_1_rd0_select_out;
  fused_level_1_rd0_select selector_fused_level_1_rd0_select(.clk(selector_fused_level_1_rd0_select_clk), .rst(selector_fused_level_1_rd0_select_rst), .d0(selector_fused_level_1_rd0_select_d0), .d1(selector_fused_level_1_rd0_select_d1), .out(selector_fused_level_1_rd0_select_out));
  assign selector_fused_level_1_rd0_select_clk = clk;
  assign selector_fused_level_1_rd0_select_rst = rst;
  // Bindings to selector_fused_level_1_rd0_select

  // selector_bright_weights_normed_gauss_blur_2_rd3_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd3_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd3_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd3_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd3_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd3_select_out;
  bright_weights_normed_gauss_blur_2_rd3_select selector_bright_weights_normed_gauss_blur_2_rd3_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd3_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd3_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd3_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd3_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd3_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd3_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd3_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd3_select

  // selector_bright_weights_normed_gauss_blur_2_rd4_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd4_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd4_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd4_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd4_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd4_select_out;
  bright_weights_normed_gauss_blur_2_rd4_select selector_bright_weights_normed_gauss_blur_2_rd4_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd4_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd4_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd4_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd4_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd4_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd4_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd4_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd4_select

  // selector_bright_weights_normed_gauss_blur_2_rd6_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd6_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd6_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd6_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd6_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd6_select_out;
  bright_weights_normed_gauss_blur_2_rd6_select selector_bright_weights_normed_gauss_blur_2_rd6_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd6_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd6_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd6_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd6_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd6_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd6_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd6_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd6_select

  // selector_bright_weights_normed_gauss_blur_2_rd5_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd5_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd5_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd5_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd5_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd5_select_out;
  bright_weights_normed_gauss_blur_2_rd5_select selector_bright_weights_normed_gauss_blur_2_rd5_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd5_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd5_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd5_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd5_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd5_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd5_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd5_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd5_select

  // Bindings to bright_weights_normed_gauss_ds_1_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_normed_gauss_ds_1_update_0_write_wen;

  // selector_bright_weights_normed_gauss_blur_2_rd7_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd7_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd7_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd7_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd7_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd7_select_out;
  bright_weights_normed_gauss_blur_2_rd7_select selector_bright_weights_normed_gauss_blur_2_rd7_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd7_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd7_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd7_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd7_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd7_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd7_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd7_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd7_select

  // selector_bright_weights_normed_gauss_blur_2_rd8_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd8_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd8_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd8_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd8_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd8_select_out;
  bright_weights_normed_gauss_blur_2_rd8_select selector_bright_weights_normed_gauss_blur_2_rd8_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd8_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd8_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd8_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd8_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd8_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd8_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd8_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd8_select

  // Bindings to bright_weights_normed_gauss_ds_1_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_normed_gauss_ds_1_update_0_write_wdata;

  // Bindings to bright_weights_normed_gauss_blur_2_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_gauss_blur_2_update_0_read_rdata = rd_2;

  // Bindings to fused_level_1_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_1_update_0_read_dummy;

  // Bindings to fused_level_1_update_0_read_rdata
    // wr_5
  assign fused_level_1_update_0_read_rdata = rd_4;



endmodule


module bright_weights_normed_gauss_blur_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 56;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_3_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 29;
    end
  end

endmodule


module bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_24 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_24 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16



endmodule


module in_wire_bright_weights_normed_gauss_ds_2_update_0_write_wen(output [0:0] bright_weights_normed_gauss_ds_2_update_0_write_wen);

endmodule


module bright_weights_normed_gauss_blur_3_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (23 - d0 >= 0) ? (54) : (-24 + d0 == 0) ? (54) : 0;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_3_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_3_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 55;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_3_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 28;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_3_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_3_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_3_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (23 - d0 >= 0) ? (27) : (-24 + d0 == 0) ? (27) : 0;
    end
  end

endmodule


module in_wire_bright_weights_normed_gauss_ds_2_update_0_write_wdata(output [31:0] bright_weights_normed_gauss_ds_2_update_0_write_wdata);

endmodule


module in_wire_bright_weights_normed_gauss_blur_3_update_0_read_dummy(output [287:0] bright_weights_normed_gauss_blur_3_update_0_read_dummy);

endmodule


module out_wire_bright_weights_normed_gauss_blur_3_update_0_read_rdata(input [287:0] bright_weights_normed_gauss_blur_3_update_0_read_rdata);

endmodule


module bright_weights_normed_gauss_ds_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [287:0] bright_weights_normed_gauss_blur_3_update_0_read_dummy, input [31:0] bright_weights_normed_gauss_ds_2_update_0_write_wdata, input [0:0] bright_weights_normed_gauss_ds_2_update_0_write_wen, output [287:0] bright_weights_normed_gauss_blur_3_update_0_read_rdata, input [31:0] fused_level_2_update_0_read_dummy, output [31:0] fused_level_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10
  logic [0:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_clk;
  logic [0:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_rst;
  logic [0:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_start;
  logic [0:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_done;
  bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10 bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10(.clk(bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_clk), .rst(bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_rst), .start(bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_start), .done(bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_done));
  assign bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_clk = clk;
  assign bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10

  // Bindings to bright_weights_normed_gauss_blur_3_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_gauss_blur_3_update_0_read_dummy;

  // selector_bright_weights_normed_gauss_blur_3_rd0_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd0_select_out;
  bright_weights_normed_gauss_blur_3_rd0_select selector_bright_weights_normed_gauss_blur_3_rd0_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd0_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd0_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd0_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd0_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd0_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd0_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd0_select

  // selector_bright_weights_normed_gauss_blur_3_rd1_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd1_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd1_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd1_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd1_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd1_select_out;
  bright_weights_normed_gauss_blur_3_rd1_select selector_bright_weights_normed_gauss_blur_3_rd1_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd1_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd1_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd1_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd1_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd1_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd1_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd1_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd1_select

  // selector_bright_weights_normed_gauss_blur_3_rd2_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd2_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd2_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd2_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd2_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd2_select_out;
  bright_weights_normed_gauss_blur_3_rd2_select selector_bright_weights_normed_gauss_blur_3_rd2_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd2_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd2_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd2_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd2_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd2_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd2_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd2_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd2_select

  // selector_bright_weights_normed_gauss_blur_3_rd3_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd3_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd3_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd3_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd3_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd3_select_out;
  bright_weights_normed_gauss_blur_3_rd3_select selector_bright_weights_normed_gauss_blur_3_rd3_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd3_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd3_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd3_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd3_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd3_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd3_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd3_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd3_select

  // selector_bright_weights_normed_gauss_blur_3_rd4_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd4_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd4_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd4_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd4_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd4_select_out;
  bright_weights_normed_gauss_blur_3_rd4_select selector_bright_weights_normed_gauss_blur_3_rd4_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd4_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd4_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd4_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd4_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd4_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd4_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd4_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd4_select

  // selector_bright_weights_normed_gauss_blur_3_rd6_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd6_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd6_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd6_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd6_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd6_select_out;
  bright_weights_normed_gauss_blur_3_rd6_select selector_bright_weights_normed_gauss_blur_3_rd6_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd6_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd6_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd6_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd6_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd6_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd6_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd6_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd6_select

  // selector_bright_weights_normed_gauss_blur_3_rd5_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd5_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd5_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd5_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd5_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd5_select_out;
  bright_weights_normed_gauss_blur_3_rd5_select selector_bright_weights_normed_gauss_blur_3_rd5_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd5_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd5_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd5_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd5_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd5_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd5_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd5_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd5_select

  // selector_fused_level_2_rd0_select
  logic [0:0] selector_fused_level_2_rd0_select_clk;
  logic [0:0] selector_fused_level_2_rd0_select_rst;
  logic [31:0] selector_fused_level_2_rd0_select_d0;
  logic [31:0] selector_fused_level_2_rd0_select_d1;
  logic [31:0] selector_fused_level_2_rd0_select_out;
  fused_level_2_rd0_select selector_fused_level_2_rd0_select(.clk(selector_fused_level_2_rd0_select_clk), .rst(selector_fused_level_2_rd0_select_rst), .d0(selector_fused_level_2_rd0_select_d0), .d1(selector_fused_level_2_rd0_select_d1), .out(selector_fused_level_2_rd0_select_out));
  assign selector_fused_level_2_rd0_select_clk = clk;
  assign selector_fused_level_2_rd0_select_rst = rst;
  // Bindings to selector_fused_level_2_rd0_select

  // selector_bright_weights_normed_gauss_blur_3_rd7_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd7_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd7_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd7_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd7_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd7_select_out;
  bright_weights_normed_gauss_blur_3_rd7_select selector_bright_weights_normed_gauss_blur_3_rd7_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd7_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd7_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd7_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd7_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd7_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd7_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd7_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd7_select

  // selector_bright_weights_normed_gauss_blur_3_rd8_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd8_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd8_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd8_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd8_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd8_select_out;
  bright_weights_normed_gauss_blur_3_rd8_select selector_bright_weights_normed_gauss_blur_3_rd8_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd8_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd8_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd8_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd8_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd8_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd8_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd8_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd8_select

  // Bindings to bright_weights_normed_gauss_ds_2_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_normed_gauss_ds_2_update_0_write_wdata;

  // Bindings to bright_weights_normed_gauss_ds_2_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_normed_gauss_ds_2_update_0_write_wen;

  // Bindings to bright_weights_normed_gauss_blur_3_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_gauss_blur_3_update_0_read_rdata = rd_2;

  // Bindings to fused_level_2_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_2_update_0_read_dummy;

  // Bindings to fused_level_2_update_0_read_rdata
    // wr_5
  assign fused_level_2_update_0_read_rdata = rd_4;



endmodule


module dark_dark_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_108 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_108 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2



endmodule


module dark_gauss_blur_1_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (107 - d0 >= 0) ? (222) : (-108 + d0 == 0) ? (222) : 0;
    end
  end

endmodule


module dark_gauss_blur_1_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 113;
    end
  end

endmodule


module dark_gauss_blur_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 224;
    end
  end

endmodule


module dark_gauss_blur_1_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module dark_gauss_blur_1_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 223;
    end
  end

endmodule


module dark_gauss_blur_1_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 112;
    end
  end

endmodule


module dark_gauss_blur_1_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module in_wire_dark_update_0_write_wen(output [0:0] dark_update_0_write_wen);

endmodule


module dark_gauss_blur_1_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (107 - d0 >= 0) ? (111) : (-108 + d0 == 0) ? (111) : 0;
    end
  end

endmodule


module dark_gauss_blur_1_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module bright(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_update_0_write_wen, input [31:0] bright_weights_update_0_read_dummy, input [31:0] bright_update_0_write_wdata, input [287:0] bright_gauss_blur_1_update_0_read_dummy, output [287:0] bright_gauss_blur_1_update_0_read_rdata, input [31:0] bright_laplace_diff_0_update_0_read_dummy, output [31:0] bright_laplace_diff_0_update_0_read_rdata, output [31:0] bright_weights_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;
  logic [31:0] rd_6;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;
  reg [31:0] rd_6_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;
      rd_6_stage_1 <= rd_6;


    end

  end


  // Data processing units...
  // Bindings to bright_update_0_write_wen
    // rd_0
  assign rd_0 = bright_update_0_write_wen;

  // selector_bright_weights_rd0_select
  logic [0:0] selector_bright_weights_rd0_select_clk;
  logic [0:0] selector_bright_weights_rd0_select_rst;
  logic [31:0] selector_bright_weights_rd0_select_d0;
  logic [31:0] selector_bright_weights_rd0_select_d1;
  logic [31:0] selector_bright_weights_rd0_select_out;
  bright_weights_rd0_select selector_bright_weights_rd0_select(.clk(selector_bright_weights_rd0_select_clk), .rst(selector_bright_weights_rd0_select_rst), .d0(selector_bright_weights_rd0_select_d0), .d1(selector_bright_weights_rd0_select_d1), .out(selector_bright_weights_rd0_select_out));
  assign selector_bright_weights_rd0_select_clk = clk;
  assign selector_bright_weights_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_rd0_select

  // selector_bright_gauss_blur_1_rd1_select
  logic [0:0] selector_bright_gauss_blur_1_rd1_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd1_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd1_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd1_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd1_select_out;
  bright_gauss_blur_1_rd1_select selector_bright_gauss_blur_1_rd1_select(.clk(selector_bright_gauss_blur_1_rd1_select_clk), .rst(selector_bright_gauss_blur_1_rd1_select_rst), .d0(selector_bright_gauss_blur_1_rd1_select_d0), .d1(selector_bright_gauss_blur_1_rd1_select_d1), .out(selector_bright_gauss_blur_1_rd1_select_out));
  assign selector_bright_gauss_blur_1_rd1_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd1_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd1_select

  // bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0
  logic [0:0] bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_clk;
  logic [0:0] bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_rst;
  logic [0:0] bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_start;
  logic [0:0] bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_done;
  bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0 bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0(.clk(bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_clk), .rst(bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_rst), .start(bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_start), .done(bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_done));
  assign bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_clk = clk;
  assign bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_rst = rst;
  // Bindings to bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0

  // Bindings to bright_weights_update_0_read_dummy
    // rd_6
  assign rd_6 = bright_weights_update_0_read_dummy;

  // selector_bright_gauss_blur_1_rd0_select
  logic [0:0] selector_bright_gauss_blur_1_rd0_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd0_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd0_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd0_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd0_select_out;
  bright_gauss_blur_1_rd0_select selector_bright_gauss_blur_1_rd0_select(.clk(selector_bright_gauss_blur_1_rd0_select_clk), .rst(selector_bright_gauss_blur_1_rd0_select_rst), .d0(selector_bright_gauss_blur_1_rd0_select_d0), .d1(selector_bright_gauss_blur_1_rd0_select_d1), .out(selector_bright_gauss_blur_1_rd0_select_out));
  assign selector_bright_gauss_blur_1_rd0_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd0_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd0_select

  // selector_bright_gauss_blur_1_rd2_select
  logic [0:0] selector_bright_gauss_blur_1_rd2_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd2_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd2_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd2_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd2_select_out;
  bright_gauss_blur_1_rd2_select selector_bright_gauss_blur_1_rd2_select(.clk(selector_bright_gauss_blur_1_rd2_select_clk), .rst(selector_bright_gauss_blur_1_rd2_select_rst), .d0(selector_bright_gauss_blur_1_rd2_select_d0), .d1(selector_bright_gauss_blur_1_rd2_select_d1), .out(selector_bright_gauss_blur_1_rd2_select_out));
  assign selector_bright_gauss_blur_1_rd2_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd2_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd2_select

  // selector_bright_gauss_blur_1_rd3_select
  logic [0:0] selector_bright_gauss_blur_1_rd3_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd3_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd3_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd3_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd3_select_out;
  bright_gauss_blur_1_rd3_select selector_bright_gauss_blur_1_rd3_select(.clk(selector_bright_gauss_blur_1_rd3_select_clk), .rst(selector_bright_gauss_blur_1_rd3_select_rst), .d0(selector_bright_gauss_blur_1_rd3_select_d0), .d1(selector_bright_gauss_blur_1_rd3_select_d1), .out(selector_bright_gauss_blur_1_rd3_select_out));
  assign selector_bright_gauss_blur_1_rd3_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd3_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd3_select

  // selector_bright_gauss_blur_1_rd4_select
  logic [0:0] selector_bright_gauss_blur_1_rd4_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd4_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd4_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd4_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd4_select_out;
  bright_gauss_blur_1_rd4_select selector_bright_gauss_blur_1_rd4_select(.clk(selector_bright_gauss_blur_1_rd4_select_clk), .rst(selector_bright_gauss_blur_1_rd4_select_rst), .d0(selector_bright_gauss_blur_1_rd4_select_d0), .d1(selector_bright_gauss_blur_1_rd4_select_d1), .out(selector_bright_gauss_blur_1_rd4_select_out));
  assign selector_bright_gauss_blur_1_rd4_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd4_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd4_select

  // selector_bright_gauss_blur_1_rd5_select
  logic [0:0] selector_bright_gauss_blur_1_rd5_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd5_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd5_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd5_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd5_select_out;
  bright_gauss_blur_1_rd5_select selector_bright_gauss_blur_1_rd5_select(.clk(selector_bright_gauss_blur_1_rd5_select_clk), .rst(selector_bright_gauss_blur_1_rd5_select_rst), .d0(selector_bright_gauss_blur_1_rd5_select_d0), .d1(selector_bright_gauss_blur_1_rd5_select_d1), .out(selector_bright_gauss_blur_1_rd5_select_out));
  assign selector_bright_gauss_blur_1_rd5_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd5_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd5_select

  // selector_bright_gauss_blur_1_rd6_select
  logic [0:0] selector_bright_gauss_blur_1_rd6_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd6_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd6_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd6_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd6_select_out;
  bright_gauss_blur_1_rd6_select selector_bright_gauss_blur_1_rd6_select(.clk(selector_bright_gauss_blur_1_rd6_select_clk), .rst(selector_bright_gauss_blur_1_rd6_select_rst), .d0(selector_bright_gauss_blur_1_rd6_select_d0), .d1(selector_bright_gauss_blur_1_rd6_select_d1), .out(selector_bright_gauss_blur_1_rd6_select_out));
  assign selector_bright_gauss_blur_1_rd6_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd6_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd6_select

  // selector_bright_gauss_blur_1_rd7_select
  logic [0:0] selector_bright_gauss_blur_1_rd7_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd7_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd7_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd7_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd7_select_out;
  bright_gauss_blur_1_rd7_select selector_bright_gauss_blur_1_rd7_select(.clk(selector_bright_gauss_blur_1_rd7_select_clk), .rst(selector_bright_gauss_blur_1_rd7_select_rst), .d0(selector_bright_gauss_blur_1_rd7_select_d0), .d1(selector_bright_gauss_blur_1_rd7_select_d1), .out(selector_bright_gauss_blur_1_rd7_select_out));
  assign selector_bright_gauss_blur_1_rd7_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd7_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd7_select

  // selector_bright_gauss_blur_1_rd8_select
  logic [0:0] selector_bright_gauss_blur_1_rd8_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd8_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd8_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd8_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd8_select_out;
  bright_gauss_blur_1_rd8_select selector_bright_gauss_blur_1_rd8_select(.clk(selector_bright_gauss_blur_1_rd8_select_clk), .rst(selector_bright_gauss_blur_1_rd8_select_rst), .d0(selector_bright_gauss_blur_1_rd8_select_d0), .d1(selector_bright_gauss_blur_1_rd8_select_d1), .out(selector_bright_gauss_blur_1_rd8_select_out));
  assign selector_bright_gauss_blur_1_rd8_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd8_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd8_select

  // Bindings to bright_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_update_0_write_wdata;

  // selector_bright_laplace_diff_0_rd0_select
  logic [0:0] selector_bright_laplace_diff_0_rd0_select_clk;
  logic [0:0] selector_bright_laplace_diff_0_rd0_select_rst;
  logic [31:0] selector_bright_laplace_diff_0_rd0_select_d0;
  logic [31:0] selector_bright_laplace_diff_0_rd0_select_d1;
  logic [31:0] selector_bright_laplace_diff_0_rd0_select_out;
  bright_laplace_diff_0_rd0_select selector_bright_laplace_diff_0_rd0_select(.clk(selector_bright_laplace_diff_0_rd0_select_clk), .rst(selector_bright_laplace_diff_0_rd0_select_rst), .d0(selector_bright_laplace_diff_0_rd0_select_d0), .d1(selector_bright_laplace_diff_0_rd0_select_d1), .out(selector_bright_laplace_diff_0_rd0_select_out));
  assign selector_bright_laplace_diff_0_rd0_select_clk = clk;
  assign selector_bright_laplace_diff_0_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_diff_0_rd0_select

  // Bindings to bright_gauss_blur_1_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_gauss_blur_1_update_0_read_dummy;

  // Bindings to bright_gauss_blur_1_update_0_read_rdata
    // wr_3
  assign bright_gauss_blur_1_update_0_read_rdata = rd_2;

  // Bindings to bright_laplace_diff_0_update_0_read_dummy
    // rd_4
  assign rd_4 = bright_laplace_diff_0_update_0_read_dummy;

  // Bindings to bright_laplace_diff_0_update_0_read_rdata
    // wr_5
  assign bright_laplace_diff_0_update_0_read_rdata = rd_4;

  // Bindings to bright_weights_update_0_read_rdata
    // wr_7
  assign bright_weights_update_0_read_rdata = rd_6;

  // bright_bright_update_0_write0_merged_banks_10
  logic [0:0] bright_bright_update_0_write0_merged_banks_10_clk;
  logic [0:0] bright_bright_update_0_write0_merged_banks_10_rst;
  logic [0:0] bright_bright_update_0_write0_merged_banks_10_start;
  logic [0:0] bright_bright_update_0_write0_merged_banks_10_done;
  bright_bright_update_0_write0_merged_banks_10 bright_bright_update_0_write0_merged_banks_10(.clk(bright_bright_update_0_write0_merged_banks_10_clk), .rst(bright_bright_update_0_write0_merged_banks_10_rst), .start(bright_bright_update_0_write0_merged_banks_10_start), .done(bright_bright_update_0_write0_merged_banks_10_done));
  assign bright_bright_update_0_write0_merged_banks_10_clk = clk;
  assign bright_bright_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to bright_bright_update_0_write0_merged_banks_10



endmodule


module bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_gauss_blur_1_update_0_write_wen(output [0:0] bright_gauss_blur_1_update_0_write_wen);

endmodule


module bright_gauss_ds_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_gauss_blur_1_update_0_write_wdata(output [31:0] bright_gauss_blur_1_update_0_write_wdata);

endmodule


module in_wire_bright_gauss_ds_1_update_0_read_dummy(output [31:0] bright_gauss_ds_1_update_0_read_dummy);

endmodule


module out_wire_bright_gauss_ds_1_update_0_read_rdata(input [31:0] bright_gauss_ds_1_update_0_read_rdata);

endmodule


module bright_gauss_blur_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_gauss_blur_3_update_0_write_wen, input [31:0] bright_gauss_blur_3_update_0_write_wdata, input [31:0] bright_gauss_ds_3_update_0_read_dummy, output [31:0] bright_gauss_ds_3_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1
  logic [0:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_done;
  bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1 bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1(.clk(bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_clk), .rst(bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_rst), .start(bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_start), .done(bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_done));
  assign bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_clk = clk;
  assign bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1

  // Bindings to bright_gauss_blur_3_update_0_write_wen
    // rd_0
  assign rd_0 = bright_gauss_blur_3_update_0_write_wen;

  // Bindings to bright_gauss_blur_3_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_gauss_blur_3_update_0_write_wdata;

  // selector_bright_gauss_ds_3_rd0_select
  logic [0:0] selector_bright_gauss_ds_3_rd0_select_clk;
  logic [0:0] selector_bright_gauss_ds_3_rd0_select_rst;
  logic [31:0] selector_bright_gauss_ds_3_rd0_select_d0;
  logic [31:0] selector_bright_gauss_ds_3_rd0_select_d1;
  logic [31:0] selector_bright_gauss_ds_3_rd0_select_out;
  bright_gauss_ds_3_rd0_select selector_bright_gauss_ds_3_rd0_select(.clk(selector_bright_gauss_ds_3_rd0_select_clk), .rst(selector_bright_gauss_ds_3_rd0_select_rst), .d0(selector_bright_gauss_ds_3_rd0_select_d0), .d1(selector_bright_gauss_ds_3_rd0_select_d1), .out(selector_bright_gauss_ds_3_rd0_select_out));
  assign selector_bright_gauss_ds_3_rd0_select_clk = clk;
  assign selector_bright_gauss_ds_3_rd0_select_rst = rst;
  // Bindings to selector_bright_gauss_ds_3_rd0_select

  // Bindings to bright_gauss_ds_3_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_gauss_ds_3_update_0_read_dummy;

  // Bindings to bright_gauss_ds_3_update_0_read_rdata
    // wr_3
  assign bright_gauss_ds_3_update_0_read_rdata = rd_2;



endmodule


module sr_buffer_32_279(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 279;

  reg [31:0] data [278:0];

  reg [31:0] rdata_d;

  reg [8:0] waddr;

  wire [8:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module sr_buffer_32_52(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 52;

  reg [31:0] data [51:0];

  reg [31:0] rdata_d;

  reg [5:0] waddr;

  wire [5:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_52 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_52 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16



endmodule


module bright_gauss_ds_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [287:0] bright_gauss_blur_2_update_0_read_dummy, input [0:0] bright_gauss_ds_1_update_0_write_wen, input [31:0] bright_gauss_ds_1_update_0_write_wdata, output [287:0] bright_gauss_blur_2_update_0_read_rdata, input [31:0] bright_laplace_diff_1_update_0_read_dummy, output [31:0] bright_laplace_diff_1_update_0_read_rdata, input [31:0] bright_laplace_us_0_update_0_read_dummy, output [31:0] bright_laplace_us_0_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;
  logic [31:0] rd_6;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;
  reg [31:0] rd_6_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;
      rd_6_stage_1 <= rd_6;


    end

  end


  // Data processing units...
  // selector_bright_gauss_blur_2_rd0_select
  logic [0:0] selector_bright_gauss_blur_2_rd0_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd0_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd0_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd0_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd0_select_out;
  bright_gauss_blur_2_rd0_select selector_bright_gauss_blur_2_rd0_select(.clk(selector_bright_gauss_blur_2_rd0_select_clk), .rst(selector_bright_gauss_blur_2_rd0_select_rst), .d0(selector_bright_gauss_blur_2_rd0_select_d0), .d1(selector_bright_gauss_blur_2_rd0_select_d1), .out(selector_bright_gauss_blur_2_rd0_select_out));
  assign selector_bright_gauss_blur_2_rd0_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd0_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd0_select

  // selector_bright_gauss_blur_2_rd1_select
  logic [0:0] selector_bright_gauss_blur_2_rd1_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd1_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd1_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd1_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd1_select_out;
  bright_gauss_blur_2_rd1_select selector_bright_gauss_blur_2_rd1_select(.clk(selector_bright_gauss_blur_2_rd1_select_clk), .rst(selector_bright_gauss_blur_2_rd1_select_rst), .d0(selector_bright_gauss_blur_2_rd1_select_d0), .d1(selector_bright_gauss_blur_2_rd1_select_d1), .out(selector_bright_gauss_blur_2_rd1_select_out));
  assign selector_bright_gauss_blur_2_rd1_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd1_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd1_select

  // selector_bright_gauss_blur_2_rd2_select
  logic [0:0] selector_bright_gauss_blur_2_rd2_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd2_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd2_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd2_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd2_select_out;
  bright_gauss_blur_2_rd2_select selector_bright_gauss_blur_2_rd2_select(.clk(selector_bright_gauss_blur_2_rd2_select_clk), .rst(selector_bright_gauss_blur_2_rd2_select_rst), .d0(selector_bright_gauss_blur_2_rd2_select_d0), .d1(selector_bright_gauss_blur_2_rd2_select_d1), .out(selector_bright_gauss_blur_2_rd2_select_out));
  assign selector_bright_gauss_blur_2_rd2_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd2_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd2_select

  // Bindings to bright_gauss_blur_2_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_gauss_blur_2_update_0_read_dummy;

  // bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_clk;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_rst;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_start;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_done;
  bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0 bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0(.clk(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_clk), .rst(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_rst), .start(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_start), .done(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_done));
  assign bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_clk = clk;
  assign bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_rst = rst;
  // Bindings to bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0

  // selector_bright_gauss_blur_2_rd3_select
  logic [0:0] selector_bright_gauss_blur_2_rd3_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd3_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd3_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd3_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd3_select_out;
  bright_gauss_blur_2_rd3_select selector_bright_gauss_blur_2_rd3_select(.clk(selector_bright_gauss_blur_2_rd3_select_clk), .rst(selector_bright_gauss_blur_2_rd3_select_rst), .d0(selector_bright_gauss_blur_2_rd3_select_d0), .d1(selector_bright_gauss_blur_2_rd3_select_d1), .out(selector_bright_gauss_blur_2_rd3_select_out));
  assign selector_bright_gauss_blur_2_rd3_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd3_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd3_select

  // Bindings to bright_gauss_ds_1_update_0_write_wen
    // rd_0
  assign rd_0 = bright_gauss_ds_1_update_0_write_wen;

  // selector_bright_gauss_blur_2_rd4_select
  logic [0:0] selector_bright_gauss_blur_2_rd4_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd4_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd4_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd4_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd4_select_out;
  bright_gauss_blur_2_rd4_select selector_bright_gauss_blur_2_rd4_select(.clk(selector_bright_gauss_blur_2_rd4_select_clk), .rst(selector_bright_gauss_blur_2_rd4_select_rst), .d0(selector_bright_gauss_blur_2_rd4_select_d0), .d1(selector_bright_gauss_blur_2_rd4_select_d1), .out(selector_bright_gauss_blur_2_rd4_select_out));
  assign selector_bright_gauss_blur_2_rd4_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd4_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd4_select

  // selector_bright_laplace_diff_1_rd0_select
  logic [0:0] selector_bright_laplace_diff_1_rd0_select_clk;
  logic [0:0] selector_bright_laplace_diff_1_rd0_select_rst;
  logic [31:0] selector_bright_laplace_diff_1_rd0_select_d0;
  logic [31:0] selector_bright_laplace_diff_1_rd0_select_d1;
  logic [31:0] selector_bright_laplace_diff_1_rd0_select_out;
  bright_laplace_diff_1_rd0_select selector_bright_laplace_diff_1_rd0_select(.clk(selector_bright_laplace_diff_1_rd0_select_clk), .rst(selector_bright_laplace_diff_1_rd0_select_rst), .d0(selector_bright_laplace_diff_1_rd0_select_d0), .d1(selector_bright_laplace_diff_1_rd0_select_d1), .out(selector_bright_laplace_diff_1_rd0_select_out));
  assign selector_bright_laplace_diff_1_rd0_select_clk = clk;
  assign selector_bright_laplace_diff_1_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_diff_1_rd0_select

  // selector_bright_gauss_blur_2_rd5_select
  logic [0:0] selector_bright_gauss_blur_2_rd5_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd5_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd5_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd5_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd5_select_out;
  bright_gauss_blur_2_rd5_select selector_bright_gauss_blur_2_rd5_select(.clk(selector_bright_gauss_blur_2_rd5_select_clk), .rst(selector_bright_gauss_blur_2_rd5_select_rst), .d0(selector_bright_gauss_blur_2_rd5_select_d0), .d1(selector_bright_gauss_blur_2_rd5_select_d1), .out(selector_bright_gauss_blur_2_rd5_select_out));
  assign selector_bright_gauss_blur_2_rd5_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd5_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd5_select

  // selector_bright_gauss_blur_2_rd6_select
  logic [0:0] selector_bright_gauss_blur_2_rd6_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd6_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd6_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd6_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd6_select_out;
  bright_gauss_blur_2_rd6_select selector_bright_gauss_blur_2_rd6_select(.clk(selector_bright_gauss_blur_2_rd6_select_clk), .rst(selector_bright_gauss_blur_2_rd6_select_rst), .d0(selector_bright_gauss_blur_2_rd6_select_d0), .d1(selector_bright_gauss_blur_2_rd6_select_d1), .out(selector_bright_gauss_blur_2_rd6_select_out));
  assign selector_bright_gauss_blur_2_rd6_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd6_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd6_select

  // selector_bright_gauss_blur_2_rd7_select
  logic [0:0] selector_bright_gauss_blur_2_rd7_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd7_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd7_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd7_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd7_select_out;
  bright_gauss_blur_2_rd7_select selector_bright_gauss_blur_2_rd7_select(.clk(selector_bright_gauss_blur_2_rd7_select_clk), .rst(selector_bright_gauss_blur_2_rd7_select_rst), .d0(selector_bright_gauss_blur_2_rd7_select_d0), .d1(selector_bright_gauss_blur_2_rd7_select_d1), .out(selector_bright_gauss_blur_2_rd7_select_out));
  assign selector_bright_gauss_blur_2_rd7_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd7_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd7_select

  // selector_bright_gauss_blur_2_rd8_select
  logic [0:0] selector_bright_gauss_blur_2_rd8_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd8_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd8_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd8_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd8_select_out;
  bright_gauss_blur_2_rd8_select selector_bright_gauss_blur_2_rd8_select(.clk(selector_bright_gauss_blur_2_rd8_select_clk), .rst(selector_bright_gauss_blur_2_rd8_select_rst), .d0(selector_bright_gauss_blur_2_rd8_select_d0), .d1(selector_bright_gauss_blur_2_rd8_select_d1), .out(selector_bright_gauss_blur_2_rd8_select_out));
  assign selector_bright_gauss_blur_2_rd8_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd8_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd8_select

  // Bindings to bright_gauss_ds_1_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_gauss_ds_1_update_0_write_wdata;

  // selector_bright_laplace_us_0_rd0_select
  logic [0:0] selector_bright_laplace_us_0_rd0_select_clk;
  logic [0:0] selector_bright_laplace_us_0_rd0_select_rst;
  logic [31:0] selector_bright_laplace_us_0_rd0_select_d0;
  logic [31:0] selector_bright_laplace_us_0_rd0_select_d1;
  logic [31:0] selector_bright_laplace_us_0_rd0_select_out;
  bright_laplace_us_0_rd0_select selector_bright_laplace_us_0_rd0_select(.clk(selector_bright_laplace_us_0_rd0_select_clk), .rst(selector_bright_laplace_us_0_rd0_select_rst), .d0(selector_bright_laplace_us_0_rd0_select_d0), .d1(selector_bright_laplace_us_0_rd0_select_d1), .out(selector_bright_laplace_us_0_rd0_select_out));
  assign selector_bright_laplace_us_0_rd0_select_clk = clk;
  assign selector_bright_laplace_us_0_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_us_0_rd0_select

  // Bindings to bright_gauss_blur_2_update_0_read_rdata
    // wr_3
  assign bright_gauss_blur_2_update_0_read_rdata = rd_2;

  // Bindings to bright_laplace_diff_1_update_0_read_dummy
    // rd_4
  assign rd_4 = bright_laplace_diff_1_update_0_read_dummy;

  // Bindings to bright_laplace_diff_1_update_0_read_rdata
    // wr_5
  assign bright_laplace_diff_1_update_0_read_rdata = rd_4;

  // Bindings to bright_laplace_us_0_update_0_read_dummy
    // rd_6
  assign rd_6 = bright_laplace_us_0_update_0_read_dummy;

  // Bindings to bright_laplace_us_0_update_0_read_rdata
    // wr_7
  assign bright_laplace_us_0_update_0_read_rdata = rd_6;

  // bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9_clk;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9_rst;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9_start;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9_done;
  bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9 bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9(.clk(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9_clk), .rst(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9_rst), .start(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9_start), .done(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9_done));
  assign bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9_clk = clk;
  assign bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9_rst = rst;
  // Bindings to bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_9

  // bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0_clk;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0_rst;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0_start;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0_done;
  bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0 bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0(.clk(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0_clk), .rst(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0_rst), .start(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0_start), .done(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0_done));
  assign bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0_clk = clk;
  assign bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0_rst = rst;
  // Bindings to bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0



endmodule


module sr_buffer_32_24(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 24;

  reg [31:0] data [23:0];

  reg [31:0] rdata_d;

  reg [4:0] waddr;

  wire [4:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module bright_gauss_blur_3_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 29;
    end
  end

endmodule


module bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_24 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_24 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16



endmodule


module sr_buffer_32_54(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 54;

  reg [31:0] data [53:0];

  reg [31:0] rdata_d;

  reg [5:0] waddr;

  wire [5:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module bright_gauss_blur_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 56;
    end
  end

endmodule


module bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_54 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52



endmodule


module bright_gauss_blur_3_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module bright_gauss_blur_3_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 55;
    end
  end

endmodule


module bright_gauss_blur_3_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 28;
    end
  end

endmodule


module bright_gauss_blur_3_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module bright_gauss_blur_3_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_gauss_ds_2_update_0_write_wen(output [0:0] bright_gauss_ds_2_update_0_write_wen);

endmodule


module bright_laplace_us_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (-1 + d1 == 0) ? ((80 - floord(d0, 2))) : (d1 == 0) ? (56) : ((-1 - d1) % 2 == 0 && -3 + d1 >= 0) ? ((80 - floord(d0, 2))) : ((-d1) % 2 == 0 && -2 + d1 >= 0) ? (56) : 0;
    end
  end

endmodule


module bright_gauss_blur_3_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (23 - d0 >= 0) ? (27) : (-24 + d0 == 0) ? (27) : 0;
    end
  end

endmodule


module bright_gauss_blur_3_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (23 - d0 >= 0) ? (54) : (-24 + d0 == 0) ? (54) : 0;
    end
  end

endmodule


module in_wire_bright_gauss_ds_2_update_0_write_wdata(output [31:0] bright_gauss_ds_2_update_0_write_wdata);

endmodule


module in_wire_bright_gauss_blur_3_update_0_read_dummy(output [287:0] bright_gauss_blur_3_update_0_read_dummy);

endmodule


module out_wire_bright_gauss_blur_3_update_0_read_rdata(input [287:0] bright_gauss_blur_3_update_0_read_rdata);

endmodule


module in_wire_bright_laplace_diff_2_update_0_read_dummy(output [31:0] bright_laplace_diff_2_update_0_read_dummy);

endmodule


module out_wire_bright_laplace_diff_2_update_0_read_rdata(input [31:0] bright_laplace_diff_2_update_0_read_rdata);

endmodule


module in_wire_bright_laplace_us_1_update_0_read_dummy(output [31:0] bright_laplace_us_1_update_0_read_dummy);

endmodule


module out_wire_bright_laplace_us_1_update_0_read_rdata(input [31:0] bright_laplace_us_1_update_0_read_rdata);

endmodule


module bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24



endmodule


module bright_gauss_ds_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_gauss_ds_2_update_0_write_wen, input [31:0] bright_gauss_ds_2_update_0_write_wdata, input [287:0] bright_gauss_blur_3_update_0_read_dummy, output [287:0] bright_gauss_blur_3_update_0_read_rdata, input [31:0] bright_laplace_diff_2_update_0_read_dummy, output [31:0] bright_laplace_diff_2_update_0_read_rdata, input [31:0] bright_laplace_us_1_update_0_read_dummy, output [31:0] bright_laplace_us_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;
  logic [31:0] rd_6;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;
  reg [31:0] rd_6_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;
      rd_6_stage_1 <= rd_6;


    end

  end


  // Data processing units...
  // bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_clk;
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_rst;
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_start;
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_done;
  bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10 bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10(.clk(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_clk), .rst(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_rst), .start(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_start), .done(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_done));
  assign bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_clk = clk;
  assign bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10

  // selector_bright_gauss_blur_3_rd3_select
  logic [0:0] selector_bright_gauss_blur_3_rd3_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd3_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd3_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd3_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd3_select_out;
  bright_gauss_blur_3_rd3_select selector_bright_gauss_blur_3_rd3_select(.clk(selector_bright_gauss_blur_3_rd3_select_clk), .rst(selector_bright_gauss_blur_3_rd3_select_rst), .d0(selector_bright_gauss_blur_3_rd3_select_d0), .d1(selector_bright_gauss_blur_3_rd3_select_d1), .out(selector_bright_gauss_blur_3_rd3_select_out));
  assign selector_bright_gauss_blur_3_rd3_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd3_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd3_select

  // selector_bright_gauss_blur_3_rd2_select
  logic [0:0] selector_bright_gauss_blur_3_rd2_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd2_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd2_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd2_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd2_select_out;
  bright_gauss_blur_3_rd2_select selector_bright_gauss_blur_3_rd2_select(.clk(selector_bright_gauss_blur_3_rd2_select_clk), .rst(selector_bright_gauss_blur_3_rd2_select_rst), .d0(selector_bright_gauss_blur_3_rd2_select_d0), .d1(selector_bright_gauss_blur_3_rd2_select_d1), .out(selector_bright_gauss_blur_3_rd2_select_out));
  assign selector_bright_gauss_blur_3_rd2_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd2_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd2_select

  // selector_bright_gauss_blur_3_rd1_select
  logic [0:0] selector_bright_gauss_blur_3_rd1_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd1_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd1_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd1_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd1_select_out;
  bright_gauss_blur_3_rd1_select selector_bright_gauss_blur_3_rd1_select(.clk(selector_bright_gauss_blur_3_rd1_select_clk), .rst(selector_bright_gauss_blur_3_rd1_select_rst), .d0(selector_bright_gauss_blur_3_rd1_select_d0), .d1(selector_bright_gauss_blur_3_rd1_select_d1), .out(selector_bright_gauss_blur_3_rd1_select_out));
  assign selector_bright_gauss_blur_3_rd1_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd1_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd1_select

  // selector_bright_gauss_blur_3_rd0_select
  logic [0:0] selector_bright_gauss_blur_3_rd0_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd0_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd0_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd0_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd0_select_out;
  bright_gauss_blur_3_rd0_select selector_bright_gauss_blur_3_rd0_select(.clk(selector_bright_gauss_blur_3_rd0_select_clk), .rst(selector_bright_gauss_blur_3_rd0_select_rst), .d0(selector_bright_gauss_blur_3_rd0_select_d0), .d1(selector_bright_gauss_blur_3_rd0_select_d1), .out(selector_bright_gauss_blur_3_rd0_select_out));
  assign selector_bright_gauss_blur_3_rd0_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd0_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd0_select

  // bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_clk;
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_rst;
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_start;
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_done;
  bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0 bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0(.clk(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_clk), .rst(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_rst), .start(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_start), .done(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_done));
  assign bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_clk = clk;
  assign bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_rst = rst;
  // Bindings to bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0

  // selector_bright_gauss_blur_3_rd4_select
  logic [0:0] selector_bright_gauss_blur_3_rd4_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd4_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd4_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd4_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd4_select_out;
  bright_gauss_blur_3_rd4_select selector_bright_gauss_blur_3_rd4_select(.clk(selector_bright_gauss_blur_3_rd4_select_clk), .rst(selector_bright_gauss_blur_3_rd4_select_rst), .d0(selector_bright_gauss_blur_3_rd4_select_d0), .d1(selector_bright_gauss_blur_3_rd4_select_d1), .out(selector_bright_gauss_blur_3_rd4_select_out));
  assign selector_bright_gauss_blur_3_rd4_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd4_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd4_select

  // selector_bright_gauss_blur_3_rd6_select
  logic [0:0] selector_bright_gauss_blur_3_rd6_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd6_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd6_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd6_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd6_select_out;
  bright_gauss_blur_3_rd6_select selector_bright_gauss_blur_3_rd6_select(.clk(selector_bright_gauss_blur_3_rd6_select_clk), .rst(selector_bright_gauss_blur_3_rd6_select_rst), .d0(selector_bright_gauss_blur_3_rd6_select_d0), .d1(selector_bright_gauss_blur_3_rd6_select_d1), .out(selector_bright_gauss_blur_3_rd6_select_out));
  assign selector_bright_gauss_blur_3_rd6_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd6_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd6_select

  // selector_bright_gauss_blur_3_rd5_select
  logic [0:0] selector_bright_gauss_blur_3_rd5_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd5_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd5_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd5_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd5_select_out;
  bright_gauss_blur_3_rd5_select selector_bright_gauss_blur_3_rd5_select(.clk(selector_bright_gauss_blur_3_rd5_select_clk), .rst(selector_bright_gauss_blur_3_rd5_select_rst), .d0(selector_bright_gauss_blur_3_rd5_select_d0), .d1(selector_bright_gauss_blur_3_rd5_select_d1), .out(selector_bright_gauss_blur_3_rd5_select_out));
  assign selector_bright_gauss_blur_3_rd5_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd5_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd5_select

  // selector_bright_gauss_blur_3_rd7_select
  logic [0:0] selector_bright_gauss_blur_3_rd7_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd7_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd7_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd7_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd7_select_out;
  bright_gauss_blur_3_rd7_select selector_bright_gauss_blur_3_rd7_select(.clk(selector_bright_gauss_blur_3_rd7_select_clk), .rst(selector_bright_gauss_blur_3_rd7_select_rst), .d0(selector_bright_gauss_blur_3_rd7_select_d0), .d1(selector_bright_gauss_blur_3_rd7_select_d1), .out(selector_bright_gauss_blur_3_rd7_select_out));
  assign selector_bright_gauss_blur_3_rd7_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd7_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd7_select

  // selector_bright_gauss_blur_3_rd8_select
  logic [0:0] selector_bright_gauss_blur_3_rd8_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd8_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd8_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd8_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd8_select_out;
  bright_gauss_blur_3_rd8_select selector_bright_gauss_blur_3_rd8_select(.clk(selector_bright_gauss_blur_3_rd8_select_clk), .rst(selector_bright_gauss_blur_3_rd8_select_rst), .d0(selector_bright_gauss_blur_3_rd8_select_d0), .d1(selector_bright_gauss_blur_3_rd8_select_d1), .out(selector_bright_gauss_blur_3_rd8_select_out));
  assign selector_bright_gauss_blur_3_rd8_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd8_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd8_select

  // selector_bright_laplace_us_1_rd0_select
  logic [0:0] selector_bright_laplace_us_1_rd0_select_clk;
  logic [0:0] selector_bright_laplace_us_1_rd0_select_rst;
  logic [31:0] selector_bright_laplace_us_1_rd0_select_d0;
  logic [31:0] selector_bright_laplace_us_1_rd0_select_d1;
  logic [31:0] selector_bright_laplace_us_1_rd0_select_out;
  bright_laplace_us_1_rd0_select selector_bright_laplace_us_1_rd0_select(.clk(selector_bright_laplace_us_1_rd0_select_clk), .rst(selector_bright_laplace_us_1_rd0_select_rst), .d0(selector_bright_laplace_us_1_rd0_select_d0), .d1(selector_bright_laplace_us_1_rd0_select_d1), .out(selector_bright_laplace_us_1_rd0_select_out));
  assign selector_bright_laplace_us_1_rd0_select_clk = clk;
  assign selector_bright_laplace_us_1_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_us_1_rd0_select

  // Bindings to bright_gauss_ds_2_update_0_write_wen
    // rd_0
  assign rd_0 = bright_gauss_ds_2_update_0_write_wen;

  // selector_bright_laplace_diff_2_rd0_select
  logic [0:0] selector_bright_laplace_diff_2_rd0_select_clk;
  logic [0:0] selector_bright_laplace_diff_2_rd0_select_rst;
  logic [31:0] selector_bright_laplace_diff_2_rd0_select_d0;
  logic [31:0] selector_bright_laplace_diff_2_rd0_select_d1;
  logic [31:0] selector_bright_laplace_diff_2_rd0_select_out;
  bright_laplace_diff_2_rd0_select selector_bright_laplace_diff_2_rd0_select(.clk(selector_bright_laplace_diff_2_rd0_select_clk), .rst(selector_bright_laplace_diff_2_rd0_select_rst), .d0(selector_bright_laplace_diff_2_rd0_select_d0), .d1(selector_bright_laplace_diff_2_rd0_select_d1), .out(selector_bright_laplace_diff_2_rd0_select_out));
  assign selector_bright_laplace_diff_2_rd0_select_clk = clk;
  assign selector_bright_laplace_diff_2_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_diff_2_rd0_select

  // Bindings to bright_gauss_ds_2_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_gauss_ds_2_update_0_write_wdata;

  // Bindings to bright_gauss_blur_3_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_gauss_blur_3_update_0_read_dummy;

  // Bindings to bright_gauss_blur_3_update_0_read_rdata
    // wr_3
  assign bright_gauss_blur_3_update_0_read_rdata = rd_2;

  // Bindings to bright_laplace_diff_2_update_0_read_dummy
    // rd_4
  assign rd_4 = bright_laplace_diff_2_update_0_read_dummy;

  // Bindings to bright_laplace_diff_2_update_0_read_rdata
    // wr_5
  assign bright_laplace_diff_2_update_0_read_rdata = rd_4;

  // Bindings to bright_laplace_us_1_update_0_read_dummy
    // rd_6
  assign rd_6 = bright_laplace_us_1_update_0_read_dummy;

  // Bindings to bright_laplace_us_1_update_0_read_rdata
    // wr_7
  assign bright_laplace_us_1_update_0_read_rdata = rd_6;



endmodule


module bright_laplace_us_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = ((-1 - d1) % 2 == 0 && 23 - d0 >= 0) ? ((12 - floord(2*d0, 4))) : 0;
    end
  end

endmodule


module in_wire_bright_gauss_ds_3_update_0_write_wen(output [0:0] bright_gauss_ds_3_update_0_write_wen);

endmodule


module bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_gauss_ds_3_update_0_write_wdata(output [31:0] bright_gauss_ds_3_update_0_write_wdata);

endmodule


module in_wire_bright_laplace_us_2_update_0_read_dummy(output [31:0] bright_laplace_us_2_update_0_read_dummy);

endmodule


module out_wire_bright_laplace_us_2_update_0_read_rdata(input [31:0] bright_laplace_us_2_update_0_read_rdata);

endmodule


module in_wire_fused_level_3_update_0_read_dummy(output [31:0] fused_level_3_update_0_read_dummy);

endmodule


module out_wire_fused_level_3_update_0_read_rdata(input [31:0] fused_level_3_update_0_read_rdata);

endmodule


module bright_gauss_ds_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] fused_level_3_update_0_read_dummy, input [0:0] bright_gauss_ds_3_update_0_write_wen, input [31:0] bright_gauss_ds_3_update_0_write_wdata, input [31:0] bright_laplace_us_2_update_0_read_dummy, output [31:0] bright_laplace_us_2_update_0_read_rdata, output [31:0] fused_level_3_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_clk;
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_rst;
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_start;
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_done;
  bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0 bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0(.clk(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_clk), .rst(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_rst), .start(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_start), .done(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_done));
  assign bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_clk = clk;
  assign bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_rst = rst;
  // Bindings to bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0

  // bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_done;
  bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1 bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1(.clk(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_clk), .rst(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_rst), .start(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_start), .done(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_done));
  assign bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_clk = clk;
  assign bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1

  // selector_bright_laplace_us_2_rd0_select
  logic [0:0] selector_bright_laplace_us_2_rd0_select_clk;
  logic [0:0] selector_bright_laplace_us_2_rd0_select_rst;
  logic [31:0] selector_bright_laplace_us_2_rd0_select_d0;
  logic [31:0] selector_bright_laplace_us_2_rd0_select_d1;
  logic [31:0] selector_bright_laplace_us_2_rd0_select_out;
  bright_laplace_us_2_rd0_select selector_bright_laplace_us_2_rd0_select(.clk(selector_bright_laplace_us_2_rd0_select_clk), .rst(selector_bright_laplace_us_2_rd0_select_rst), .d0(selector_bright_laplace_us_2_rd0_select_d0), .d1(selector_bright_laplace_us_2_rd0_select_d1), .out(selector_bright_laplace_us_2_rd0_select_out));
  assign selector_bright_laplace_us_2_rd0_select_clk = clk;
  assign selector_bright_laplace_us_2_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_us_2_rd0_select

  // Bindings to fused_level_3_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_3_update_0_read_dummy;

  // Bindings to bright_gauss_ds_3_update_0_write_wen
    // rd_0
  assign rd_0 = bright_gauss_ds_3_update_0_write_wen;

  // selector_fused_level_3_rd0_select
  logic [0:0] selector_fused_level_3_rd0_select_clk;
  logic [0:0] selector_fused_level_3_rd0_select_rst;
  logic [31:0] selector_fused_level_3_rd0_select_d0;
  logic [31:0] selector_fused_level_3_rd0_select_d1;
  logic [31:0] selector_fused_level_3_rd0_select_out;
  fused_level_3_rd0_select selector_fused_level_3_rd0_select(.clk(selector_fused_level_3_rd0_select_clk), .rst(selector_fused_level_3_rd0_select_rst), .d0(selector_fused_level_3_rd0_select_d0), .d1(selector_fused_level_3_rd0_select_d1), .out(selector_fused_level_3_rd0_select_out));
  assign selector_fused_level_3_rd0_select_clk = clk;
  assign selector_fused_level_3_rd0_select_rst = rst;
  // Bindings to selector_fused_level_3_rd0_select

  // Bindings to bright_gauss_ds_3_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_gauss_ds_3_update_0_write_wdata;

  // Bindings to bright_laplace_us_2_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_laplace_us_2_update_0_read_dummy;

  // Bindings to bright_laplace_us_2_update_0_read_rdata
    // wr_3
  assign bright_laplace_us_2_update_0_read_rdata = rd_2;

  // Bindings to fused_level_3_update_0_read_rdata
    // wr_5
  assign fused_level_3_update_0_read_rdata = rd_4;



endmodule


module bright_weights_normed(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] fused_level_0_update_0_read_dummy, output [31:0] fused_level_0_update_0_read_rdata, input [0:0] bright_weights_normed_update_0_write_wen, input [31:0] bright_weights_normed_update_0_write_wdata, input [287:0] bright_weights_normed_gauss_blur_1_update_0_read_dummy, output [287:0] bright_weights_normed_gauss_blur_1_update_0_read_rdata);

  logic [31:0] rd_4;
  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_4_stage_1;
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_4_stage_1 <= rd_4;
      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to fused_level_0_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_0_update_0_read_dummy;

  // Bindings to fused_level_0_update_0_read_rdata
    // wr_5
  assign fused_level_0_update_0_read_rdata = rd_4;

  // bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_clk;
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_rst;
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_start;
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_done;
  bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9 bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9(.clk(bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_clk), .rst(bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_rst), .start(bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_start), .done(bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_done));
  assign bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_clk = clk;
  assign bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_rst = rst;
  // Bindings to bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9

  // bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_clk;
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_rst;
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_start;
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_done;
  bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0 bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0(.clk(bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_clk), .rst(bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_rst), .start(bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_start), .done(bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_done));
  assign bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_clk = clk;
  assign bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_rst = rst;
  // Bindings to bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0

  // selector_fused_level_0_rd0_select
  logic [0:0] selector_fused_level_0_rd0_select_clk;
  logic [0:0] selector_fused_level_0_rd0_select_rst;
  logic [31:0] selector_fused_level_0_rd0_select_d0;
  logic [31:0] selector_fused_level_0_rd0_select_d1;
  logic [31:0] selector_fused_level_0_rd0_select_out;
  fused_level_0_rd0_select selector_fused_level_0_rd0_select(.clk(selector_fused_level_0_rd0_select_clk), .rst(selector_fused_level_0_rd0_select_rst), .d0(selector_fused_level_0_rd0_select_d0), .d1(selector_fused_level_0_rd0_select_d1), .out(selector_fused_level_0_rd0_select_out));
  assign selector_fused_level_0_rd0_select_clk = clk;
  assign selector_fused_level_0_rd0_select_rst = rst;
  // Bindings to selector_fused_level_0_rd0_select

  // selector_bright_weights_normed_gauss_blur_1_rd0_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd0_select_out;
  bright_weights_normed_gauss_blur_1_rd0_select selector_bright_weights_normed_gauss_blur_1_rd0_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd0_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd0_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd0_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd0_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd0_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd0_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd0_select

  // selector_bright_weights_normed_gauss_blur_1_rd1_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd1_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd1_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd1_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd1_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd1_select_out;
  bright_weights_normed_gauss_blur_1_rd1_select selector_bright_weights_normed_gauss_blur_1_rd1_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd1_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd1_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd1_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd1_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd1_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd1_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd1_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd1_select

  // selector_bright_weights_normed_gauss_blur_1_rd2_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd2_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd2_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd2_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd2_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd2_select_out;
  bright_weights_normed_gauss_blur_1_rd2_select selector_bright_weights_normed_gauss_blur_1_rd2_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd2_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd2_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd2_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd2_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd2_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd2_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd2_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd2_select

  // selector_bright_weights_normed_gauss_blur_1_rd3_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd3_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd3_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd3_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd3_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd3_select_out;
  bright_weights_normed_gauss_blur_1_rd3_select selector_bright_weights_normed_gauss_blur_1_rd3_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd3_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd3_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd3_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd3_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd3_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd3_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd3_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd3_select

  // selector_bright_weights_normed_gauss_blur_1_rd4_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd4_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd4_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd4_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd4_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd4_select_out;
  bright_weights_normed_gauss_blur_1_rd4_select selector_bright_weights_normed_gauss_blur_1_rd4_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd4_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd4_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd4_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd4_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd4_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd4_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd4_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd4_select

  // selector_bright_weights_normed_gauss_blur_1_rd6_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd6_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd6_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd6_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd6_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd6_select_out;
  bright_weights_normed_gauss_blur_1_rd6_select selector_bright_weights_normed_gauss_blur_1_rd6_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd6_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd6_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd6_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd6_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd6_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd6_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd6_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd6_select

  // selector_bright_weights_normed_gauss_blur_1_rd5_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd5_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd5_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd5_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd5_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd5_select_out;
  bright_weights_normed_gauss_blur_1_rd5_select selector_bright_weights_normed_gauss_blur_1_rd5_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd5_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd5_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd5_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd5_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd5_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd5_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd5_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd5_select

  // Bindings to bright_weights_normed_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_normed_update_0_write_wen;

  // selector_bright_weights_normed_gauss_blur_1_rd7_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd7_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd7_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd7_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd7_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd7_select_out;
  bright_weights_normed_gauss_blur_1_rd7_select selector_bright_weights_normed_gauss_blur_1_rd7_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd7_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd7_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd7_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd7_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd7_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd7_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd7_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd7_select

  // selector_bright_weights_normed_gauss_blur_1_rd8_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd8_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd8_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd8_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd8_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd8_select_out;
  bright_weights_normed_gauss_blur_1_rd8_select selector_bright_weights_normed_gauss_blur_1_rd8_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd8_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd8_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd8_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd8_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd8_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd8_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd8_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd8_select

  // Bindings to bright_weights_normed_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_normed_update_0_write_wdata;

  // Bindings to bright_weights_normed_gauss_blur_1_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_gauss_blur_1_update_0_read_dummy;

  // Bindings to bright_weights_normed_gauss_blur_1_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_gauss_blur_1_update_0_read_rdata = rd_2;



endmodule


module bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_weights_normed_gauss_blur_1_update_0_write_wen(output [0:0] bright_weights_normed_gauss_blur_1_update_0_write_wen);

endmodule


module bright_weights_normed_gauss_ds_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_weights_normed_gauss_blur_1_update_0_write_wdata(output [31:0] bright_weights_normed_gauss_blur_1_update_0_write_wdata);

endmodule


module in_wire_bright_weights_normed_gauss_ds_1_update_0_read_dummy(output [31:0] bright_weights_normed_gauss_ds_1_update_0_read_dummy);

endmodule


module out_wire_bright_weights_normed_gauss_ds_1_update_0_read_rdata(input [31:0] bright_weights_normed_gauss_ds_1_update_0_read_rdata);

endmodule


module bright_weights_normed_gauss_blur_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] bright_weights_normed_gauss_blur_1_update_0_write_wdata, input [0:0] bright_weights_normed_gauss_blur_1_update_0_write_wen, input [31:0] bright_weights_normed_gauss_ds_1_update_0_read_dummy, output [31:0] bright_weights_normed_gauss_ds_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1
  logic [0:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_done;
  bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1 bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1(.clk(bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_clk), .rst(bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_rst), .start(bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_start), .done(bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_done));
  assign bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_clk = clk;
  assign bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1

  // selector_bright_weights_normed_gauss_ds_1_rd0_select
  logic [0:0] selector_bright_weights_normed_gauss_ds_1_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_ds_1_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_ds_1_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_ds_1_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_ds_1_rd0_select_out;
  bright_weights_normed_gauss_ds_1_rd0_select selector_bright_weights_normed_gauss_ds_1_rd0_select(.clk(selector_bright_weights_normed_gauss_ds_1_rd0_select_clk), .rst(selector_bright_weights_normed_gauss_ds_1_rd0_select_rst), .d0(selector_bright_weights_normed_gauss_ds_1_rd0_select_d0), .d1(selector_bright_weights_normed_gauss_ds_1_rd0_select_d1), .out(selector_bright_weights_normed_gauss_ds_1_rd0_select_out));
  assign selector_bright_weights_normed_gauss_ds_1_rd0_select_clk = clk;
  assign selector_bright_weights_normed_gauss_ds_1_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_ds_1_rd0_select

  // Bindings to bright_weights_normed_gauss_blur_1_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_normed_gauss_blur_1_update_0_write_wdata;

  // Bindings to bright_weights_normed_gauss_blur_1_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_normed_gauss_blur_1_update_0_write_wen;

  // Bindings to bright_weights_normed_gauss_ds_1_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_gauss_ds_1_update_0_read_dummy;

  // Bindings to bright_weights_normed_gauss_ds_1_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_gauss_ds_1_update_0_read_rdata = rd_2;



endmodule


module bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_weights_normed_gauss_blur_2_update_0_write_wen(output [0:0] bright_weights_normed_gauss_blur_2_update_0_write_wen);

endmodule


module bright_weights_normed_gauss_ds_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_weights_normed_gauss_blur_2_update_0_write_wdata(output [31:0] bright_weights_normed_gauss_blur_2_update_0_write_wdata);

endmodule


module in_wire_bright_weights_normed_gauss_ds_2_update_0_read_dummy(output [31:0] bright_weights_normed_gauss_ds_2_update_0_read_dummy);

endmodule


module out_wire_bright_weights_normed_gauss_ds_2_update_0_read_rdata(input [31:0] bright_weights_normed_gauss_ds_2_update_0_read_rdata);

endmodule


module bright_weights_normed_gauss_blur_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_weights_normed_gauss_blur_2_update_0_write_wen, input [31:0] bright_weights_normed_gauss_blur_2_update_0_write_wdata, input [31:0] bright_weights_normed_gauss_ds_2_update_0_read_dummy, output [31:0] bright_weights_normed_gauss_ds_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to bright_weights_normed_gauss_blur_2_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_normed_gauss_blur_2_update_0_write_wen;

  // Bindings to bright_weights_normed_gauss_blur_2_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_normed_gauss_blur_2_update_0_write_wdata;

  // bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1
  logic [0:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_done;
  bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1 bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1(.clk(bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_clk), .rst(bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_rst), .start(bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_start), .done(bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_done));
  assign bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_clk = clk;
  assign bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1

  // selector_bright_weights_normed_gauss_ds_2_rd0_select
  logic [0:0] selector_bright_weights_normed_gauss_ds_2_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_ds_2_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_ds_2_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_ds_2_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_ds_2_rd0_select_out;
  bright_weights_normed_gauss_ds_2_rd0_select selector_bright_weights_normed_gauss_ds_2_rd0_select(.clk(selector_bright_weights_normed_gauss_ds_2_rd0_select_clk), .rst(selector_bright_weights_normed_gauss_ds_2_rd0_select_rst), .d0(selector_bright_weights_normed_gauss_ds_2_rd0_select_d0), .d1(selector_bright_weights_normed_gauss_ds_2_rd0_select_d1), .out(selector_bright_weights_normed_gauss_ds_2_rd0_select_out));
  assign selector_bright_weights_normed_gauss_ds_2_rd0_select_clk = clk;
  assign selector_bright_weights_normed_gauss_ds_2_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_ds_2_rd0_select

  // Bindings to bright_weights_normed_gauss_ds_2_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_gauss_ds_2_update_0_read_dummy;

  // Bindings to bright_weights_normed_gauss_ds_2_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_gauss_ds_2_update_0_read_rdata = rd_2;



endmodule


module in_wire_bright_weights_normed_gauss_blur_3_update_0_write_wen(output [0:0] bright_weights_normed_gauss_blur_3_update_0_write_wen);

endmodule


module bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module bright_weights_normed_gauss_ds_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_weights_normed_gauss_blur_3_update_0_write_wdata(output [31:0] bright_weights_normed_gauss_blur_3_update_0_write_wdata);

endmodule


module in_wire_bright_weights_normed_gauss_ds_3_update_0_read_dummy(output [31:0] bright_weights_normed_gauss_ds_3_update_0_read_dummy);

endmodule


module out_wire_bright_weights_normed_gauss_ds_3_update_0_read_rdata(input [31:0] bright_weights_normed_gauss_ds_3_update_0_read_rdata);

endmodule


module bright_weights_normed_gauss_blur_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_weights_normed_gauss_blur_3_update_0_write_wen, input [31:0] bright_weights_normed_gauss_blur_3_update_0_write_wdata, input [31:0] bright_weights_normed_gauss_ds_3_update_0_read_dummy, output [31:0] bright_weights_normed_gauss_ds_3_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to bright_weights_normed_gauss_blur_3_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_normed_gauss_blur_3_update_0_write_wen;

  // Bindings to bright_weights_normed_gauss_blur_3_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_normed_gauss_blur_3_update_0_write_wdata;

  // bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1
  logic [0:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_done;
  bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1 bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1(.clk(bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_clk), .rst(bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_rst), .start(bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_start), .done(bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_done));
  assign bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_clk = clk;
  assign bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1

  // selector_bright_weights_normed_gauss_ds_3_rd0_select
  logic [0:0] selector_bright_weights_normed_gauss_ds_3_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_ds_3_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_ds_3_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_ds_3_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_ds_3_rd0_select_out;
  bright_weights_normed_gauss_ds_3_rd0_select selector_bright_weights_normed_gauss_ds_3_rd0_select(.clk(selector_bright_weights_normed_gauss_ds_3_rd0_select_clk), .rst(selector_bright_weights_normed_gauss_ds_3_rd0_select_rst), .d0(selector_bright_weights_normed_gauss_ds_3_rd0_select_d0), .d1(selector_bright_weights_normed_gauss_ds_3_rd0_select_d1), .out(selector_bright_weights_normed_gauss_ds_3_rd0_select_out));
  assign selector_bright_weights_normed_gauss_ds_3_rd0_select_clk = clk;
  assign selector_bright_weights_normed_gauss_ds_3_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_ds_3_rd0_select

  // Bindings to bright_weights_normed_gauss_ds_3_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_gauss_ds_3_update_0_read_dummy;

  // Bindings to bright_weights_normed_gauss_ds_3_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_gauss_ds_3_update_0_read_rdata = rd_2;



endmodule


module in_wire_bright_weights_normed_gauss_ds_3_update_0_write_wdata(output [31:0] bright_weights_normed_gauss_ds_3_update_0_write_wdata);

endmodule


module bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_52 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_52 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16



endmodule


module in_wire_bright_weights_normed_gauss_ds_3_update_0_write_wen(output [0:0] bright_weights_normed_gauss_ds_3_update_0_write_wen);

endmodule


module dark(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] dark_update_0_write_wdata, output [31:0] dark_weights_update_0_read_rdata, output [31:0] dark_laplace_diff_0_update_0_read_rdata, output [287:0] dark_gauss_blur_1_update_0_read_rdata, input [31:0] dark_laplace_diff_0_update_0_read_dummy, input [31:0] dark_weights_update_0_read_dummy, input [287:0] dark_gauss_blur_1_update_0_read_dummy, input [0:0] dark_update_0_write_wen);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;
  logic [31:0] rd_6;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;
  reg [31:0] rd_6_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;
      rd_6_stage_1 <= rd_6;


    end

  end


  // Data processing units...
  // dark_dark_update_0_write0_merged_banks_10
  logic [0:0] dark_dark_update_0_write0_merged_banks_10_clk;
  logic [0:0] dark_dark_update_0_write0_merged_banks_10_rst;
  logic [0:0] dark_dark_update_0_write0_merged_banks_10_start;
  logic [0:0] dark_dark_update_0_write0_merged_banks_10_done;
  dark_dark_update_0_write0_merged_banks_10 dark_dark_update_0_write0_merged_banks_10(.clk(dark_dark_update_0_write0_merged_banks_10_clk), .rst(dark_dark_update_0_write0_merged_banks_10_rst), .start(dark_dark_update_0_write0_merged_banks_10_start), .done(dark_dark_update_0_write0_merged_banks_10_done));
  assign dark_dark_update_0_write0_merged_banks_10_clk = clk;
  assign dark_dark_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to dark_dark_update_0_write0_merged_banks_10

  // Bindings to dark_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_update_0_write_wdata;

  // selector_dark_gauss_blur_1_rd0_select
  logic [0:0] selector_dark_gauss_blur_1_rd0_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd0_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd0_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd0_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd0_select_out;
  dark_gauss_blur_1_rd0_select selector_dark_gauss_blur_1_rd0_select(.clk(selector_dark_gauss_blur_1_rd0_select_clk), .rst(selector_dark_gauss_blur_1_rd0_select_rst), .d0(selector_dark_gauss_blur_1_rd0_select_d0), .d1(selector_dark_gauss_blur_1_rd0_select_d1), .out(selector_dark_gauss_blur_1_rd0_select_out));
  assign selector_dark_gauss_blur_1_rd0_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd0_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd0_select

  // selector_dark_gauss_blur_1_rd3_select
  logic [0:0] selector_dark_gauss_blur_1_rd3_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd3_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd3_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd3_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd3_select_out;
  dark_gauss_blur_1_rd3_select selector_dark_gauss_blur_1_rd3_select(.clk(selector_dark_gauss_blur_1_rd3_select_clk), .rst(selector_dark_gauss_blur_1_rd3_select_rst), .d0(selector_dark_gauss_blur_1_rd3_select_d0), .d1(selector_dark_gauss_blur_1_rd3_select_d1), .out(selector_dark_gauss_blur_1_rd3_select_out));
  assign selector_dark_gauss_blur_1_rd3_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd3_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd3_select

  // selector_dark_gauss_blur_1_rd2_select
  logic [0:0] selector_dark_gauss_blur_1_rd2_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd2_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd2_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd2_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd2_select_out;
  dark_gauss_blur_1_rd2_select selector_dark_gauss_blur_1_rd2_select(.clk(selector_dark_gauss_blur_1_rd2_select_clk), .rst(selector_dark_gauss_blur_1_rd2_select_rst), .d0(selector_dark_gauss_blur_1_rd2_select_d0), .d1(selector_dark_gauss_blur_1_rd2_select_d1), .out(selector_dark_gauss_blur_1_rd2_select_out));
  assign selector_dark_gauss_blur_1_rd2_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd2_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd2_select

  // Bindings to dark_weights_update_0_read_rdata
    // wr_7
  assign dark_weights_update_0_read_rdata = rd_6;

  // Bindings to dark_laplace_diff_0_update_0_read_rdata
    // wr_5
  assign dark_laplace_diff_0_update_0_read_rdata = rd_4;

  // Bindings to dark_gauss_blur_1_update_0_read_rdata
    // wr_3
  assign dark_gauss_blur_1_update_0_read_rdata = rd_2;

  // Bindings to dark_laplace_diff_0_update_0_read_dummy
    // rd_4
  assign rd_4 = dark_laplace_diff_0_update_0_read_dummy;

  // Bindings to dark_weights_update_0_read_dummy
    // rd_6
  assign rd_6 = dark_weights_update_0_read_dummy;

  // Bindings to dark_gauss_blur_1_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_gauss_blur_1_update_0_read_dummy;

  // Bindings to dark_update_0_write_wen
    // rd_0
  assign rd_0 = dark_update_0_write_wen;

  // selector_dark_weights_rd0_select
  logic [0:0] selector_dark_weights_rd0_select_clk;
  logic [0:0] selector_dark_weights_rd0_select_rst;
  logic [31:0] selector_dark_weights_rd0_select_d0;
  logic [31:0] selector_dark_weights_rd0_select_d1;
  logic [31:0] selector_dark_weights_rd0_select_out;
  dark_weights_rd0_select selector_dark_weights_rd0_select(.clk(selector_dark_weights_rd0_select_clk), .rst(selector_dark_weights_rd0_select_rst), .d0(selector_dark_weights_rd0_select_d0), .d1(selector_dark_weights_rd0_select_d1), .out(selector_dark_weights_rd0_select_out));
  assign selector_dark_weights_rd0_select_clk = clk;
  assign selector_dark_weights_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_rd0_select

  // selector_dark_laplace_diff_0_rd0_select
  logic [0:0] selector_dark_laplace_diff_0_rd0_select_clk;
  logic [0:0] selector_dark_laplace_diff_0_rd0_select_rst;
  logic [31:0] selector_dark_laplace_diff_0_rd0_select_d0;
  logic [31:0] selector_dark_laplace_diff_0_rd0_select_d1;
  logic [31:0] selector_dark_laplace_diff_0_rd0_select_out;
  dark_laplace_diff_0_rd0_select selector_dark_laplace_diff_0_rd0_select(.clk(selector_dark_laplace_diff_0_rd0_select_clk), .rst(selector_dark_laplace_diff_0_rd0_select_rst), .d0(selector_dark_laplace_diff_0_rd0_select_d0), .d1(selector_dark_laplace_diff_0_rd0_select_d1), .out(selector_dark_laplace_diff_0_rd0_select_out));
  assign selector_dark_laplace_diff_0_rd0_select_clk = clk;
  assign selector_dark_laplace_diff_0_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_diff_0_rd0_select

  // selector_dark_gauss_blur_1_rd8_select
  logic [0:0] selector_dark_gauss_blur_1_rd8_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd8_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd8_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd8_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd8_select_out;
  dark_gauss_blur_1_rd8_select selector_dark_gauss_blur_1_rd8_select(.clk(selector_dark_gauss_blur_1_rd8_select_clk), .rst(selector_dark_gauss_blur_1_rd8_select_rst), .d0(selector_dark_gauss_blur_1_rd8_select_d0), .d1(selector_dark_gauss_blur_1_rd8_select_d1), .out(selector_dark_gauss_blur_1_rd8_select_out));
  assign selector_dark_gauss_blur_1_rd8_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd8_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd8_select

  // selector_dark_gauss_blur_1_rd7_select
  logic [0:0] selector_dark_gauss_blur_1_rd7_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd7_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd7_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd7_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd7_select_out;
  dark_gauss_blur_1_rd7_select selector_dark_gauss_blur_1_rd7_select(.clk(selector_dark_gauss_blur_1_rd7_select_clk), .rst(selector_dark_gauss_blur_1_rd7_select_rst), .d0(selector_dark_gauss_blur_1_rd7_select_d0), .d1(selector_dark_gauss_blur_1_rd7_select_d1), .out(selector_dark_gauss_blur_1_rd7_select_out));
  assign selector_dark_gauss_blur_1_rd7_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd7_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd7_select

  // selector_dark_gauss_blur_1_rd6_select
  logic [0:0] selector_dark_gauss_blur_1_rd6_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd6_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd6_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd6_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd6_select_out;
  dark_gauss_blur_1_rd6_select selector_dark_gauss_blur_1_rd6_select(.clk(selector_dark_gauss_blur_1_rd6_select_clk), .rst(selector_dark_gauss_blur_1_rd6_select_rst), .d0(selector_dark_gauss_blur_1_rd6_select_d0), .d1(selector_dark_gauss_blur_1_rd6_select_d1), .out(selector_dark_gauss_blur_1_rd6_select_out));
  assign selector_dark_gauss_blur_1_rd6_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd6_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd6_select

  // selector_dark_gauss_blur_1_rd5_select
  logic [0:0] selector_dark_gauss_blur_1_rd5_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd5_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd5_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd5_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd5_select_out;
  dark_gauss_blur_1_rd5_select selector_dark_gauss_blur_1_rd5_select(.clk(selector_dark_gauss_blur_1_rd5_select_clk), .rst(selector_dark_gauss_blur_1_rd5_select_rst), .d0(selector_dark_gauss_blur_1_rd5_select_d0), .d1(selector_dark_gauss_blur_1_rd5_select_d1), .out(selector_dark_gauss_blur_1_rd5_select_out));
  assign selector_dark_gauss_blur_1_rd5_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd5_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd5_select

  // selector_dark_gauss_blur_1_rd4_select
  logic [0:0] selector_dark_gauss_blur_1_rd4_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd4_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd4_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd4_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd4_select_out;
  dark_gauss_blur_1_rd4_select selector_dark_gauss_blur_1_rd4_select(.clk(selector_dark_gauss_blur_1_rd4_select_clk), .rst(selector_dark_gauss_blur_1_rd4_select_rst), .d0(selector_dark_gauss_blur_1_rd4_select_d0), .d1(selector_dark_gauss_blur_1_rd4_select_d1), .out(selector_dark_gauss_blur_1_rd4_select_out));
  assign selector_dark_gauss_blur_1_rd4_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd4_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd4_select

  // selector_dark_gauss_blur_1_rd1_select
  logic [0:0] selector_dark_gauss_blur_1_rd1_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd1_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd1_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd1_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd1_select_out;
  dark_gauss_blur_1_rd1_select selector_dark_gauss_blur_1_rd1_select(.clk(selector_dark_gauss_blur_1_rd1_select_clk), .rst(selector_dark_gauss_blur_1_rd1_select_rst), .d0(selector_dark_gauss_blur_1_rd1_select_d0), .d1(selector_dark_gauss_blur_1_rd1_select_d1), .out(selector_dark_gauss_blur_1_rd1_select_out));
  assign selector_dark_gauss_blur_1_rd1_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd1_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd1_select

  // dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0
  logic [0:0] dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_clk;
  logic [0:0] dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_rst;
  logic [0:0] dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_start;
  logic [0:0] dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_done;
  dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0 dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0(.clk(dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_clk), .rst(dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_rst), .start(dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_start), .done(dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_done));
  assign dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_clk = clk;
  assign dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_rst = rst;
  // Bindings to dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0



endmodule


module dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_gauss_blur_1_update_0_write_wen(output [0:0] dark_gauss_blur_1_update_0_write_wen);

endmodule


module dark_gauss_ds_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_gauss_blur_1_update_0_write_wdata(output [31:0] dark_gauss_blur_1_update_0_write_wdata);

endmodule


module in_wire_dark_gauss_ds_1_update_0_read_dummy(output [31:0] dark_gauss_ds_1_update_0_read_dummy);

endmodule


module out_wire_dark_gauss_ds_1_update_0_read_rdata(input [31:0] dark_gauss_ds_1_update_0_read_rdata);

endmodule


module dark_weights(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_weights_update_0_write_wen, input [31:0] dark_weights_update_0_write_wdata, input [31:0] weight_sums_update_0_read_dummy, input [31:0] dark_weights_normed_update_0_read_dummy, output [31:0] dark_weights_normed_update_0_read_rdata, output [31:0] weight_sums_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // dark_weights_dark_weights_update_0_write0_merged_banks_2
  logic [0:0] dark_weights_dark_weights_update_0_write0_merged_banks_2_clk;
  logic [0:0] dark_weights_dark_weights_update_0_write0_merged_banks_2_rst;
  logic [0:0] dark_weights_dark_weights_update_0_write0_merged_banks_2_start;
  logic [0:0] dark_weights_dark_weights_update_0_write0_merged_banks_2_done;
  dark_weights_dark_weights_update_0_write0_merged_banks_2 dark_weights_dark_weights_update_0_write0_merged_banks_2(.clk(dark_weights_dark_weights_update_0_write0_merged_banks_2_clk), .rst(dark_weights_dark_weights_update_0_write0_merged_banks_2_rst), .start(dark_weights_dark_weights_update_0_write0_merged_banks_2_start), .done(dark_weights_dark_weights_update_0_write0_merged_banks_2_done));
  assign dark_weights_dark_weights_update_0_write0_merged_banks_2_clk = clk;
  assign dark_weights_dark_weights_update_0_write0_merged_banks_2_rst = rst;
  // Bindings to dark_weights_dark_weights_update_0_write0_merged_banks_2

  // Bindings to dark_weights_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_update_0_write_wen;

  // selector_dark_weights_normed_rd0_select
  logic [0:0] selector_dark_weights_normed_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_rd0_select_out;
  dark_weights_normed_rd0_select selector_dark_weights_normed_rd0_select(.clk(selector_dark_weights_normed_rd0_select_clk), .rst(selector_dark_weights_normed_rd0_select_rst), .d0(selector_dark_weights_normed_rd0_select_d0), .d1(selector_dark_weights_normed_rd0_select_d1), .out(selector_dark_weights_normed_rd0_select_out));
  assign selector_dark_weights_normed_rd0_select_clk = clk;
  assign selector_dark_weights_normed_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_rd0_select

  // selector_weight_sums_rd0_select
  logic [0:0] selector_weight_sums_rd0_select_clk;
  logic [0:0] selector_weight_sums_rd0_select_rst;
  logic [31:0] selector_weight_sums_rd0_select_d0;
  logic [31:0] selector_weight_sums_rd0_select_d1;
  logic [31:0] selector_weight_sums_rd0_select_out;
  weight_sums_rd0_select selector_weight_sums_rd0_select(.clk(selector_weight_sums_rd0_select_clk), .rst(selector_weight_sums_rd0_select_rst), .d0(selector_weight_sums_rd0_select_d0), .d1(selector_weight_sums_rd0_select_d1), .out(selector_weight_sums_rd0_select_out));
  assign selector_weight_sums_rd0_select_clk = clk;
  assign selector_weight_sums_rd0_select_rst = rst;
  // Bindings to selector_weight_sums_rd0_select

  // Bindings to dark_weights_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_update_0_write_wdata;

  // Bindings to weight_sums_update_0_read_dummy
    // rd_4
  assign rd_4 = weight_sums_update_0_read_dummy;

  // Bindings to dark_weights_normed_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_weights_normed_update_0_read_dummy;

  // Bindings to dark_weights_normed_update_0_read_rdata
    // wr_3
  assign dark_weights_normed_update_0_read_rdata = rd_2;

  // Bindings to weight_sums_update_0_read_rdata
    // wr_5
  assign weight_sums_update_0_read_rdata = rd_4;



endmodule


module dark_weights_normed_gauss_ds_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] fused_level_1_update_0_read_rdata, input [31:0] fused_level_1_update_0_read_dummy, output [287:0] dark_weights_normed_gauss_blur_2_update_0_read_rdata, input [31:0] dark_weights_normed_gauss_ds_1_update_0_write_wdata, input [0:0] dark_weights_normed_gauss_ds_1_update_0_write_wen, input [287:0] dark_weights_normed_gauss_blur_2_update_0_read_dummy);

  logic [31:0] rd_4;
  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_4_stage_1;
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_4_stage_1 <= rd_4;
      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0
  logic [0:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_clk;
  logic [0:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_rst;
  logic [0:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_start;
  logic [0:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_done;
  dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0 dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0(.clk(dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_clk), .rst(dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_rst), .start(dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_start), .done(dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_done));
  assign dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_clk = clk;
  assign dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0_rst = rst;
  // Bindings to dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0

  // selector_dark_weights_normed_gauss_blur_2_rd4_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd4_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd4_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd4_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd4_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd4_select_out;
  dark_weights_normed_gauss_blur_2_rd4_select selector_dark_weights_normed_gauss_blur_2_rd4_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd4_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd4_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd4_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd4_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd4_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd4_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd4_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd4_select

  // selector_dark_weights_normed_gauss_blur_2_rd7_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd7_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd7_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd7_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd7_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd7_select_out;
  dark_weights_normed_gauss_blur_2_rd7_select selector_dark_weights_normed_gauss_blur_2_rd7_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd7_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd7_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd7_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd7_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd7_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd7_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd7_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd7_select

  // Bindings to fused_level_1_update_0_read_rdata
    // wr_5
  assign fused_level_1_update_0_read_rdata = rd_4;

  // selector_dark_weights_normed_gauss_blur_2_rd8_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd8_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd8_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd8_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd8_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd8_select_out;
  dark_weights_normed_gauss_blur_2_rd8_select selector_dark_weights_normed_gauss_blur_2_rd8_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd8_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd8_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd8_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd8_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd8_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd8_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd8_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd8_select

  // Bindings to fused_level_1_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_1_update_0_read_dummy;

  // Bindings to dark_weights_normed_gauss_blur_2_update_0_read_rdata
    // wr_3
  assign dark_weights_normed_gauss_blur_2_update_0_read_rdata = rd_2;

  // Bindings to dark_weights_normed_gauss_ds_1_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_normed_gauss_ds_1_update_0_write_wdata;

  // Bindings to dark_weights_normed_gauss_ds_1_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_normed_gauss_ds_1_update_0_write_wen;

  // selector_dark_weights_normed_gauss_blur_2_rd6_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd6_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd6_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd6_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd6_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd6_select_out;
  dark_weights_normed_gauss_blur_2_rd6_select selector_dark_weights_normed_gauss_blur_2_rd6_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd6_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd6_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd6_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd6_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd6_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd6_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd6_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd6_select

  // Bindings to dark_weights_normed_gauss_blur_2_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_weights_normed_gauss_blur_2_update_0_read_dummy;

  // selector_dark_weights_normed_gauss_blur_2_rd0_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd0_select_out;
  dark_weights_normed_gauss_blur_2_rd0_select selector_dark_weights_normed_gauss_blur_2_rd0_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd0_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd0_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd0_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd0_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd0_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd0_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd0_select

  // selector_fused_level_1_rd0_select
  logic [0:0] selector_fused_level_1_rd0_select_clk;
  logic [0:0] selector_fused_level_1_rd0_select_rst;
  logic [31:0] selector_fused_level_1_rd0_select_d0;
  logic [31:0] selector_fused_level_1_rd0_select_d1;
  logic [31:0] selector_fused_level_1_rd0_select_out;
  fused_level_1_rd0_select selector_fused_level_1_rd0_select(.clk(selector_fused_level_1_rd0_select_clk), .rst(selector_fused_level_1_rd0_select_rst), .d0(selector_fused_level_1_rd0_select_d0), .d1(selector_fused_level_1_rd0_select_d1), .out(selector_fused_level_1_rd0_select_out));
  assign selector_fused_level_1_rd0_select_clk = clk;
  assign selector_fused_level_1_rd0_select_rst = rst;
  // Bindings to selector_fused_level_1_rd0_select

  // selector_dark_weights_normed_gauss_blur_2_rd1_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd1_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd1_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd1_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd1_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd1_select_out;
  dark_weights_normed_gauss_blur_2_rd1_select selector_dark_weights_normed_gauss_blur_2_rd1_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd1_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd1_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd1_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd1_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd1_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd1_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd1_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd1_select

  // selector_dark_weights_normed_gauss_blur_2_rd2_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd2_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd2_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd2_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd2_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd2_select_out;
  dark_weights_normed_gauss_blur_2_rd2_select selector_dark_weights_normed_gauss_blur_2_rd2_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd2_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd2_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd2_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd2_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd2_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd2_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd2_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd2_select

  // selector_dark_weights_normed_gauss_blur_2_rd3_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd3_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd3_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd3_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd3_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd3_select_out;
  dark_weights_normed_gauss_blur_2_rd3_select selector_dark_weights_normed_gauss_blur_2_rd3_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd3_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd3_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd3_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd3_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd3_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd3_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd3_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd3_select

  // selector_dark_weights_normed_gauss_blur_2_rd5_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd5_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd5_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd5_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd5_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd5_select_out;
  dark_weights_normed_gauss_blur_2_rd5_select selector_dark_weights_normed_gauss_blur_2_rd5_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd5_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd5_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd5_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd5_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd5_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd5_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd5_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd5_select

  // dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9
  logic [0:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_clk;
  logic [0:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_rst;
  logic [0:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_start;
  logic [0:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_done;
  dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9 dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9(.clk(dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_clk), .rst(dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_rst), .start(dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_start), .done(dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_done));
  assign dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_clk = clk;
  assign dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9_rst = rst;
  // Bindings to dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9



endmodule


module final_merged_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] final_merged_1_update_0_write_wen, input [31:0] final_merged_1_update_0_write_wdata, input [31:0] final_merged_0_update_0_read_dummy, output [31:0] final_merged_0_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to final_merged_1_update_0_write_wen
    // rd_0
  assign rd_0 = final_merged_1_update_0_write_wen;

  // final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0
  logic [0:0] final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_clk;
  logic [0:0] final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_rst;
  logic [0:0] final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_start;
  logic [0:0] final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_done;
  final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0 final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0(.clk(final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_clk), .rst(final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_rst), .start(final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_start), .done(final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_done));
  assign final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_clk = clk;
  assign final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_rst = rst;
  // Bindings to final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0

  // Bindings to final_merged_1_update_0_write_wdata
    // rd_1
  assign rd_1 = final_merged_1_update_0_write_wdata;

  // selector_final_merged_0_rd0_select
  logic [0:0] selector_final_merged_0_rd0_select_clk;
  logic [0:0] selector_final_merged_0_rd0_select_rst;
  logic [31:0] selector_final_merged_0_rd0_select_d0;
  logic [31:0] selector_final_merged_0_rd0_select_d1;
  logic [31:0] selector_final_merged_0_rd0_select_out;
  final_merged_0_rd0_select selector_final_merged_0_rd0_select(.clk(selector_final_merged_0_rd0_select_clk), .rst(selector_final_merged_0_rd0_select_rst), .d0(selector_final_merged_0_rd0_select_d0), .d1(selector_final_merged_0_rd0_select_d1), .out(selector_final_merged_0_rd0_select_out));
  assign selector_final_merged_0_rd0_select_clk = clk;
  assign selector_final_merged_0_rd0_select_rst = rst;
  // Bindings to selector_final_merged_0_rd0_select

  // Bindings to final_merged_0_update_0_read_dummy
    // rd_2
  assign rd_2 = final_merged_0_update_0_read_dummy;

  // Bindings to final_merged_0_update_0_read_rdata
    // wr_3
  assign final_merged_0_update_0_read_rdata = rd_2;



endmodule


module final_merged_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] final_merged_2_update_0_write_wdata, input [0:0] final_merged_2_update_0_write_wen, input [31:0] final_merged_1_update_0_read_dummy, output [31:0] final_merged_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0
  logic [0:0] final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_clk;
  logic [0:0] final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_rst;
  logic [0:0] final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_start;
  logic [0:0] final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_done;
  final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0 final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0(.clk(final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_clk), .rst(final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_rst), .start(final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_start), .done(final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_done));
  assign final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_clk = clk;
  assign final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_rst = rst;
  // Bindings to final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0

  // selector_final_merged_1_rd0_select
  logic [0:0] selector_final_merged_1_rd0_select_clk;
  logic [0:0] selector_final_merged_1_rd0_select_rst;
  logic [31:0] selector_final_merged_1_rd0_select_d0;
  logic [31:0] selector_final_merged_1_rd0_select_d1;
  logic [31:0] selector_final_merged_1_rd0_select_out;
  final_merged_1_rd0_select selector_final_merged_1_rd0_select(.clk(selector_final_merged_1_rd0_select_clk), .rst(selector_final_merged_1_rd0_select_rst), .d0(selector_final_merged_1_rd0_select_d0), .d1(selector_final_merged_1_rd0_select_d1), .out(selector_final_merged_1_rd0_select_out));
  assign selector_final_merged_1_rd0_select_clk = clk;
  assign selector_final_merged_1_rd0_select_rst = rst;
  // Bindings to selector_final_merged_1_rd0_select

  // Bindings to final_merged_2_update_0_write_wdata
    // rd_1
  assign rd_1 = final_merged_2_update_0_write_wdata;

  // Bindings to final_merged_2_update_0_write_wen
    // rd_0
  assign rd_0 = final_merged_2_update_0_write_wen;

  // Bindings to final_merged_1_update_0_read_dummy
    // rd_2
  assign rd_2 = final_merged_1_update_0_read_dummy;

  // Bindings to final_merged_1_update_0_read_rdata
    // wr_3
  assign final_merged_1_update_0_read_rdata = rd_2;



endmodule


module fused_level_0_fused_level_0_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module fused_level_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_weights_normed_gauss_blur_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module dark_gauss_ds_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module dark_weights_normed_gauss_ds_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_weights_normed_gauss_ds_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module dark_laplace_us_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module fused_level_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module final_merged_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module final_merged_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module final_merged_0_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module pyramid_synthetic_exposure_fusion_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module sr_buffer_32_1(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 1;

  reg [31:0] data [0:0];

  reg [31:0] rdata_d;

  reg [0:0] waddr;

  wire [0:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module sr_buffer_32_108(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 108;

  reg [31:0] data [107:0];

  reg [31:0] rdata_d;

  reg [6:0] waddr;

  wire [6:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module bright_laplace_diff_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] fused_level_1_update_0_read_dummy, input [0:0] bright_laplace_diff_1_update_0_write_wen, input [31:0] bright_laplace_diff_1_update_0_write_wdata, output [31:0] fused_level_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to fused_level_1_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_1_update_0_read_dummy;

  // bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1
  logic [0:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_done;
  bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1 bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1(.clk(bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_clk), .rst(bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_rst), .start(bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_start), .done(bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_done));
  assign bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_clk = clk;
  assign bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1

  // selector_fused_level_1_rd0_select
  logic [0:0] selector_fused_level_1_rd0_select_clk;
  logic [0:0] selector_fused_level_1_rd0_select_rst;
  logic [31:0] selector_fused_level_1_rd0_select_d0;
  logic [31:0] selector_fused_level_1_rd0_select_d1;
  logic [31:0] selector_fused_level_1_rd0_select_out;
  fused_level_1_rd0_select selector_fused_level_1_rd0_select(.clk(selector_fused_level_1_rd0_select_clk), .rst(selector_fused_level_1_rd0_select_rst), .d0(selector_fused_level_1_rd0_select_d0), .d1(selector_fused_level_1_rd0_select_d1), .out(selector_fused_level_1_rd0_select_out));
  assign selector_fused_level_1_rd0_select_clk = clk;
  assign selector_fused_level_1_rd0_select_rst = rst;
  // Bindings to selector_fused_level_1_rd0_select

  // Bindings to bright_laplace_diff_1_update_0_write_wen
    // rd_0
  assign rd_0 = bright_laplace_diff_1_update_0_write_wen;

  // Bindings to bright_laplace_diff_1_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_laplace_diff_1_update_0_write_wdata;

  // Bindings to fused_level_1_update_0_read_rdata
    // wr_3
  assign fused_level_1_update_0_read_rdata = rd_2;



endmodule


module bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_laplace_diff_2_update_0_write_wen(output [0:0] bright_laplace_diff_2_update_0_write_wen);

endmodule


module in_wire_bright_laplace_diff_2_update_0_write_wdata(output [31:0] bright_laplace_diff_2_update_0_write_wdata);

endmodule


module in_wire_fused_level_2_update_0_read_dummy(output [31:0] fused_level_2_update_0_read_dummy);

endmodule


module out_wire_fused_level_2_update_0_read_rdata(input [31:0] fused_level_2_update_0_read_rdata);

endmodule


module bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_108 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_108 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16



endmodule


module bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_278 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212



endmodule


module bright_weights_normed_gauss_ds_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] bright_weights_normed_gauss_ds_3_update_0_write_wdata, output [31:0] fused_level_3_update_0_read_rdata, input [31:0] fused_level_3_update_0_read_dummy, input [0:0] bright_weights_normed_gauss_ds_3_update_0_write_wen);

  logic [0:0] rd_0;
  logic [31:0] rd_2;
  logic [31:0] rd_1;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_2_stage_1;
  reg [31:0] rd_1_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_2_stage_1 <= rd_2;
      rd_1_stage_1 <= rd_1;


    end

  end


  // Data processing units...
  // Bindings to bright_weights_normed_gauss_ds_3_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_normed_gauss_ds_3_update_0_write_wdata;

  // Bindings to fused_level_3_update_0_read_rdata
    // wr_3
  assign fused_level_3_update_0_read_rdata = rd_2;

  // Bindings to fused_level_3_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_3_update_0_read_dummy;

  // selector_fused_level_3_rd0_select
  logic [0:0] selector_fused_level_3_rd0_select_clk;
  logic [0:0] selector_fused_level_3_rd0_select_rst;
  logic [31:0] selector_fused_level_3_rd0_select_d0;
  logic [31:0] selector_fused_level_3_rd0_select_d1;
  logic [31:0] selector_fused_level_3_rd0_select_out;
  fused_level_3_rd0_select selector_fused_level_3_rd0_select(.clk(selector_fused_level_3_rd0_select_clk), .rst(selector_fused_level_3_rd0_select_rst), .d0(selector_fused_level_3_rd0_select_d0), .d1(selector_fused_level_3_rd0_select_d1), .out(selector_fused_level_3_rd0_select_out));
  assign selector_fused_level_3_rd0_select_clk = clk;
  assign selector_fused_level_3_rd0_select_rst = rst;
  // Bindings to selector_fused_level_3_rd0_select

  // Bindings to bright_weights_normed_gauss_ds_3_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_normed_gauss_ds_3_update_0_write_wen;

  // bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1
  logic [0:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_done;
  bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1 bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1(.clk(bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_clk), .rst(bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_rst), .start(bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_start), .done(bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_done));
  assign bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_clk = clk;
  assign bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1



endmodule


module dark_gauss_blur_2_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (51 - d0 >= 0) ? (110) : (-52 + d0 == 0) ? (110) : 0;
    end
  end

endmodule


module dark_gauss_blur_2_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 57;
    end
  end

endmodule


module dark_gauss_blur_2_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module dark_gauss_blur_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 112;
    end
  end

endmodule


module dark_gauss_blur_2_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 111;
    end
  end

endmodule


module dark_laplace_us_0_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (d1 == 0 && -98 + d0 >= 0) ? (335) : (-98 + d1 >= 0) ? ((329 - floord(d0, 2))) : (-1 + d1 == 0) ? ((384 - floord(d0, 2))) : (d1 == 0 && 97 - d0 >= 0) ? (336) : ((-d1) % 2 == 0 && -98 + d0 >= 0 && -2 + d1 >= 0 && 96 - d1 >= 0) ? (335) : ((-1 - d1) % 2 == 0 && -3 + d1 >= 0 && 97 - d1 >= 0) ? ((384 - floord(d0, 2))) : ((-d1) % 2 == 0 && 97 - d0 >= 0 && -2 + d1 >= 0 && 96 - d1 >= 0) ? (336) : 0;
    end
  end

endmodule


module dark_gauss_blur_2_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 56;
    end
  end

endmodule


module dark_gauss_blur_2_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module dark_gauss_blur_2_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_gauss_ds_1_update_0_write_wen(output [0:0] dark_gauss_ds_1_update_0_write_wen);

endmodule


module dark_gauss_blur_2_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (51 - d0 >= 0) ? (55) : (-52 + d0 == 0) ? (55) : 0;
    end
  end

endmodule


module dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_24 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_24 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0



endmodule


module in_wire_dark_gauss_blur_2_update_0_read_dummy(output [287:0] dark_gauss_blur_2_update_0_read_dummy);

endmodule


module out_wire_dark_gauss_blur_2_update_0_read_rdata(input [287:0] dark_gauss_blur_2_update_0_read_rdata);

endmodule


module in_wire_dark_gauss_ds_1_update_0_write_wdata(output [31:0] dark_gauss_ds_1_update_0_write_wdata);

endmodule


module in_wire_dark_laplace_diff_1_update_0_read_dummy(output [31:0] dark_laplace_diff_1_update_0_read_dummy);

endmodule


module out_wire_dark_laplace_diff_1_update_0_read_rdata(input [31:0] dark_laplace_diff_1_update_0_read_rdata);

endmodule


module in_wire_dark_laplace_us_0_update_0_read_dummy(output [31:0] dark_laplace_us_0_update_0_read_dummy);

endmodule


module out_wire_dark_laplace_us_0_update_0_read_rdata(input [31:0] dark_laplace_us_0_update_0_read_rdata);

endmodule


module dark_gauss_blur_3_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (23 - d0 >= 0) ? (54) : (-24 + d0 == 0) ? (54) : 0;
    end
  end

endmodule


module dark_gauss_blur_3_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_gauss_blur_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 56;
    end
  end

endmodule


module dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_54 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52



endmodule


module dark_gauss_blur_3_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 29;
    end
  end

endmodule


module dark_gauss_blur_3_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module dark_gauss_blur_3_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 55;
    end
  end

endmodule


module dark_gauss_blur_3_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 28;
    end
  end

endmodule


module dark_gauss_blur_3_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (23 - d0 >= 0) ? (27) : (-24 + d0 == 0) ? (27) : 0;
    end
  end

endmodule


module dark_gauss_blur_3_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module in_wire_dark_gauss_ds_2_update_0_write_wen(output [0:0] dark_gauss_ds_2_update_0_write_wen);

endmodule


module dark_laplace_us_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (-1 + d1 == 0) ? ((80 - floord(d0, 2))) : (d1 == 0) ? (56) : ((-1 - d1) % 2 == 0 && -3 + d1 >= 0) ? ((80 - floord(d0, 2))) : ((-d1) % 2 == 0 && -2 + d1 >= 0) ? (56) : 0;
    end
  end

endmodule


module in_wire_dark_gauss_ds_2_update_0_write_wdata(output [31:0] dark_gauss_ds_2_update_0_write_wdata);

endmodule


module dark_gauss_ds_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_gauss_ds_2_update_0_write_wen, input [31:0] dark_gauss_ds_2_update_0_write_wdata, input [287:0] dark_gauss_blur_3_update_0_read_dummy, output [287:0] dark_gauss_blur_3_update_0_read_rdata, input [31:0] dark_laplace_diff_2_update_0_read_dummy, output [31:0] dark_laplace_diff_2_update_0_read_rdata, input [31:0] dark_laplace_us_1_update_0_read_dummy, output [31:0] dark_laplace_us_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;
  logic [31:0] rd_6;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;
  reg [31:0] rd_6_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;
      rd_6_stage_1 <= rd_6;


    end

  end


  // Data processing units...
  // selector_dark_gauss_blur_3_rd2_select
  logic [0:0] selector_dark_gauss_blur_3_rd2_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd2_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd2_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd2_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd2_select_out;
  dark_gauss_blur_3_rd2_select selector_dark_gauss_blur_3_rd2_select(.clk(selector_dark_gauss_blur_3_rd2_select_clk), .rst(selector_dark_gauss_blur_3_rd2_select_rst), .d0(selector_dark_gauss_blur_3_rd2_select_d0), .d1(selector_dark_gauss_blur_3_rd2_select_d1), .out(selector_dark_gauss_blur_3_rd2_select_out));
  assign selector_dark_gauss_blur_3_rd2_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd2_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd2_select

  // dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_clk;
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_rst;
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_start;
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_done;
  dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10 dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10(.clk(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_clk), .rst(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_rst), .start(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_start), .done(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_done));
  assign dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_clk = clk;
  assign dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10

  // selector_dark_gauss_blur_3_rd3_select
  logic [0:0] selector_dark_gauss_blur_3_rd3_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd3_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd3_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd3_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd3_select_out;
  dark_gauss_blur_3_rd3_select selector_dark_gauss_blur_3_rd3_select(.clk(selector_dark_gauss_blur_3_rd3_select_clk), .rst(selector_dark_gauss_blur_3_rd3_select_rst), .d0(selector_dark_gauss_blur_3_rd3_select_d0), .d1(selector_dark_gauss_blur_3_rd3_select_d1), .out(selector_dark_gauss_blur_3_rd3_select_out));
  assign selector_dark_gauss_blur_3_rd3_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd3_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd3_select

  // selector_dark_gauss_blur_3_rd1_select
  logic [0:0] selector_dark_gauss_blur_3_rd1_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd1_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd1_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd1_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd1_select_out;
  dark_gauss_blur_3_rd1_select selector_dark_gauss_blur_3_rd1_select(.clk(selector_dark_gauss_blur_3_rd1_select_clk), .rst(selector_dark_gauss_blur_3_rd1_select_rst), .d0(selector_dark_gauss_blur_3_rd1_select_d0), .d1(selector_dark_gauss_blur_3_rd1_select_d1), .out(selector_dark_gauss_blur_3_rd1_select_out));
  assign selector_dark_gauss_blur_3_rd1_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd1_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd1_select

  // selector_dark_gauss_blur_3_rd0_select
  logic [0:0] selector_dark_gauss_blur_3_rd0_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd0_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd0_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd0_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd0_select_out;
  dark_gauss_blur_3_rd0_select selector_dark_gauss_blur_3_rd0_select(.clk(selector_dark_gauss_blur_3_rd0_select_clk), .rst(selector_dark_gauss_blur_3_rd0_select_rst), .d0(selector_dark_gauss_blur_3_rd0_select_d0), .d1(selector_dark_gauss_blur_3_rd0_select_d1), .out(selector_dark_gauss_blur_3_rd0_select_out));
  assign selector_dark_gauss_blur_3_rd0_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd0_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd0_select

  // dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_clk;
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_rst;
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_start;
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_done;
  dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0 dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0(.clk(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_clk), .rst(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_rst), .start(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_start), .done(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_done));
  assign dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_clk = clk;
  assign dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_rst = rst;
  // Bindings to dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0

  // Bindings to dark_gauss_ds_2_update_0_write_wen
    // rd_0
  assign rd_0 = dark_gauss_ds_2_update_0_write_wen;

  // selector_dark_gauss_blur_3_rd4_select
  logic [0:0] selector_dark_gauss_blur_3_rd4_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd4_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd4_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd4_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd4_select_out;
  dark_gauss_blur_3_rd4_select selector_dark_gauss_blur_3_rd4_select(.clk(selector_dark_gauss_blur_3_rd4_select_clk), .rst(selector_dark_gauss_blur_3_rd4_select_rst), .d0(selector_dark_gauss_blur_3_rd4_select_d0), .d1(selector_dark_gauss_blur_3_rd4_select_d1), .out(selector_dark_gauss_blur_3_rd4_select_out));
  assign selector_dark_gauss_blur_3_rd4_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd4_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd4_select

  // selector_dark_gauss_blur_3_rd7_select
  logic [0:0] selector_dark_gauss_blur_3_rd7_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd7_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd7_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd7_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd7_select_out;
  dark_gauss_blur_3_rd7_select selector_dark_gauss_blur_3_rd7_select(.clk(selector_dark_gauss_blur_3_rd7_select_clk), .rst(selector_dark_gauss_blur_3_rd7_select_rst), .d0(selector_dark_gauss_blur_3_rd7_select_d0), .d1(selector_dark_gauss_blur_3_rd7_select_d1), .out(selector_dark_gauss_blur_3_rd7_select_out));
  assign selector_dark_gauss_blur_3_rd7_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd7_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd7_select

  // selector_dark_gauss_blur_3_rd6_select
  logic [0:0] selector_dark_gauss_blur_3_rd6_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd6_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd6_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd6_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd6_select_out;
  dark_gauss_blur_3_rd6_select selector_dark_gauss_blur_3_rd6_select(.clk(selector_dark_gauss_blur_3_rd6_select_clk), .rst(selector_dark_gauss_blur_3_rd6_select_rst), .d0(selector_dark_gauss_blur_3_rd6_select_d0), .d1(selector_dark_gauss_blur_3_rd6_select_d1), .out(selector_dark_gauss_blur_3_rd6_select_out));
  assign selector_dark_gauss_blur_3_rd6_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd6_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd6_select

  // selector_dark_gauss_blur_3_rd5_select
  logic [0:0] selector_dark_gauss_blur_3_rd5_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd5_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd5_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd5_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd5_select_out;
  dark_gauss_blur_3_rd5_select selector_dark_gauss_blur_3_rd5_select(.clk(selector_dark_gauss_blur_3_rd5_select_clk), .rst(selector_dark_gauss_blur_3_rd5_select_rst), .d0(selector_dark_gauss_blur_3_rd5_select_d0), .d1(selector_dark_gauss_blur_3_rd5_select_d1), .out(selector_dark_gauss_blur_3_rd5_select_out));
  assign selector_dark_gauss_blur_3_rd5_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd5_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd5_select

  // selector_dark_laplace_us_1_rd0_select
  logic [0:0] selector_dark_laplace_us_1_rd0_select_clk;
  logic [0:0] selector_dark_laplace_us_1_rd0_select_rst;
  logic [31:0] selector_dark_laplace_us_1_rd0_select_d0;
  logic [31:0] selector_dark_laplace_us_1_rd0_select_d1;
  logic [31:0] selector_dark_laplace_us_1_rd0_select_out;
  dark_laplace_us_1_rd0_select selector_dark_laplace_us_1_rd0_select(.clk(selector_dark_laplace_us_1_rd0_select_clk), .rst(selector_dark_laplace_us_1_rd0_select_rst), .d0(selector_dark_laplace_us_1_rd0_select_d0), .d1(selector_dark_laplace_us_1_rd0_select_d1), .out(selector_dark_laplace_us_1_rd0_select_out));
  assign selector_dark_laplace_us_1_rd0_select_clk = clk;
  assign selector_dark_laplace_us_1_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_us_1_rd0_select

  // selector_dark_gauss_blur_3_rd8_select
  logic [0:0] selector_dark_gauss_blur_3_rd8_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd8_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd8_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd8_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd8_select_out;
  dark_gauss_blur_3_rd8_select selector_dark_gauss_blur_3_rd8_select(.clk(selector_dark_gauss_blur_3_rd8_select_clk), .rst(selector_dark_gauss_blur_3_rd8_select_rst), .d0(selector_dark_gauss_blur_3_rd8_select_d0), .d1(selector_dark_gauss_blur_3_rd8_select_d1), .out(selector_dark_gauss_blur_3_rd8_select_out));
  assign selector_dark_gauss_blur_3_rd8_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd8_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd8_select

  // selector_dark_laplace_diff_2_rd0_select
  logic [0:0] selector_dark_laplace_diff_2_rd0_select_clk;
  logic [0:0] selector_dark_laplace_diff_2_rd0_select_rst;
  logic [31:0] selector_dark_laplace_diff_2_rd0_select_d0;
  logic [31:0] selector_dark_laplace_diff_2_rd0_select_d1;
  logic [31:0] selector_dark_laplace_diff_2_rd0_select_out;
  dark_laplace_diff_2_rd0_select selector_dark_laplace_diff_2_rd0_select(.clk(selector_dark_laplace_diff_2_rd0_select_clk), .rst(selector_dark_laplace_diff_2_rd0_select_rst), .d0(selector_dark_laplace_diff_2_rd0_select_d0), .d1(selector_dark_laplace_diff_2_rd0_select_d1), .out(selector_dark_laplace_diff_2_rd0_select_out));
  assign selector_dark_laplace_diff_2_rd0_select_clk = clk;
  assign selector_dark_laplace_diff_2_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_diff_2_rd0_select

  // Bindings to dark_gauss_ds_2_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_gauss_ds_2_update_0_write_wdata;

  // Bindings to dark_gauss_blur_3_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_gauss_blur_3_update_0_read_dummy;

  // Bindings to dark_gauss_blur_3_update_0_read_rdata
    // wr_3
  assign dark_gauss_blur_3_update_0_read_rdata = rd_2;

  // Bindings to dark_laplace_diff_2_update_0_read_dummy
    // rd_4
  assign rd_4 = dark_laplace_diff_2_update_0_read_dummy;

  // Bindings to dark_laplace_diff_2_update_0_read_rdata
    // wr_5
  assign dark_laplace_diff_2_update_0_read_rdata = rd_4;

  // Bindings to dark_laplace_us_1_update_0_read_dummy
    // rd_6
  assign rd_6 = dark_laplace_us_1_update_0_read_dummy;

  // Bindings to dark_laplace_us_1_update_0_read_rdata
    // wr_7
  assign dark_laplace_us_1_update_0_read_rdata = rd_6;



endmodule


module in_wire_dark_gauss_blur_3_update_0_read_dummy(output [287:0] dark_gauss_blur_3_update_0_read_dummy);

endmodule


module out_wire_dark_gauss_blur_3_update_0_read_rdata(input [287:0] dark_gauss_blur_3_update_0_read_rdata);

endmodule


module in_wire_dark_laplace_diff_2_update_0_read_dummy(output [31:0] dark_laplace_diff_2_update_0_read_dummy);

endmodule


module out_wire_dark_laplace_diff_2_update_0_read_rdata(input [31:0] dark_laplace_diff_2_update_0_read_rdata);

endmodule


module in_wire_dark_laplace_us_1_update_0_read_dummy(output [31:0] dark_laplace_us_1_update_0_read_dummy);

endmodule


module out_wire_dark_laplace_us_1_update_0_read_rdata(input [31:0] dark_laplace_us_1_update_0_read_rdata);

endmodule


module dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24



endmodule


module in_wire_dark_laplace_diff_0_update_0_write_wen(output [0:0] dark_laplace_diff_0_update_0_write_wen);

endmodule


module dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_laplace_diff_0_update_0_write_wdata(output [31:0] dark_laplace_diff_0_update_0_write_wdata);

endmodule


module dark_laplace_diff_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] fused_level_0_update_0_read_dummy, input [0:0] dark_laplace_diff_0_update_0_write_wen, input [31:0] dark_laplace_diff_0_update_0_write_wdata, output [31:0] fused_level_0_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to fused_level_0_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_0_update_0_read_dummy;

  // selector_fused_level_0_rd0_select
  logic [0:0] selector_fused_level_0_rd0_select_clk;
  logic [0:0] selector_fused_level_0_rd0_select_rst;
  logic [31:0] selector_fused_level_0_rd0_select_d0;
  logic [31:0] selector_fused_level_0_rd0_select_d1;
  logic [31:0] selector_fused_level_0_rd0_select_out;
  fused_level_0_rd0_select selector_fused_level_0_rd0_select(.clk(selector_fused_level_0_rd0_select_clk), .rst(selector_fused_level_0_rd0_select_rst), .d0(selector_fused_level_0_rd0_select_d0), .d1(selector_fused_level_0_rd0_select_d1), .out(selector_fused_level_0_rd0_select_out));
  assign selector_fused_level_0_rd0_select_clk = clk;
  assign selector_fused_level_0_rd0_select_rst = rst;
  // Bindings to selector_fused_level_0_rd0_select

  // Bindings to dark_laplace_diff_0_update_0_write_wen
    // rd_0
  assign rd_0 = dark_laplace_diff_0_update_0_write_wen;

  // dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1
  logic [0:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_done;
  dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1 dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1(.clk(dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_clk), .rst(dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_rst), .start(dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_start), .done(dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_done));
  assign dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_clk = clk;
  assign dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1

  // Bindings to dark_laplace_diff_0_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_laplace_diff_0_update_0_write_wdata;

  // Bindings to fused_level_0_update_0_read_rdata
    // wr_3
  assign fused_level_0_update_0_read_rdata = rd_2;



endmodule


module dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module dark_laplace_diff_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_laplace_diff_1_update_0_write_wen, input [31:0] fused_level_1_update_0_read_dummy, input [31:0] dark_laplace_diff_1_update_0_write_wdata, output [31:0] fused_level_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1
  logic [0:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_done;
  dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1 dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1(.clk(dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_clk), .rst(dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_rst), .start(dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_start), .done(dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_done));
  assign dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_clk = clk;
  assign dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1

  // Bindings to dark_laplace_diff_1_update_0_write_wen
    // rd_0
  assign rd_0 = dark_laplace_diff_1_update_0_write_wen;

  // Bindings to fused_level_1_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_1_update_0_read_dummy;

  // selector_fused_level_1_rd0_select
  logic [0:0] selector_fused_level_1_rd0_select_clk;
  logic [0:0] selector_fused_level_1_rd0_select_rst;
  logic [31:0] selector_fused_level_1_rd0_select_d0;
  logic [31:0] selector_fused_level_1_rd0_select_d1;
  logic [31:0] selector_fused_level_1_rd0_select_out;
  fused_level_1_rd0_select selector_fused_level_1_rd0_select(.clk(selector_fused_level_1_rd0_select_clk), .rst(selector_fused_level_1_rd0_select_rst), .d0(selector_fused_level_1_rd0_select_d0), .d1(selector_fused_level_1_rd0_select_d1), .out(selector_fused_level_1_rd0_select_out));
  assign selector_fused_level_1_rd0_select_clk = clk;
  assign selector_fused_level_1_rd0_select_rst = rst;
  // Bindings to selector_fused_level_1_rd0_select

  // Bindings to dark_laplace_diff_1_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_laplace_diff_1_update_0_write_wdata;

  // Bindings to fused_level_1_update_0_read_rdata
    // wr_3
  assign fused_level_1_update_0_read_rdata = rd_2;



endmodule


module dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_laplace_diff_2_update_0_write_wen(output [0:0] dark_laplace_diff_2_update_0_write_wen);

endmodule


module in_wire_dark_laplace_diff_2_update_0_write_wdata(output [31:0] dark_laplace_diff_2_update_0_write_wdata);

endmodule


module dark_laplace_diff_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] fused_level_2_update_0_read_dummy, input [0:0] dark_laplace_diff_2_update_0_write_wen, input [31:0] dark_laplace_diff_2_update_0_write_wdata, output [31:0] fused_level_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to fused_level_2_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_2_update_0_read_dummy;

  // Bindings to dark_laplace_diff_2_update_0_write_wen
    // rd_0
  assign rd_0 = dark_laplace_diff_2_update_0_write_wen;

  // dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1
  logic [0:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_done;
  dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1 dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1(.clk(dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_clk), .rst(dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_rst), .start(dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_start), .done(dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_done));
  assign dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_clk = clk;
  assign dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1

  // selector_fused_level_2_rd0_select
  logic [0:0] selector_fused_level_2_rd0_select_clk;
  logic [0:0] selector_fused_level_2_rd0_select_rst;
  logic [31:0] selector_fused_level_2_rd0_select_d0;
  logic [31:0] selector_fused_level_2_rd0_select_d1;
  logic [31:0] selector_fused_level_2_rd0_select_out;
  fused_level_2_rd0_select selector_fused_level_2_rd0_select(.clk(selector_fused_level_2_rd0_select_clk), .rst(selector_fused_level_2_rd0_select_rst), .d0(selector_fused_level_2_rd0_select_d0), .d1(selector_fused_level_2_rd0_select_d1), .out(selector_fused_level_2_rd0_select_out));
  assign selector_fused_level_2_rd0_select_clk = clk;
  assign selector_fused_level_2_rd0_select_rst = rst;
  // Bindings to selector_fused_level_2_rd0_select

  // Bindings to dark_laplace_diff_2_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_laplace_diff_2_update_0_write_wdata;

  // Bindings to fused_level_2_update_0_read_rdata
    // wr_3
  assign fused_level_2_update_0_read_rdata = rd_2;



endmodule


module in_wire_dark_laplace_us_0_update_0_write_wen(output [0:0] dark_laplace_us_0_update_0_write_wen);

endmodule


module in_wire_dark_laplace_us_0_update_0_write_wdata(output [31:0] dark_laplace_us_0_update_0_write_wdata);

endmodule


module dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module dark_laplace_diff_0_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_laplace_us_1_update_0_write_wen(output [0:0] dark_laplace_us_1_update_0_write_wen);

endmodule


module dark_laplace_us_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_laplace_us_0_update_0_write_wen, input [31:0] dark_laplace_us_0_update_0_write_wdata, input [31:0] dark_laplace_diff_0_update_0_read_dummy, output [31:0] dark_laplace_diff_0_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_laplace_us_0_update_0_write_wen
    // rd_0
  assign rd_0 = dark_laplace_us_0_update_0_write_wen;

  // dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1
  logic [0:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_done;
  dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1 dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1(.clk(dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_clk), .rst(dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_rst), .start(dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_start), .done(dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_done));
  assign dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_clk = clk;
  assign dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1

  // selector_dark_laplace_diff_0_rd0_select
  logic [0:0] selector_dark_laplace_diff_0_rd0_select_clk;
  logic [0:0] selector_dark_laplace_diff_0_rd0_select_rst;
  logic [31:0] selector_dark_laplace_diff_0_rd0_select_d0;
  logic [31:0] selector_dark_laplace_diff_0_rd0_select_d1;
  logic [31:0] selector_dark_laplace_diff_0_rd0_select_out;
  dark_laplace_diff_0_rd0_select selector_dark_laplace_diff_0_rd0_select(.clk(selector_dark_laplace_diff_0_rd0_select_clk), .rst(selector_dark_laplace_diff_0_rd0_select_rst), .d0(selector_dark_laplace_diff_0_rd0_select_d0), .d1(selector_dark_laplace_diff_0_rd0_select_d1), .out(selector_dark_laplace_diff_0_rd0_select_out));
  assign selector_dark_laplace_diff_0_rd0_select_clk = clk;
  assign selector_dark_laplace_diff_0_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_diff_0_rd0_select

  // Bindings to dark_laplace_us_0_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_laplace_us_0_update_0_write_wdata;

  // Bindings to dark_laplace_diff_0_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_laplace_diff_0_update_0_read_dummy;

  // Bindings to dark_laplace_diff_0_update_0_read_rdata
    // wr_3
  assign dark_laplace_diff_0_update_0_read_rdata = rd_2;



endmodule


module dark_laplace_diff_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_laplace_us_1_update_0_write_wdata(output [31:0] dark_laplace_us_1_update_0_write_wdata);

endmodule


module dark_laplace_us_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_laplace_us_1_update_0_write_wen, input [31:0] dark_laplace_us_1_update_0_write_wdata, input [31:0] dark_laplace_diff_1_update_0_read_dummy, output [31:0] dark_laplace_diff_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_laplace_us_1_update_0_write_wen
    // rd_0
  assign rd_0 = dark_laplace_us_1_update_0_write_wen;

  // dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1
  logic [0:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_done;
  dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1 dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1(.clk(dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_clk), .rst(dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_rst), .start(dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_start), .done(dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_done));
  assign dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_clk = clk;
  assign dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1

  // selector_dark_laplace_diff_1_rd0_select
  logic [0:0] selector_dark_laplace_diff_1_rd0_select_clk;
  logic [0:0] selector_dark_laplace_diff_1_rd0_select_rst;
  logic [31:0] selector_dark_laplace_diff_1_rd0_select_d0;
  logic [31:0] selector_dark_laplace_diff_1_rd0_select_d1;
  logic [31:0] selector_dark_laplace_diff_1_rd0_select_out;
  dark_laplace_diff_1_rd0_select selector_dark_laplace_diff_1_rd0_select(.clk(selector_dark_laplace_diff_1_rd0_select_clk), .rst(selector_dark_laplace_diff_1_rd0_select_rst), .d0(selector_dark_laplace_diff_1_rd0_select_d0), .d1(selector_dark_laplace_diff_1_rd0_select_d1), .out(selector_dark_laplace_diff_1_rd0_select_out));
  assign selector_dark_laplace_diff_1_rd0_select_clk = clk;
  assign selector_dark_laplace_diff_1_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_diff_1_rd0_select

  // Bindings to dark_laplace_us_1_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_laplace_us_1_update_0_write_wdata;

  // Bindings to dark_laplace_diff_1_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_laplace_diff_1_update_0_read_dummy;

  // Bindings to dark_laplace_diff_1_update_0_read_rdata
    // wr_3
  assign dark_laplace_diff_1_update_0_read_rdata = rd_2;



endmodule


module in_wire_dark_laplace_us_2_update_0_write_wdata(output [31:0] dark_laplace_us_2_update_0_write_wdata);

endmodule


module dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_laplace_us_2_update_0_write_wen(output [0:0] dark_laplace_us_2_update_0_write_wen);

endmodule


module dark_laplace_diff_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_weights_update_0_write_wen(output [0:0] dark_weights_update_0_write_wen);

endmodule


module dark_weights_dark_weights_update_0_write0_merged_banks_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module dark_laplace_us_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_laplace_us_2_update_0_write_wen, input [31:0] dark_laplace_us_2_update_0_write_wdata, input [31:0] dark_laplace_diff_2_update_0_read_dummy, output [31:0] dark_laplace_diff_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_laplace_us_2_update_0_write_wen
    // rd_0
  assign rd_0 = dark_laplace_us_2_update_0_write_wen;

  // dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1
  logic [0:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_done;
  dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1 dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1(.clk(dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_clk), .rst(dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_rst), .start(dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_start), .done(dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_done));
  assign dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_clk = clk;
  assign dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1

  // selector_dark_laplace_diff_2_rd0_select
  logic [0:0] selector_dark_laplace_diff_2_rd0_select_clk;
  logic [0:0] selector_dark_laplace_diff_2_rd0_select_rst;
  logic [31:0] selector_dark_laplace_diff_2_rd0_select_d0;
  logic [31:0] selector_dark_laplace_diff_2_rd0_select_d1;
  logic [31:0] selector_dark_laplace_diff_2_rd0_select_out;
  dark_laplace_diff_2_rd0_select selector_dark_laplace_diff_2_rd0_select(.clk(selector_dark_laplace_diff_2_rd0_select_clk), .rst(selector_dark_laplace_diff_2_rd0_select_rst), .d0(selector_dark_laplace_diff_2_rd0_select_d0), .d1(selector_dark_laplace_diff_2_rd0_select_d1), .out(selector_dark_laplace_diff_2_rd0_select_out));
  assign selector_dark_laplace_diff_2_rd0_select_clk = clk;
  assign selector_dark_laplace_diff_2_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_diff_2_rd0_select

  // Bindings to dark_laplace_us_2_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_laplace_us_2_update_0_write_wdata;

  // Bindings to dark_laplace_diff_2_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_laplace_diff_2_update_0_read_dummy;

  // Bindings to dark_laplace_diff_2_update_0_read_rdata
    // wr_3
  assign dark_laplace_diff_2_update_0_read_rdata = rd_2;



endmodule


module weight_sums_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_weights_update_0_write_wdata(output [31:0] dark_weights_update_0_write_wdata);

endmodule


module in_wire_dark_weights_normed_update_0_read_dummy(output [31:0] dark_weights_normed_update_0_read_dummy);

endmodule


module out_wire_dark_weights_normed_update_0_read_rdata(input [31:0] dark_weights_normed_update_0_read_rdata);

endmodule


module dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1231 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f314
  logic [0:0] f314_wen;
  logic [31:0] f314_wdata;
  logic [0:0] f314_clk;
  logic [0:0] f314_rst;
  logic [31:0] f314_rdata;
  sr_buffer_32_1 f314(.wen(f314_wen), .wdata(f314_wdata), .clk(f314_clk), .rst(f314_rst), .rdata(f314_rdata));
  assign f314_clk = clk;
  assign f314_rst = rst;
  // Bindings to f314

  // f316
  logic [0:0] f316_wen;
  logic [31:0] f316_wdata;
  logic [0:0] f316_clk;
  logic [0:0] f316_rst;
  logic [31:0] f316_rdata;
  sr_buffer_32_1 f316(.wen(f316_wen), .wdata(f316_wdata), .clk(f316_clk), .rst(f316_rst), .rdata(f316_rdata));
  assign f316_clk = clk;
  assign f316_rst = rst;
  // Bindings to f316

  // f318
  logic [0:0] f318_wen;
  logic [31:0] f318_wdata;
  logic [0:0] f318_clk;
  logic [0:0] f318_rst;
  logic [31:0] f318_rdata;
  sr_buffer_32_1 f318(.wen(f318_wen), .wdata(f318_wdata), .clk(f318_clk), .rst(f318_rst), .rdata(f318_rdata));
  assign f318_clk = clk;
  assign f318_rst = rst;
  // Bindings to f318

  // f320
  logic [0:0] f320_wen;
  logic [31:0] f320_wdata;
  logic [0:0] f320_clk;
  logic [0:0] f320_rst;
  logic [31:0] f320_rdata;
  sr_buffer_32_1 f320(.wen(f320_wen), .wdata(f320_wdata), .clk(f320_clk), .rst(f320_rst), .rdata(f320_rdata));
  assign f320_clk = clk;
  assign f320_rst = rst;
  // Bindings to f320

  // f322
  logic [0:0] f322_wen;
  logic [31:0] f322_wdata;
  logic [0:0] f322_clk;
  logic [0:0] f322_rst;
  logic [31:0] f322_rdata;
  sr_buffer_32_1 f322(.wen(f322_wen), .wdata(f322_wdata), .clk(f322_clk), .rst(f322_rst), .rdata(f322_rdata));
  assign f322_clk = clk;
  assign f322_rst = rst;
  // Bindings to f322

  // f324
  logic [0:0] f324_wen;
  logic [31:0] f324_wdata;
  logic [0:0] f324_clk;
  logic [0:0] f324_rst;
  logic [31:0] f324_rdata;
  sr_buffer_32_1 f324(.wen(f324_wen), .wdata(f324_wdata), .clk(f324_clk), .rst(f324_rst), .rdata(f324_rdata));
  assign f324_clk = clk;
  assign f324_rst = rst;
  // Bindings to f324

  // f326
  logic [0:0] f326_wen;
  logic [31:0] f326_wdata;
  logic [0:0] f326_clk;
  logic [0:0] f326_rst;
  logic [31:0] f326_rdata;
  sr_buffer_32_1 f326(.wen(f326_wen), .wdata(f326_wdata), .clk(f326_clk), .rst(f326_rst), .rdata(f326_rdata));
  assign f326_clk = clk;
  assign f326_rst = rst;
  // Bindings to f326

  // f328
  logic [0:0] f328_wen;
  logic [31:0] f328_wdata;
  logic [0:0] f328_clk;
  logic [0:0] f328_rst;
  logic [31:0] f328_rdata;
  sr_buffer_32_1 f328(.wen(f328_wen), .wdata(f328_wdata), .clk(f328_clk), .rst(f328_rst), .rdata(f328_rdata));
  assign f328_clk = clk;
  assign f328_rst = rst;
  // Bindings to f328

  // f330
  logic [0:0] f330_wen;
  logic [31:0] f330_wdata;
  logic [0:0] f330_clk;
  logic [0:0] f330_rst;
  logic [31:0] f330_rdata;
  sr_buffer_32_1 f330(.wen(f330_wen), .wdata(f330_wdata), .clk(f330_clk), .rst(f330_rst), .rdata(f330_rdata));
  assign f330_clk = clk;
  assign f330_rst = rst;
  // Bindings to f330

  // f332
  logic [0:0] f332_wen;
  logic [31:0] f332_wdata;
  logic [0:0] f332_clk;
  logic [0:0] f332_rst;
  logic [31:0] f332_rdata;
  sr_buffer_32_1 f332(.wen(f332_wen), .wdata(f332_wdata), .clk(f332_clk), .rst(f332_rst), .rdata(f332_rdata));
  assign f332_clk = clk;
  assign f332_rst = rst;
  // Bindings to f332

  // f334
  logic [0:0] f334_wen;
  logic [31:0] f334_wdata;
  logic [0:0] f334_clk;
  logic [0:0] f334_rst;
  logic [31:0] f334_rdata;
  sr_buffer_32_1 f334(.wen(f334_wen), .wdata(f334_wdata), .clk(f334_clk), .rst(f334_rst), .rdata(f334_rdata));
  assign f334_clk = clk;
  assign f334_rst = rst;
  // Bindings to f334

  // f336
  logic [0:0] f336_wen;
  logic [31:0] f336_wdata;
  logic [0:0] f336_clk;
  logic [0:0] f336_rst;
  logic [31:0] f336_rdata;
  sr_buffer_32_1 f336(.wen(f336_wen), .wdata(f336_wdata), .clk(f336_clk), .rst(f336_rst), .rdata(f336_rdata));
  assign f336_clk = clk;
  assign f336_rst = rst;
  // Bindings to f336

  // f338
  logic [0:0] f338_wen;
  logic [31:0] f338_wdata;
  logic [0:0] f338_clk;
  logic [0:0] f338_rst;
  logic [31:0] f338_rdata;
  sr_buffer_32_1 f338(.wen(f338_wen), .wdata(f338_wdata), .clk(f338_clk), .rst(f338_rst), .rdata(f338_rdata));
  assign f338_clk = clk;
  assign f338_rst = rst;
  // Bindings to f338

  // f340
  logic [0:0] f340_wen;
  logic [31:0] f340_wdata;
  logic [0:0] f340_clk;
  logic [0:0] f340_rst;
  logic [31:0] f340_rdata;
  sr_buffer_32_1 f340(.wen(f340_wen), .wdata(f340_wdata), .clk(f340_clk), .rst(f340_rst), .rdata(f340_rdata));
  assign f340_clk = clk;
  assign f340_rst = rst;
  // Bindings to f340

  // f342
  logic [0:0] f342_wen;
  logic [31:0] f342_wdata;
  logic [0:0] f342_clk;
  logic [0:0] f342_rst;
  logic [31:0] f342_rdata;
  sr_buffer_32_1 f342(.wen(f342_wen), .wdata(f342_wdata), .clk(f342_clk), .rst(f342_rst), .rdata(f342_rdata));
  assign f342_clk = clk;
  assign f342_rst = rst;
  // Bindings to f342

  // f344
  logic [0:0] f344_wen;
  logic [31:0] f344_wdata;
  logic [0:0] f344_clk;
  logic [0:0] f344_rst;
  logic [31:0] f344_rdata;
  sr_buffer_32_1 f344(.wen(f344_wen), .wdata(f344_wdata), .clk(f344_clk), .rst(f344_rst), .rdata(f344_rdata));
  assign f344_clk = clk;
  assign f344_rst = rst;
  // Bindings to f344

  // f346
  logic [0:0] f346_wen;
  logic [31:0] f346_wdata;
  logic [0:0] f346_clk;
  logic [0:0] f346_rst;
  logic [31:0] f346_rdata;
  sr_buffer_32_1 f346(.wen(f346_wen), .wdata(f346_wdata), .clk(f346_clk), .rst(f346_rst), .rdata(f346_rdata));
  assign f346_clk = clk;
  assign f346_rst = rst;
  // Bindings to f346

  // f348
  logic [0:0] f348_wen;
  logic [31:0] f348_wdata;
  logic [0:0] f348_clk;
  logic [0:0] f348_rst;
  logic [31:0] f348_rdata;
  sr_buffer_32_1 f348(.wen(f348_wen), .wdata(f348_wdata), .clk(f348_clk), .rst(f348_rst), .rdata(f348_rdata));
  assign f348_clk = clk;
  assign f348_rst = rst;
  // Bindings to f348

  // f350
  logic [0:0] f350_wen;
  logic [31:0] f350_wdata;
  logic [0:0] f350_clk;
  logic [0:0] f350_rst;
  logic [31:0] f350_rdata;
  sr_buffer_32_1 f350(.wen(f350_wen), .wdata(f350_wdata), .clk(f350_clk), .rst(f350_rst), .rdata(f350_rdata));
  assign f350_clk = clk;
  assign f350_rst = rst;
  // Bindings to f350

  // f352
  logic [0:0] f352_wen;
  logic [31:0] f352_wdata;
  logic [0:0] f352_clk;
  logic [0:0] f352_rst;
  logic [31:0] f352_rdata;
  sr_buffer_32_1 f352(.wen(f352_wen), .wdata(f352_wdata), .clk(f352_clk), .rst(f352_rst), .rdata(f352_rdata));
  assign f352_clk = clk;
  assign f352_rst = rst;
  // Bindings to f352

  // f354
  logic [0:0] f354_wen;
  logic [31:0] f354_wdata;
  logic [0:0] f354_clk;
  logic [0:0] f354_rst;
  logic [31:0] f354_rdata;
  sr_buffer_32_1 f354(.wen(f354_wen), .wdata(f354_wdata), .clk(f354_clk), .rst(f354_rst), .rdata(f354_rdata));
  assign f354_clk = clk;
  assign f354_rst = rst;
  // Bindings to f354

  // f356
  logic [0:0] f356_wen;
  logic [31:0] f356_wdata;
  logic [0:0] f356_clk;
  logic [0:0] f356_rst;
  logic [31:0] f356_rdata;
  sr_buffer_32_1 f356(.wen(f356_wen), .wdata(f356_wdata), .clk(f356_clk), .rst(f356_rst), .rdata(f356_rdata));
  assign f356_clk = clk;
  assign f356_rst = rst;
  // Bindings to f356

  // f358
  logic [0:0] f358_wen;
  logic [31:0] f358_wdata;
  logic [0:0] f358_clk;
  logic [0:0] f358_rst;
  logic [31:0] f358_rdata;
  sr_buffer_32_1 f358(.wen(f358_wen), .wdata(f358_wdata), .clk(f358_clk), .rst(f358_rst), .rdata(f358_rdata));
  assign f358_clk = clk;
  assign f358_rst = rst;
  // Bindings to f358

  // f360
  logic [0:0] f360_wen;
  logic [31:0] f360_wdata;
  logic [0:0] f360_clk;
  logic [0:0] f360_rst;
  logic [31:0] f360_rdata;
  sr_buffer_32_1 f360(.wen(f360_wen), .wdata(f360_wdata), .clk(f360_clk), .rst(f360_rst), .rdata(f360_rdata));
  assign f360_clk = clk;
  assign f360_rst = rst;
  // Bindings to f360

  // f362
  logic [0:0] f362_wen;
  logic [31:0] f362_wdata;
  logic [0:0] f362_clk;
  logic [0:0] f362_rst;
  logic [31:0] f362_rdata;
  sr_buffer_32_1 f362(.wen(f362_wen), .wdata(f362_wdata), .clk(f362_clk), .rst(f362_rst), .rdata(f362_rdata));
  assign f362_clk = clk;
  assign f362_rst = rst;
  // Bindings to f362

  // f364
  logic [0:0] f364_wen;
  logic [31:0] f364_wdata;
  logic [0:0] f364_clk;
  logic [0:0] f364_rst;
  logic [31:0] f364_rdata;
  sr_buffer_32_1 f364(.wen(f364_wen), .wdata(f364_wdata), .clk(f364_clk), .rst(f364_rst), .rdata(f364_rdata));
  assign f364_clk = clk;
  assign f364_rst = rst;
  // Bindings to f364

  // f366
  logic [0:0] f366_wen;
  logic [31:0] f366_wdata;
  logic [0:0] f366_clk;
  logic [0:0] f366_rst;
  logic [31:0] f366_rdata;
  sr_buffer_32_1 f366(.wen(f366_wen), .wdata(f366_wdata), .clk(f366_clk), .rst(f366_rst), .rdata(f366_rdata));
  assign f366_clk = clk;
  assign f366_rst = rst;
  // Bindings to f366

  // f368
  logic [0:0] f368_wen;
  logic [31:0] f368_wdata;
  logic [0:0] f368_clk;
  logic [0:0] f368_rst;
  logic [31:0] f368_rdata;
  sr_buffer_32_1 f368(.wen(f368_wen), .wdata(f368_wdata), .clk(f368_clk), .rst(f368_rst), .rdata(f368_rdata));
  assign f368_clk = clk;
  assign f368_rst = rst;
  // Bindings to f368

  // f370
  logic [0:0] f370_wen;
  logic [31:0] f370_wdata;
  logic [0:0] f370_clk;
  logic [0:0] f370_rst;
  logic [31:0] f370_rdata;
  sr_buffer_32_1 f370(.wen(f370_wen), .wdata(f370_wdata), .clk(f370_clk), .rst(f370_rst), .rdata(f370_rdata));
  assign f370_clk = clk;
  assign f370_rst = rst;
  // Bindings to f370

  // f372
  logic [0:0] f372_wen;
  logic [31:0] f372_wdata;
  logic [0:0] f372_clk;
  logic [0:0] f372_rst;
  logic [31:0] f372_rdata;
  sr_buffer_32_1 f372(.wen(f372_wen), .wdata(f372_wdata), .clk(f372_clk), .rst(f372_rst), .rdata(f372_rdata));
  assign f372_clk = clk;
  assign f372_rst = rst;
  // Bindings to f372

  // f374
  logic [0:0] f374_wen;
  logic [31:0] f374_wdata;
  logic [0:0] f374_clk;
  logic [0:0] f374_rst;
  logic [31:0] f374_rdata;
  sr_buffer_32_1 f374(.wen(f374_wen), .wdata(f374_wdata), .clk(f374_clk), .rst(f374_rst), .rdata(f374_rdata));
  assign f374_clk = clk;
  assign f374_rst = rst;
  // Bindings to f374

  // f376
  logic [0:0] f376_wen;
  logic [31:0] f376_wdata;
  logic [0:0] f376_clk;
  logic [0:0] f376_rst;
  logic [31:0] f376_rdata;
  sr_buffer_32_1 f376(.wen(f376_wen), .wdata(f376_wdata), .clk(f376_clk), .rst(f376_rst), .rdata(f376_rdata));
  assign f376_clk = clk;
  assign f376_rst = rst;
  // Bindings to f376

  // f378
  logic [0:0] f378_wen;
  logic [31:0] f378_wdata;
  logic [0:0] f378_clk;
  logic [0:0] f378_rst;
  logic [31:0] f378_rdata;
  sr_buffer_32_1 f378(.wen(f378_wen), .wdata(f378_wdata), .clk(f378_clk), .rst(f378_rst), .rdata(f378_rdata));
  assign f378_clk = clk;
  assign f378_rst = rst;
  // Bindings to f378

  // f380
  logic [0:0] f380_wen;
  logic [31:0] f380_wdata;
  logic [0:0] f380_clk;
  logic [0:0] f380_rst;
  logic [31:0] f380_rdata;
  sr_buffer_32_1 f380(.wen(f380_wen), .wdata(f380_wdata), .clk(f380_clk), .rst(f380_rst), .rdata(f380_rdata));
  assign f380_clk = clk;
  assign f380_rst = rst;
  // Bindings to f380

  // f382
  logic [0:0] f382_wen;
  logic [31:0] f382_wdata;
  logic [0:0] f382_clk;
  logic [0:0] f382_rst;
  logic [31:0] f382_rdata;
  sr_buffer_32_1 f382(.wen(f382_wen), .wdata(f382_wdata), .clk(f382_clk), .rst(f382_rst), .rdata(f382_rdata));
  assign f382_clk = clk;
  assign f382_rst = rst;
  // Bindings to f382

  // f384
  logic [0:0] f384_wen;
  logic [31:0] f384_wdata;
  logic [0:0] f384_clk;
  logic [0:0] f384_rst;
  logic [31:0] f384_rdata;
  sr_buffer_32_1 f384(.wen(f384_wen), .wdata(f384_wdata), .clk(f384_clk), .rst(f384_rst), .rdata(f384_rdata));
  assign f384_clk = clk;
  assign f384_rst = rst;
  // Bindings to f384

  // f386
  logic [0:0] f386_wen;
  logic [31:0] f386_wdata;
  logic [0:0] f386_clk;
  logic [0:0] f386_rst;
  logic [31:0] f386_rdata;
  sr_buffer_32_1 f386(.wen(f386_wen), .wdata(f386_wdata), .clk(f386_clk), .rst(f386_rst), .rdata(f386_rdata));
  assign f386_clk = clk;
  assign f386_rst = rst;
  // Bindings to f386

  // f388
  logic [0:0] f388_wen;
  logic [31:0] f388_wdata;
  logic [0:0] f388_clk;
  logic [0:0] f388_rst;
  logic [31:0] f388_rdata;
  sr_buffer_32_1 f388(.wen(f388_wen), .wdata(f388_wdata), .clk(f388_clk), .rst(f388_rst), .rdata(f388_rdata));
  assign f388_clk = clk;
  assign f388_rst = rst;
  // Bindings to f388

  // f390
  logic [0:0] f390_wen;
  logic [31:0] f390_wdata;
  logic [0:0] f390_clk;
  logic [0:0] f390_rst;
  logic [31:0] f390_rdata;
  sr_buffer_32_1 f390(.wen(f390_wen), .wdata(f390_wdata), .clk(f390_clk), .rst(f390_rst), .rdata(f390_rdata));
  assign f390_clk = clk;
  assign f390_rst = rst;
  // Bindings to f390

  // f392
  logic [0:0] f392_wen;
  logic [31:0] f392_wdata;
  logic [0:0] f392_clk;
  logic [0:0] f392_rst;
  logic [31:0] f392_rdata;
  sr_buffer_32_1 f392(.wen(f392_wen), .wdata(f392_wdata), .clk(f392_clk), .rst(f392_rst), .rdata(f392_rdata));
  assign f392_clk = clk;
  assign f392_rst = rst;
  // Bindings to f392

  // f394
  logic [0:0] f394_wen;
  logic [31:0] f394_wdata;
  logic [0:0] f394_clk;
  logic [0:0] f394_rst;
  logic [31:0] f394_rdata;
  sr_buffer_32_1 f394(.wen(f394_wen), .wdata(f394_wdata), .clk(f394_clk), .rst(f394_rst), .rdata(f394_rdata));
  assign f394_clk = clk;
  assign f394_rst = rst;
  // Bindings to f394

  // f396
  logic [0:0] f396_wen;
  logic [31:0] f396_wdata;
  logic [0:0] f396_clk;
  logic [0:0] f396_rst;
  logic [31:0] f396_rdata;
  sr_buffer_32_1 f396(.wen(f396_wen), .wdata(f396_wdata), .clk(f396_clk), .rst(f396_rst), .rdata(f396_rdata));
  assign f396_clk = clk;
  assign f396_rst = rst;
  // Bindings to f396

  // f398
  logic [0:0] f398_wen;
  logic [31:0] f398_wdata;
  logic [0:0] f398_clk;
  logic [0:0] f398_rst;
  logic [31:0] f398_rdata;
  sr_buffer_32_1 f398(.wen(f398_wen), .wdata(f398_wdata), .clk(f398_clk), .rst(f398_rst), .rdata(f398_rdata));
  assign f398_clk = clk;
  assign f398_rst = rst;
  // Bindings to f398

  // f400
  logic [0:0] f400_wen;
  logic [31:0] f400_wdata;
  logic [0:0] f400_clk;
  logic [0:0] f400_rst;
  logic [31:0] f400_rdata;
  sr_buffer_32_1 f400(.wen(f400_wen), .wdata(f400_wdata), .clk(f400_clk), .rst(f400_rst), .rdata(f400_rdata));
  assign f400_clk = clk;
  assign f400_rst = rst;
  // Bindings to f400

  // f402
  logic [0:0] f402_wen;
  logic [31:0] f402_wdata;
  logic [0:0] f402_clk;
  logic [0:0] f402_rst;
  logic [31:0] f402_rdata;
  sr_buffer_32_1 f402(.wen(f402_wen), .wdata(f402_wdata), .clk(f402_clk), .rst(f402_rst), .rdata(f402_rdata));
  assign f402_clk = clk;
  assign f402_rst = rst;
  // Bindings to f402

  // f404
  logic [0:0] f404_wen;
  logic [31:0] f404_wdata;
  logic [0:0] f404_clk;
  logic [0:0] f404_rst;
  logic [31:0] f404_rdata;
  sr_buffer_32_1 f404(.wen(f404_wen), .wdata(f404_wdata), .clk(f404_clk), .rst(f404_rst), .rdata(f404_rdata));
  assign f404_clk = clk;
  assign f404_rst = rst;
  // Bindings to f404

  // f406
  logic [0:0] f406_wen;
  logic [31:0] f406_wdata;
  logic [0:0] f406_clk;
  logic [0:0] f406_rst;
  logic [31:0] f406_rdata;
  sr_buffer_32_1 f406(.wen(f406_wen), .wdata(f406_wdata), .clk(f406_clk), .rst(f406_rst), .rdata(f406_rdata));
  assign f406_clk = clk;
  assign f406_rst = rst;
  // Bindings to f406

  // f408
  logic [0:0] f408_wen;
  logic [31:0] f408_wdata;
  logic [0:0] f408_clk;
  logic [0:0] f408_rst;
  logic [31:0] f408_rdata;
  sr_buffer_32_1 f408(.wen(f408_wen), .wdata(f408_wdata), .clk(f408_clk), .rst(f408_rst), .rdata(f408_rdata));
  assign f408_clk = clk;
  assign f408_rst = rst;
  // Bindings to f408

  // f410
  logic [0:0] f410_wen;
  logic [31:0] f410_wdata;
  logic [0:0] f410_clk;
  logic [0:0] f410_rst;
  logic [31:0] f410_rdata;
  sr_buffer_32_1 f410(.wen(f410_wen), .wdata(f410_wdata), .clk(f410_clk), .rst(f410_rst), .rdata(f410_rdata));
  assign f410_clk = clk;
  assign f410_rst = rst;
  // Bindings to f410

  // f412
  logic [0:0] f412_wen;
  logic [31:0] f412_wdata;
  logic [0:0] f412_clk;
  logic [0:0] f412_rst;
  logic [31:0] f412_rdata;
  sr_buffer_32_1 f412(.wen(f412_wen), .wdata(f412_wdata), .clk(f412_clk), .rst(f412_rst), .rdata(f412_rdata));
  assign f412_clk = clk;
  assign f412_rst = rst;
  // Bindings to f412

  // f414
  logic [0:0] f414_wen;
  logic [31:0] f414_wdata;
  logic [0:0] f414_clk;
  logic [0:0] f414_rst;
  logic [31:0] f414_rdata;
  sr_buffer_32_1 f414(.wen(f414_wen), .wdata(f414_wdata), .clk(f414_clk), .rst(f414_rst), .rdata(f414_rdata));
  assign f414_clk = clk;
  assign f414_rst = rst;
  // Bindings to f414

  // f416
  logic [0:0] f416_wen;
  logic [31:0] f416_wdata;
  logic [0:0] f416_clk;
  logic [0:0] f416_rst;
  logic [31:0] f416_rdata;
  sr_buffer_32_1 f416(.wen(f416_wen), .wdata(f416_wdata), .clk(f416_clk), .rst(f416_rst), .rdata(f416_rdata));
  assign f416_clk = clk;
  assign f416_rst = rst;
  // Bindings to f416

  // f418
  logic [0:0] f418_wen;
  logic [31:0] f418_wdata;
  logic [0:0] f418_clk;
  logic [0:0] f418_rst;
  logic [31:0] f418_rdata;
  sr_buffer_32_1 f418(.wen(f418_wen), .wdata(f418_wdata), .clk(f418_clk), .rst(f418_rst), .rdata(f418_rdata));
  assign f418_clk = clk;
  assign f418_rst = rst;
  // Bindings to f418

  // f420
  logic [0:0] f420_wen;
  logic [31:0] f420_wdata;
  logic [0:0] f420_clk;
  logic [0:0] f420_rst;
  logic [31:0] f420_rdata;
  sr_buffer_32_1 f420(.wen(f420_wen), .wdata(f420_wdata), .clk(f420_clk), .rst(f420_rst), .rdata(f420_rdata));
  assign f420_clk = clk;
  assign f420_rst = rst;
  // Bindings to f420

  // f422
  logic [0:0] f422_wen;
  logic [31:0] f422_wdata;
  logic [0:0] f422_clk;
  logic [0:0] f422_rst;
  logic [31:0] f422_rdata;
  sr_buffer_32_1 f422(.wen(f422_wen), .wdata(f422_wdata), .clk(f422_clk), .rst(f422_rst), .rdata(f422_rdata));
  assign f422_clk = clk;
  assign f422_rst = rst;
  // Bindings to f422

  // f424
  logic [0:0] f424_wen;
  logic [31:0] f424_wdata;
  logic [0:0] f424_clk;
  logic [0:0] f424_rst;
  logic [31:0] f424_rdata;
  sr_buffer_32_1 f424(.wen(f424_wen), .wdata(f424_wdata), .clk(f424_clk), .rst(f424_rst), .rdata(f424_rdata));
  assign f424_clk = clk;
  assign f424_rst = rst;
  // Bindings to f424

  // f426
  logic [0:0] f426_wen;
  logic [31:0] f426_wdata;
  logic [0:0] f426_clk;
  logic [0:0] f426_rst;
  logic [31:0] f426_rdata;
  sr_buffer_32_1 f426(.wen(f426_wen), .wdata(f426_wdata), .clk(f426_clk), .rst(f426_rst), .rdata(f426_rdata));
  assign f426_clk = clk;
  assign f426_rst = rst;
  // Bindings to f426

  // f428
  logic [0:0] f428_wen;
  logic [31:0] f428_wdata;
  logic [0:0] f428_clk;
  logic [0:0] f428_rst;
  logic [31:0] f428_rdata;
  sr_buffer_32_1 f428(.wen(f428_wen), .wdata(f428_wdata), .clk(f428_clk), .rst(f428_rst), .rdata(f428_rdata));
  assign f428_clk = clk;
  assign f428_rst = rst;
  // Bindings to f428

  // f430
  logic [0:0] f430_wen;
  logic [31:0] f430_wdata;
  logic [0:0] f430_clk;
  logic [0:0] f430_rst;
  logic [31:0] f430_rdata;
  sr_buffer_32_1 f430(.wen(f430_wen), .wdata(f430_wdata), .clk(f430_clk), .rst(f430_rst), .rdata(f430_rdata));
  assign f430_clk = clk;
  assign f430_rst = rst;
  // Bindings to f430

  // f432
  logic [0:0] f432_wen;
  logic [31:0] f432_wdata;
  logic [0:0] f432_clk;
  logic [0:0] f432_rst;
  logic [31:0] f432_rdata;
  sr_buffer_32_1 f432(.wen(f432_wen), .wdata(f432_wdata), .clk(f432_clk), .rst(f432_rst), .rdata(f432_rdata));
  assign f432_clk = clk;
  assign f432_rst = rst;
  // Bindings to f432

  // f434
  logic [0:0] f434_wen;
  logic [31:0] f434_wdata;
  logic [0:0] f434_clk;
  logic [0:0] f434_rst;
  logic [31:0] f434_rdata;
  sr_buffer_32_1 f434(.wen(f434_wen), .wdata(f434_wdata), .clk(f434_clk), .rst(f434_rst), .rdata(f434_rdata));
  assign f434_clk = clk;
  assign f434_rst = rst;
  // Bindings to f434

  // f436
  logic [0:0] f436_wen;
  logic [31:0] f436_wdata;
  logic [0:0] f436_clk;
  logic [0:0] f436_rst;
  logic [31:0] f436_rdata;
  sr_buffer_32_1 f436(.wen(f436_wen), .wdata(f436_wdata), .clk(f436_clk), .rst(f436_rst), .rdata(f436_rdata));
  assign f436_clk = clk;
  assign f436_rst = rst;
  // Bindings to f436

  // f438
  logic [0:0] f438_wen;
  logic [31:0] f438_wdata;
  logic [0:0] f438_clk;
  logic [0:0] f438_rst;
  logic [31:0] f438_rdata;
  sr_buffer_32_1 f438(.wen(f438_wen), .wdata(f438_wdata), .clk(f438_clk), .rst(f438_rst), .rdata(f438_rdata));
  assign f438_clk = clk;
  assign f438_rst = rst;
  // Bindings to f438

  // f440
  logic [0:0] f440_wen;
  logic [31:0] f440_wdata;
  logic [0:0] f440_clk;
  logic [0:0] f440_rst;
  logic [31:0] f440_rdata;
  sr_buffer_32_1 f440(.wen(f440_wen), .wdata(f440_wdata), .clk(f440_clk), .rst(f440_rst), .rdata(f440_rdata));
  assign f440_clk = clk;
  assign f440_rst = rst;
  // Bindings to f440

  // f442
  logic [0:0] f442_wen;
  logic [31:0] f442_wdata;
  logic [0:0] f442_clk;
  logic [0:0] f442_rst;
  logic [31:0] f442_rdata;
  sr_buffer_32_1 f442(.wen(f442_wen), .wdata(f442_wdata), .clk(f442_clk), .rst(f442_rst), .rdata(f442_rdata));
  assign f442_clk = clk;
  assign f442_rst = rst;
  // Bindings to f442

  // f444
  logic [0:0] f444_wen;
  logic [31:0] f444_wdata;
  logic [0:0] f444_clk;
  logic [0:0] f444_rst;
  logic [31:0] f444_rdata;
  sr_buffer_32_1 f444(.wen(f444_wen), .wdata(f444_wdata), .clk(f444_clk), .rst(f444_rst), .rdata(f444_rdata));
  assign f444_clk = clk;
  assign f444_rst = rst;
  // Bindings to f444

  // f446
  logic [0:0] f446_wen;
  logic [31:0] f446_wdata;
  logic [0:0] f446_clk;
  logic [0:0] f446_rst;
  logic [31:0] f446_rdata;
  sr_buffer_32_1 f446(.wen(f446_wen), .wdata(f446_wdata), .clk(f446_clk), .rst(f446_rst), .rdata(f446_rdata));
  assign f446_clk = clk;
  assign f446_rst = rst;
  // Bindings to f446

  // f448
  logic [0:0] f448_wen;
  logic [31:0] f448_wdata;
  logic [0:0] f448_clk;
  logic [0:0] f448_rst;
  logic [31:0] f448_rdata;
  sr_buffer_32_1 f448(.wen(f448_wen), .wdata(f448_wdata), .clk(f448_clk), .rst(f448_rst), .rdata(f448_rdata));
  assign f448_clk = clk;
  assign f448_rst = rst;
  // Bindings to f448

  // f450
  logic [0:0] f450_wen;
  logic [31:0] f450_wdata;
  logic [0:0] f450_clk;
  logic [0:0] f450_rst;
  logic [31:0] f450_rdata;
  sr_buffer_32_1 f450(.wen(f450_wen), .wdata(f450_wdata), .clk(f450_clk), .rst(f450_rst), .rdata(f450_rdata));
  assign f450_clk = clk;
  assign f450_rst = rst;
  // Bindings to f450

  // f452
  logic [0:0] f452_wen;
  logic [31:0] f452_wdata;
  logic [0:0] f452_clk;
  logic [0:0] f452_rst;
  logic [31:0] f452_rdata;
  sr_buffer_32_1 f452(.wen(f452_wen), .wdata(f452_wdata), .clk(f452_clk), .rst(f452_rst), .rdata(f452_rdata));
  assign f452_clk = clk;
  assign f452_rst = rst;
  // Bindings to f452

  // f454
  logic [0:0] f454_wen;
  logic [31:0] f454_wdata;
  logic [0:0] f454_clk;
  logic [0:0] f454_rst;
  logic [31:0] f454_rdata;
  sr_buffer_32_1 f454(.wen(f454_wen), .wdata(f454_wdata), .clk(f454_clk), .rst(f454_rst), .rdata(f454_rdata));
  assign f454_clk = clk;
  assign f454_rst = rst;
  // Bindings to f454

  // f456
  logic [0:0] f456_wen;
  logic [31:0] f456_wdata;
  logic [0:0] f456_clk;
  logic [0:0] f456_rst;
  logic [31:0] f456_rdata;
  sr_buffer_32_1 f456(.wen(f456_wen), .wdata(f456_wdata), .clk(f456_clk), .rst(f456_rst), .rdata(f456_rdata));
  assign f456_clk = clk;
  assign f456_rst = rst;
  // Bindings to f456

  // f458
  logic [0:0] f458_wen;
  logic [31:0] f458_wdata;
  logic [0:0] f458_clk;
  logic [0:0] f458_rst;
  logic [31:0] f458_rdata;
  sr_buffer_32_1 f458(.wen(f458_wen), .wdata(f458_wdata), .clk(f458_clk), .rst(f458_rst), .rdata(f458_rdata));
  assign f458_clk = clk;
  assign f458_rst = rst;
  // Bindings to f458

  // f460
  logic [0:0] f460_wen;
  logic [31:0] f460_wdata;
  logic [0:0] f460_clk;
  logic [0:0] f460_rst;
  logic [31:0] f460_rdata;
  sr_buffer_32_1 f460(.wen(f460_wen), .wdata(f460_wdata), .clk(f460_clk), .rst(f460_rst), .rdata(f460_rdata));
  assign f460_clk = clk;
  assign f460_rst = rst;
  // Bindings to f460

  // f462
  logic [0:0] f462_wen;
  logic [31:0] f462_wdata;
  logic [0:0] f462_clk;
  logic [0:0] f462_rst;
  logic [31:0] f462_rdata;
  sr_buffer_32_1 f462(.wen(f462_wen), .wdata(f462_wdata), .clk(f462_clk), .rst(f462_rst), .rdata(f462_rdata));
  assign f462_clk = clk;
  assign f462_rst = rst;
  // Bindings to f462

  // f464
  logic [0:0] f464_wen;
  logic [31:0] f464_wdata;
  logic [0:0] f464_clk;
  logic [0:0] f464_rst;
  logic [31:0] f464_rdata;
  sr_buffer_32_1 f464(.wen(f464_wen), .wdata(f464_wdata), .clk(f464_clk), .rst(f464_rst), .rdata(f464_rdata));
  assign f464_clk = clk;
  assign f464_rst = rst;
  // Bindings to f464

  // f466
  logic [0:0] f466_wen;
  logic [31:0] f466_wdata;
  logic [0:0] f466_clk;
  logic [0:0] f466_rst;
  logic [31:0] f466_rdata;
  sr_buffer_32_1 f466(.wen(f466_wen), .wdata(f466_wdata), .clk(f466_clk), .rst(f466_rst), .rdata(f466_rdata));
  assign f466_clk = clk;
  assign f466_rst = rst;
  // Bindings to f466

  // f468
  logic [0:0] f468_wen;
  logic [31:0] f468_wdata;
  logic [0:0] f468_clk;
  logic [0:0] f468_rst;
  logic [31:0] f468_rdata;
  sr_buffer_32_1 f468(.wen(f468_wen), .wdata(f468_wdata), .clk(f468_clk), .rst(f468_rst), .rdata(f468_rdata));
  assign f468_clk = clk;
  assign f468_rst = rst;
  // Bindings to f468

  // f470
  logic [0:0] f470_wen;
  logic [31:0] f470_wdata;
  logic [0:0] f470_clk;
  logic [0:0] f470_rst;
  logic [31:0] f470_rdata;
  sr_buffer_32_1 f470(.wen(f470_wen), .wdata(f470_wdata), .clk(f470_clk), .rst(f470_rst), .rdata(f470_rdata));
  assign f470_clk = clk;
  assign f470_rst = rst;
  // Bindings to f470

  // f472
  logic [0:0] f472_wen;
  logic [31:0] f472_wdata;
  logic [0:0] f472_clk;
  logic [0:0] f472_rst;
  logic [31:0] f472_rdata;
  sr_buffer_32_1 f472(.wen(f472_wen), .wdata(f472_wdata), .clk(f472_clk), .rst(f472_rst), .rdata(f472_rdata));
  assign f472_clk = clk;
  assign f472_rst = rst;
  // Bindings to f472

  // f474
  logic [0:0] f474_wen;
  logic [31:0] f474_wdata;
  logic [0:0] f474_clk;
  logic [0:0] f474_rst;
  logic [31:0] f474_rdata;
  sr_buffer_32_1 f474(.wen(f474_wen), .wdata(f474_wdata), .clk(f474_clk), .rst(f474_rst), .rdata(f474_rdata));
  assign f474_clk = clk;
  assign f474_rst = rst;
  // Bindings to f474

  // f476
  logic [0:0] f476_wen;
  logic [31:0] f476_wdata;
  logic [0:0] f476_clk;
  logic [0:0] f476_rst;
  logic [31:0] f476_rdata;
  sr_buffer_32_1 f476(.wen(f476_wen), .wdata(f476_wdata), .clk(f476_clk), .rst(f476_rst), .rdata(f476_rdata));
  assign f476_clk = clk;
  assign f476_rst = rst;
  // Bindings to f476

  // f478
  logic [0:0] f478_wen;
  logic [31:0] f478_wdata;
  logic [0:0] f478_clk;
  logic [0:0] f478_rst;
  logic [31:0] f478_rdata;
  sr_buffer_32_1 f478(.wen(f478_wen), .wdata(f478_wdata), .clk(f478_clk), .rst(f478_rst), .rdata(f478_rdata));
  assign f478_clk = clk;
  assign f478_rst = rst;
  // Bindings to f478

  // f480
  logic [0:0] f480_wen;
  logic [31:0] f480_wdata;
  logic [0:0] f480_clk;
  logic [0:0] f480_rst;
  logic [31:0] f480_rdata;
  sr_buffer_32_1 f480(.wen(f480_wen), .wdata(f480_wdata), .clk(f480_clk), .rst(f480_rst), .rdata(f480_rdata));
  assign f480_clk = clk;
  assign f480_rst = rst;
  // Bindings to f480

  // f482
  logic [0:0] f482_wen;
  logic [31:0] f482_wdata;
  logic [0:0] f482_clk;
  logic [0:0] f482_rst;
  logic [31:0] f482_rdata;
  sr_buffer_32_1 f482(.wen(f482_wen), .wdata(f482_wdata), .clk(f482_clk), .rst(f482_rst), .rdata(f482_rdata));
  assign f482_clk = clk;
  assign f482_rst = rst;
  // Bindings to f482

  // f484
  logic [0:0] f484_wen;
  logic [31:0] f484_wdata;
  logic [0:0] f484_clk;
  logic [0:0] f484_rst;
  logic [31:0] f484_rdata;
  sr_buffer_32_1 f484(.wen(f484_wen), .wdata(f484_wdata), .clk(f484_clk), .rst(f484_rst), .rdata(f484_rdata));
  assign f484_clk = clk;
  assign f484_rst = rst;
  // Bindings to f484

  // f486
  logic [0:0] f486_wen;
  logic [31:0] f486_wdata;
  logic [0:0] f486_clk;
  logic [0:0] f486_rst;
  logic [31:0] f486_rdata;
  sr_buffer_32_1 f486(.wen(f486_wen), .wdata(f486_wdata), .clk(f486_clk), .rst(f486_rst), .rdata(f486_rdata));
  assign f486_clk = clk;
  assign f486_rst = rst;
  // Bindings to f486

  // f488
  logic [0:0] f488_wen;
  logic [31:0] f488_wdata;
  logic [0:0] f488_clk;
  logic [0:0] f488_rst;
  logic [31:0] f488_rdata;
  sr_buffer_32_1 f488(.wen(f488_wen), .wdata(f488_wdata), .clk(f488_clk), .rst(f488_rst), .rdata(f488_rdata));
  assign f488_clk = clk;
  assign f488_rst = rst;
  // Bindings to f488

  // f490
  logic [0:0] f490_wen;
  logic [31:0] f490_wdata;
  logic [0:0] f490_clk;
  logic [0:0] f490_rst;
  logic [31:0] f490_rdata;
  sr_buffer_32_1 f490(.wen(f490_wen), .wdata(f490_wdata), .clk(f490_clk), .rst(f490_rst), .rdata(f490_rdata));
  assign f490_clk = clk;
  assign f490_rst = rst;
  // Bindings to f490

  // f492
  logic [0:0] f492_wen;
  logic [31:0] f492_wdata;
  logic [0:0] f492_clk;
  logic [0:0] f492_rst;
  logic [31:0] f492_rdata;
  sr_buffer_32_1 f492(.wen(f492_wen), .wdata(f492_wdata), .clk(f492_clk), .rst(f492_rst), .rdata(f492_rdata));
  assign f492_clk = clk;
  assign f492_rst = rst;
  // Bindings to f492

  // f494
  logic [0:0] f494_wen;
  logic [31:0] f494_wdata;
  logic [0:0] f494_clk;
  logic [0:0] f494_rst;
  logic [31:0] f494_rdata;
  sr_buffer_32_1 f494(.wen(f494_wen), .wdata(f494_wdata), .clk(f494_clk), .rst(f494_rst), .rdata(f494_rdata));
  assign f494_clk = clk;
  assign f494_rst = rst;
  // Bindings to f494

  // f496
  logic [0:0] f496_wen;
  logic [31:0] f496_wdata;
  logic [0:0] f496_clk;
  logic [0:0] f496_rst;
  logic [31:0] f496_rdata;
  sr_buffer_32_1 f496(.wen(f496_wen), .wdata(f496_wdata), .clk(f496_clk), .rst(f496_rst), .rdata(f496_rdata));
  assign f496_clk = clk;
  assign f496_rst = rst;
  // Bindings to f496

  // f498
  logic [0:0] f498_wen;
  logic [31:0] f498_wdata;
  logic [0:0] f498_clk;
  logic [0:0] f498_rst;
  logic [31:0] f498_rdata;
  sr_buffer_32_1 f498(.wen(f498_wen), .wdata(f498_wdata), .clk(f498_clk), .rst(f498_rst), .rdata(f498_rdata));
  assign f498_clk = clk;
  assign f498_rst = rst;
  // Bindings to f498

  // f500
  logic [0:0] f500_wen;
  logic [31:0] f500_wdata;
  logic [0:0] f500_clk;
  logic [0:0] f500_rst;
  logic [31:0] f500_rdata;
  sr_buffer_32_1 f500(.wen(f500_wen), .wdata(f500_wdata), .clk(f500_clk), .rst(f500_rst), .rdata(f500_rdata));
  assign f500_clk = clk;
  assign f500_rst = rst;
  // Bindings to f500

  // f502
  logic [0:0] f502_wen;
  logic [31:0] f502_wdata;
  logic [0:0] f502_clk;
  logic [0:0] f502_rst;
  logic [31:0] f502_rdata;
  sr_buffer_32_1 f502(.wen(f502_wen), .wdata(f502_wdata), .clk(f502_clk), .rst(f502_rst), .rdata(f502_rdata));
  assign f502_clk = clk;
  assign f502_rst = rst;
  // Bindings to f502

  // f504
  logic [0:0] f504_wen;
  logic [31:0] f504_wdata;
  logic [0:0] f504_clk;
  logic [0:0] f504_rst;
  logic [31:0] f504_rdata;
  sr_buffer_32_1 f504(.wen(f504_wen), .wdata(f504_wdata), .clk(f504_clk), .rst(f504_rst), .rdata(f504_rdata));
  assign f504_clk = clk;
  assign f504_rst = rst;
  // Bindings to f504

  // f506
  logic [0:0] f506_wen;
  logic [31:0] f506_wdata;
  logic [0:0] f506_clk;
  logic [0:0] f506_rst;
  logic [31:0] f506_rdata;
  sr_buffer_32_1 f506(.wen(f506_wen), .wdata(f506_wdata), .clk(f506_clk), .rst(f506_rst), .rdata(f506_rdata));
  assign f506_clk = clk;
  assign f506_rst = rst;
  // Bindings to f506

  // f508
  logic [0:0] f508_wen;
  logic [31:0] f508_wdata;
  logic [0:0] f508_clk;
  logic [0:0] f508_rst;
  logic [31:0] f508_rdata;
  sr_buffer_32_1 f508(.wen(f508_wen), .wdata(f508_wdata), .clk(f508_clk), .rst(f508_rst), .rdata(f508_rdata));
  assign f508_clk = clk;
  assign f508_rst = rst;
  // Bindings to f508

  // f510
  logic [0:0] f510_wen;
  logic [31:0] f510_wdata;
  logic [0:0] f510_clk;
  logic [0:0] f510_rst;
  logic [31:0] f510_rdata;
  sr_buffer_32_1 f510(.wen(f510_wen), .wdata(f510_wdata), .clk(f510_clk), .rst(f510_rst), .rdata(f510_rdata));
  assign f510_clk = clk;
  assign f510_rst = rst;
  // Bindings to f510

  // f512
  logic [0:0] f512_wen;
  logic [31:0] f512_wdata;
  logic [0:0] f512_clk;
  logic [0:0] f512_rst;
  logic [31:0] f512_rdata;
  sr_buffer_32_1 f512(.wen(f512_wen), .wdata(f512_wdata), .clk(f512_clk), .rst(f512_rst), .rdata(f512_rdata));
  assign f512_clk = clk;
  assign f512_rst = rst;
  // Bindings to f512

  // f514
  logic [0:0] f514_wen;
  logic [31:0] f514_wdata;
  logic [0:0] f514_clk;
  logic [0:0] f514_rst;
  logic [31:0] f514_rdata;
  sr_buffer_32_1 f514(.wen(f514_wen), .wdata(f514_wdata), .clk(f514_clk), .rst(f514_rst), .rdata(f514_rdata));
  assign f514_clk = clk;
  assign f514_rst = rst;
  // Bindings to f514

  // f516
  logic [0:0] f516_wen;
  logic [31:0] f516_wdata;
  logic [0:0] f516_clk;
  logic [0:0] f516_rst;
  logic [31:0] f516_rdata;
  sr_buffer_32_1 f516(.wen(f516_wen), .wdata(f516_wdata), .clk(f516_clk), .rst(f516_rst), .rdata(f516_rdata));
  assign f516_clk = clk;
  assign f516_rst = rst;
  // Bindings to f516

  // f518
  logic [0:0] f518_wen;
  logic [31:0] f518_wdata;
  logic [0:0] f518_clk;
  logic [0:0] f518_rst;
  logic [31:0] f518_rdata;
  sr_buffer_32_1 f518(.wen(f518_wen), .wdata(f518_wdata), .clk(f518_clk), .rst(f518_rst), .rdata(f518_rdata));
  assign f518_clk = clk;
  assign f518_rst = rst;
  // Bindings to f518

  // f520
  logic [0:0] f520_wen;
  logic [31:0] f520_wdata;
  logic [0:0] f520_clk;
  logic [0:0] f520_rst;
  logic [31:0] f520_rdata;
  sr_buffer_32_1 f520(.wen(f520_wen), .wdata(f520_wdata), .clk(f520_clk), .rst(f520_rst), .rdata(f520_rdata));
  assign f520_clk = clk;
  assign f520_rst = rst;
  // Bindings to f520

  // f522
  logic [0:0] f522_wen;
  logic [31:0] f522_wdata;
  logic [0:0] f522_clk;
  logic [0:0] f522_rst;
  logic [31:0] f522_rdata;
  sr_buffer_32_1 f522(.wen(f522_wen), .wdata(f522_wdata), .clk(f522_clk), .rst(f522_rst), .rdata(f522_rdata));
  assign f522_clk = clk;
  assign f522_rst = rst;
  // Bindings to f522

  // f524
  logic [0:0] f524_wen;
  logic [31:0] f524_wdata;
  logic [0:0] f524_clk;
  logic [0:0] f524_rst;
  logic [31:0] f524_rdata;
  sr_buffer_32_1 f524(.wen(f524_wen), .wdata(f524_wdata), .clk(f524_clk), .rst(f524_rst), .rdata(f524_rdata));
  assign f524_clk = clk;
  assign f524_rst = rst;
  // Bindings to f524

  // f526
  logic [0:0] f526_wen;
  logic [31:0] f526_wdata;
  logic [0:0] f526_clk;
  logic [0:0] f526_rst;
  logic [31:0] f526_rdata;
  sr_buffer_32_1 f526(.wen(f526_wen), .wdata(f526_wdata), .clk(f526_clk), .rst(f526_rst), .rdata(f526_rdata));
  assign f526_clk = clk;
  assign f526_rst = rst;
  // Bindings to f526

  // f528
  logic [0:0] f528_wen;
  logic [31:0] f528_wdata;
  logic [0:0] f528_clk;
  logic [0:0] f528_rst;
  logic [31:0] f528_rdata;
  sr_buffer_32_1 f528(.wen(f528_wen), .wdata(f528_wdata), .clk(f528_clk), .rst(f528_rst), .rdata(f528_rdata));
  assign f528_clk = clk;
  assign f528_rst = rst;
  // Bindings to f528

  // f530
  logic [0:0] f530_wen;
  logic [31:0] f530_wdata;
  logic [0:0] f530_clk;
  logic [0:0] f530_rst;
  logic [31:0] f530_rdata;
  sr_buffer_32_1 f530(.wen(f530_wen), .wdata(f530_wdata), .clk(f530_clk), .rst(f530_rst), .rdata(f530_rdata));
  assign f530_clk = clk;
  assign f530_rst = rst;
  // Bindings to f530

  // f532
  logic [0:0] f532_wen;
  logic [31:0] f532_wdata;
  logic [0:0] f532_clk;
  logic [0:0] f532_rst;
  logic [31:0] f532_rdata;
  sr_buffer_32_1 f532(.wen(f532_wen), .wdata(f532_wdata), .clk(f532_clk), .rst(f532_rst), .rdata(f532_rdata));
  assign f532_clk = clk;
  assign f532_rst = rst;
  // Bindings to f532

  // f534
  logic [0:0] f534_wen;
  logic [31:0] f534_wdata;
  logic [0:0] f534_clk;
  logic [0:0] f534_rst;
  logic [31:0] f534_rdata;
  sr_buffer_32_1 f534(.wen(f534_wen), .wdata(f534_wdata), .clk(f534_clk), .rst(f534_rst), .rdata(f534_rdata));
  assign f534_clk = clk;
  assign f534_rst = rst;
  // Bindings to f534

  // f536
  logic [0:0] f536_wen;
  logic [31:0] f536_wdata;
  logic [0:0] f536_clk;
  logic [0:0] f536_rst;
  logic [31:0] f536_rdata;
  sr_buffer_32_1 f536(.wen(f536_wen), .wdata(f536_wdata), .clk(f536_clk), .rst(f536_rst), .rdata(f536_rdata));
  assign f536_clk = clk;
  assign f536_rst = rst;
  // Bindings to f536

  // f538
  logic [0:0] f538_wen;
  logic [31:0] f538_wdata;
  logic [0:0] f538_clk;
  logic [0:0] f538_rst;
  logic [31:0] f538_rdata;
  sr_buffer_32_1 f538(.wen(f538_wen), .wdata(f538_wdata), .clk(f538_clk), .rst(f538_rst), .rdata(f538_rdata));
  assign f538_clk = clk;
  assign f538_rst = rst;
  // Bindings to f538

  // f540
  logic [0:0] f540_wen;
  logic [31:0] f540_wdata;
  logic [0:0] f540_clk;
  logic [0:0] f540_rst;
  logic [31:0] f540_rdata;
  sr_buffer_32_1 f540(.wen(f540_wen), .wdata(f540_wdata), .clk(f540_clk), .rst(f540_rst), .rdata(f540_rdata));
  assign f540_clk = clk;
  assign f540_rst = rst;
  // Bindings to f540

  // f542
  logic [0:0] f542_wen;
  logic [31:0] f542_wdata;
  logic [0:0] f542_clk;
  logic [0:0] f542_rst;
  logic [31:0] f542_rdata;
  sr_buffer_32_1 f542(.wen(f542_wen), .wdata(f542_wdata), .clk(f542_clk), .rst(f542_rst), .rdata(f542_rdata));
  assign f542_clk = clk;
  assign f542_rst = rst;
  // Bindings to f542

  // f544
  logic [0:0] f544_wen;
  logic [31:0] f544_wdata;
  logic [0:0] f544_clk;
  logic [0:0] f544_rst;
  logic [31:0] f544_rdata;
  sr_buffer_32_1 f544(.wen(f544_wen), .wdata(f544_wdata), .clk(f544_clk), .rst(f544_rst), .rdata(f544_rdata));
  assign f544_clk = clk;
  assign f544_rst = rst;
  // Bindings to f544

  // f546
  logic [0:0] f546_wen;
  logic [31:0] f546_wdata;
  logic [0:0] f546_clk;
  logic [0:0] f546_rst;
  logic [31:0] f546_rdata;
  sr_buffer_32_1 f546(.wen(f546_wen), .wdata(f546_wdata), .clk(f546_clk), .rst(f546_rst), .rdata(f546_rdata));
  assign f546_clk = clk;
  assign f546_rst = rst;
  // Bindings to f546

  // f548
  logic [0:0] f548_wen;
  logic [31:0] f548_wdata;
  logic [0:0] f548_clk;
  logic [0:0] f548_rst;
  logic [31:0] f548_rdata;
  sr_buffer_32_1 f548(.wen(f548_wen), .wdata(f548_wdata), .clk(f548_clk), .rst(f548_rst), .rdata(f548_rdata));
  assign f548_clk = clk;
  assign f548_rst = rst;
  // Bindings to f548

  // f550
  logic [0:0] f550_wen;
  logic [31:0] f550_wdata;
  logic [0:0] f550_clk;
  logic [0:0] f550_rst;
  logic [31:0] f550_rdata;
  sr_buffer_32_1 f550(.wen(f550_wen), .wdata(f550_wdata), .clk(f550_clk), .rst(f550_rst), .rdata(f550_rdata));
  assign f550_clk = clk;
  assign f550_rst = rst;
  // Bindings to f550

  // f552
  logic [0:0] f552_wen;
  logic [31:0] f552_wdata;
  logic [0:0] f552_clk;
  logic [0:0] f552_rst;
  logic [31:0] f552_rdata;
  sr_buffer_32_1 f552(.wen(f552_wen), .wdata(f552_wdata), .clk(f552_clk), .rst(f552_rst), .rdata(f552_rdata));
  assign f552_clk = clk;
  assign f552_rst = rst;
  // Bindings to f552

  // f554
  logic [0:0] f554_wen;
  logic [31:0] f554_wdata;
  logic [0:0] f554_clk;
  logic [0:0] f554_rst;
  logic [31:0] f554_rdata;
  sr_buffer_32_1 f554(.wen(f554_wen), .wdata(f554_wdata), .clk(f554_clk), .rst(f554_rst), .rdata(f554_rdata));
  assign f554_clk = clk;
  assign f554_rst = rst;
  // Bindings to f554

  // f556
  logic [0:0] f556_wen;
  logic [31:0] f556_wdata;
  logic [0:0] f556_clk;
  logic [0:0] f556_rst;
  logic [31:0] f556_rdata;
  sr_buffer_32_1 f556(.wen(f556_wen), .wdata(f556_wdata), .clk(f556_clk), .rst(f556_rst), .rdata(f556_rdata));
  assign f556_clk = clk;
  assign f556_rst = rst;
  // Bindings to f556

  // f558
  logic [0:0] f558_wen;
  logic [31:0] f558_wdata;
  logic [0:0] f558_clk;
  logic [0:0] f558_rst;
  logic [31:0] f558_rdata;
  sr_buffer_32_1 f558(.wen(f558_wen), .wdata(f558_wdata), .clk(f558_clk), .rst(f558_rst), .rdata(f558_rdata));
  assign f558_clk = clk;
  assign f558_rst = rst;
  // Bindings to f558

  // f560
  logic [0:0] f560_wen;
  logic [31:0] f560_wdata;
  logic [0:0] f560_clk;
  logic [0:0] f560_rst;
  logic [31:0] f560_rdata;
  sr_buffer_32_1 f560(.wen(f560_wen), .wdata(f560_wdata), .clk(f560_clk), .rst(f560_rst), .rdata(f560_rdata));
  assign f560_clk = clk;
  assign f560_rst = rst;
  // Bindings to f560

  // f562
  logic [0:0] f562_wen;
  logic [31:0] f562_wdata;
  logic [0:0] f562_clk;
  logic [0:0] f562_rst;
  logic [31:0] f562_rdata;
  sr_buffer_32_1 f562(.wen(f562_wen), .wdata(f562_wdata), .clk(f562_clk), .rst(f562_rst), .rdata(f562_rdata));
  assign f562_clk = clk;
  assign f562_rst = rst;
  // Bindings to f562

  // f564
  logic [0:0] f564_wen;
  logic [31:0] f564_wdata;
  logic [0:0] f564_clk;
  logic [0:0] f564_rst;
  logic [31:0] f564_rdata;
  sr_buffer_32_1 f564(.wen(f564_wen), .wdata(f564_wdata), .clk(f564_clk), .rst(f564_rst), .rdata(f564_rdata));
  assign f564_clk = clk;
  assign f564_rst = rst;
  // Bindings to f564

  // f566
  logic [0:0] f566_wen;
  logic [31:0] f566_wdata;
  logic [0:0] f566_clk;
  logic [0:0] f566_rst;
  logic [31:0] f566_rdata;
  sr_buffer_32_1 f566(.wen(f566_wen), .wdata(f566_wdata), .clk(f566_clk), .rst(f566_rst), .rdata(f566_rdata));
  assign f566_clk = clk;
  assign f566_rst = rst;
  // Bindings to f566

  // f568
  logic [0:0] f568_wen;
  logic [31:0] f568_wdata;
  logic [0:0] f568_clk;
  logic [0:0] f568_rst;
  logic [31:0] f568_rdata;
  sr_buffer_32_1 f568(.wen(f568_wen), .wdata(f568_wdata), .clk(f568_clk), .rst(f568_rst), .rdata(f568_rdata));
  assign f568_clk = clk;
  assign f568_rst = rst;
  // Bindings to f568

  // f570
  logic [0:0] f570_wen;
  logic [31:0] f570_wdata;
  logic [0:0] f570_clk;
  logic [0:0] f570_rst;
  logic [31:0] f570_rdata;
  sr_buffer_32_1 f570(.wen(f570_wen), .wdata(f570_wdata), .clk(f570_clk), .rst(f570_rst), .rdata(f570_rdata));
  assign f570_clk = clk;
  assign f570_rst = rst;
  // Bindings to f570

  // f572
  logic [0:0] f572_wen;
  logic [31:0] f572_wdata;
  logic [0:0] f572_clk;
  logic [0:0] f572_rst;
  logic [31:0] f572_rdata;
  sr_buffer_32_1 f572(.wen(f572_wen), .wdata(f572_wdata), .clk(f572_clk), .rst(f572_rst), .rdata(f572_rdata));
  assign f572_clk = clk;
  assign f572_rst = rst;
  // Bindings to f572

  // f574
  logic [0:0] f574_wen;
  logic [31:0] f574_wdata;
  logic [0:0] f574_clk;
  logic [0:0] f574_rst;
  logic [31:0] f574_rdata;
  sr_buffer_32_1 f574(.wen(f574_wen), .wdata(f574_wdata), .clk(f574_clk), .rst(f574_rst), .rdata(f574_rdata));
  assign f574_clk = clk;
  assign f574_rst = rst;
  // Bindings to f574

  // f576
  logic [0:0] f576_wen;
  logic [31:0] f576_wdata;
  logic [0:0] f576_clk;
  logic [0:0] f576_rst;
  logic [31:0] f576_rdata;
  sr_buffer_32_1 f576(.wen(f576_wen), .wdata(f576_wdata), .clk(f576_clk), .rst(f576_rst), .rdata(f576_rdata));
  assign f576_clk = clk;
  assign f576_rst = rst;
  // Bindings to f576

  // f578
  logic [0:0] f578_wen;
  logic [31:0] f578_wdata;
  logic [0:0] f578_clk;
  logic [0:0] f578_rst;
  logic [31:0] f578_rdata;
  sr_buffer_32_1 f578(.wen(f578_wen), .wdata(f578_wdata), .clk(f578_clk), .rst(f578_rst), .rdata(f578_rdata));
  assign f578_clk = clk;
  assign f578_rst = rst;
  // Bindings to f578

  // f580
  logic [0:0] f580_wen;
  logic [31:0] f580_wdata;
  logic [0:0] f580_clk;
  logic [0:0] f580_rst;
  logic [31:0] f580_rdata;
  sr_buffer_32_1 f580(.wen(f580_wen), .wdata(f580_wdata), .clk(f580_clk), .rst(f580_rst), .rdata(f580_rdata));
  assign f580_clk = clk;
  assign f580_rst = rst;
  // Bindings to f580

  // f582
  logic [0:0] f582_wen;
  logic [31:0] f582_wdata;
  logic [0:0] f582_clk;
  logic [0:0] f582_rst;
  logic [31:0] f582_rdata;
  sr_buffer_32_1 f582(.wen(f582_wen), .wdata(f582_wdata), .clk(f582_clk), .rst(f582_rst), .rdata(f582_rdata));
  assign f582_clk = clk;
  assign f582_rst = rst;
  // Bindings to f582

  // f584
  logic [0:0] f584_wen;
  logic [31:0] f584_wdata;
  logic [0:0] f584_clk;
  logic [0:0] f584_rst;
  logic [31:0] f584_rdata;
  sr_buffer_32_1 f584(.wen(f584_wen), .wdata(f584_wdata), .clk(f584_clk), .rst(f584_rst), .rdata(f584_rdata));
  assign f584_clk = clk;
  assign f584_rst = rst;
  // Bindings to f584

  // f586
  logic [0:0] f586_wen;
  logic [31:0] f586_wdata;
  logic [0:0] f586_clk;
  logic [0:0] f586_rst;
  logic [31:0] f586_rdata;
  sr_buffer_32_1 f586(.wen(f586_wen), .wdata(f586_wdata), .clk(f586_clk), .rst(f586_rst), .rdata(f586_rdata));
  assign f586_clk = clk;
  assign f586_rst = rst;
  // Bindings to f586

  // f588
  logic [0:0] f588_wen;
  logic [31:0] f588_wdata;
  logic [0:0] f588_clk;
  logic [0:0] f588_rst;
  logic [31:0] f588_rdata;
  sr_buffer_32_1 f588(.wen(f588_wen), .wdata(f588_wdata), .clk(f588_clk), .rst(f588_rst), .rdata(f588_rdata));
  assign f588_clk = clk;
  assign f588_rst = rst;
  // Bindings to f588

  // f590
  logic [0:0] f590_wen;
  logic [31:0] f590_wdata;
  logic [0:0] f590_clk;
  logic [0:0] f590_rst;
  logic [31:0] f590_rdata;
  sr_buffer_32_1 f590(.wen(f590_wen), .wdata(f590_wdata), .clk(f590_clk), .rst(f590_rst), .rdata(f590_rdata));
  assign f590_clk = clk;
  assign f590_rst = rst;
  // Bindings to f590

  // f592
  logic [0:0] f592_wen;
  logic [31:0] f592_wdata;
  logic [0:0] f592_clk;
  logic [0:0] f592_rst;
  logic [31:0] f592_rdata;
  sr_buffer_32_1 f592(.wen(f592_wen), .wdata(f592_wdata), .clk(f592_clk), .rst(f592_rst), .rdata(f592_rdata));
  assign f592_clk = clk;
  assign f592_rst = rst;
  // Bindings to f592

  // f594
  logic [0:0] f594_wen;
  logic [31:0] f594_wdata;
  logic [0:0] f594_clk;
  logic [0:0] f594_rst;
  logic [31:0] f594_rdata;
  sr_buffer_32_1 f594(.wen(f594_wen), .wdata(f594_wdata), .clk(f594_clk), .rst(f594_rst), .rdata(f594_rdata));
  assign f594_clk = clk;
  assign f594_rst = rst;
  // Bindings to f594

  // f596
  logic [0:0] f596_wen;
  logic [31:0] f596_wdata;
  logic [0:0] f596_clk;
  logic [0:0] f596_rst;
  logic [31:0] f596_rdata;
  sr_buffer_32_1 f596(.wen(f596_wen), .wdata(f596_wdata), .clk(f596_clk), .rst(f596_rst), .rdata(f596_rdata));
  assign f596_clk = clk;
  assign f596_rst = rst;
  // Bindings to f596

  // f598
  logic [0:0] f598_wen;
  logic [31:0] f598_wdata;
  logic [0:0] f598_clk;
  logic [0:0] f598_rst;
  logic [31:0] f598_rdata;
  sr_buffer_32_1 f598(.wen(f598_wen), .wdata(f598_wdata), .clk(f598_clk), .rst(f598_rst), .rdata(f598_rdata));
  assign f598_clk = clk;
  assign f598_rst = rst;
  // Bindings to f598

  // f600
  logic [0:0] f600_wen;
  logic [31:0] f600_wdata;
  logic [0:0] f600_clk;
  logic [0:0] f600_rst;
  logic [31:0] f600_rdata;
  sr_buffer_32_1 f600(.wen(f600_wen), .wdata(f600_wdata), .clk(f600_clk), .rst(f600_rst), .rdata(f600_rdata));
  assign f600_clk = clk;
  assign f600_rst = rst;
  // Bindings to f600

  // f602
  logic [0:0] f602_wen;
  logic [31:0] f602_wdata;
  logic [0:0] f602_clk;
  logic [0:0] f602_rst;
  logic [31:0] f602_rdata;
  sr_buffer_32_1 f602(.wen(f602_wen), .wdata(f602_wdata), .clk(f602_clk), .rst(f602_rst), .rdata(f602_rdata));
  assign f602_clk = clk;
  assign f602_rst = rst;
  // Bindings to f602

  // f604
  logic [0:0] f604_wen;
  logic [31:0] f604_wdata;
  logic [0:0] f604_clk;
  logic [0:0] f604_rst;
  logic [31:0] f604_rdata;
  sr_buffer_32_1 f604(.wen(f604_wen), .wdata(f604_wdata), .clk(f604_clk), .rst(f604_rst), .rdata(f604_rdata));
  assign f604_clk = clk;
  assign f604_rst = rst;
  // Bindings to f604

  // f606
  logic [0:0] f606_wen;
  logic [31:0] f606_wdata;
  logic [0:0] f606_clk;
  logic [0:0] f606_rst;
  logic [31:0] f606_rdata;
  sr_buffer_32_1 f606(.wen(f606_wen), .wdata(f606_wdata), .clk(f606_clk), .rst(f606_rst), .rdata(f606_rdata));
  assign f606_clk = clk;
  assign f606_rst = rst;
  // Bindings to f606

  // f608
  logic [0:0] f608_wen;
  logic [31:0] f608_wdata;
  logic [0:0] f608_clk;
  logic [0:0] f608_rst;
  logic [31:0] f608_rdata;
  sr_buffer_32_1 f608(.wen(f608_wen), .wdata(f608_wdata), .clk(f608_clk), .rst(f608_rst), .rdata(f608_rdata));
  assign f608_clk = clk;
  assign f608_rst = rst;
  // Bindings to f608

  // f610
  logic [0:0] f610_wen;
  logic [31:0] f610_wdata;
  logic [0:0] f610_clk;
  logic [0:0] f610_rst;
  logic [31:0] f610_rdata;
  sr_buffer_32_1 f610(.wen(f610_wen), .wdata(f610_wdata), .clk(f610_clk), .rst(f610_rst), .rdata(f610_rdata));
  assign f610_clk = clk;
  assign f610_rst = rst;
  // Bindings to f610

  // f612
  logic [0:0] f612_wen;
  logic [31:0] f612_wdata;
  logic [0:0] f612_clk;
  logic [0:0] f612_rst;
  logic [31:0] f612_rdata;
  sr_buffer_32_1 f612(.wen(f612_wen), .wdata(f612_wdata), .clk(f612_clk), .rst(f612_rst), .rdata(f612_rdata));
  assign f612_clk = clk;
  assign f612_rst = rst;
  // Bindings to f612

  // f614
  logic [0:0] f614_wen;
  logic [31:0] f614_wdata;
  logic [0:0] f614_clk;
  logic [0:0] f614_rst;
  logic [31:0] f614_rdata;
  sr_buffer_32_1 f614(.wen(f614_wen), .wdata(f614_wdata), .clk(f614_clk), .rst(f614_rst), .rdata(f614_rdata));
  assign f614_clk = clk;
  assign f614_rst = rst;
  // Bindings to f614

  // f616
  logic [0:0] f616_wen;
  logic [31:0] f616_wdata;
  logic [0:0] f616_clk;
  logic [0:0] f616_rst;
  logic [31:0] f616_rdata;
  sr_buffer_32_1 f616(.wen(f616_wen), .wdata(f616_wdata), .clk(f616_clk), .rst(f616_rst), .rdata(f616_rdata));
  assign f616_clk = clk;
  assign f616_rst = rst;
  // Bindings to f616

  // f618
  logic [0:0] f618_wen;
  logic [31:0] f618_wdata;
  logic [0:0] f618_clk;
  logic [0:0] f618_rst;
  logic [31:0] f618_rdata;
  sr_buffer_32_1 f618(.wen(f618_wen), .wdata(f618_wdata), .clk(f618_clk), .rst(f618_rst), .rdata(f618_rdata));
  assign f618_clk = clk;
  assign f618_rst = rst;
  // Bindings to f618

  // f620
  logic [0:0] f620_wen;
  logic [31:0] f620_wdata;
  logic [0:0] f620_clk;
  logic [0:0] f620_rst;
  logic [31:0] f620_rdata;
  sr_buffer_32_1 f620(.wen(f620_wen), .wdata(f620_wdata), .clk(f620_clk), .rst(f620_rst), .rdata(f620_rdata));
  assign f620_clk = clk;
  assign f620_rst = rst;
  // Bindings to f620

  // f622
  logic [0:0] f622_wen;
  logic [31:0] f622_wdata;
  logic [0:0] f622_clk;
  logic [0:0] f622_rst;
  logic [31:0] f622_rdata;
  sr_buffer_32_1 f622(.wen(f622_wen), .wdata(f622_wdata), .clk(f622_clk), .rst(f622_rst), .rdata(f622_rdata));
  assign f622_clk = clk;
  assign f622_rst = rst;
  // Bindings to f622

  // f624
  logic [0:0] f624_wen;
  logic [31:0] f624_wdata;
  logic [0:0] f624_clk;
  logic [0:0] f624_rst;
  logic [31:0] f624_rdata;
  sr_buffer_32_1 f624(.wen(f624_wen), .wdata(f624_wdata), .clk(f624_clk), .rst(f624_rst), .rdata(f624_rdata));
  assign f624_clk = clk;
  assign f624_rst = rst;
  // Bindings to f624

  // f626
  logic [0:0] f626_wen;
  logic [31:0] f626_wdata;
  logic [0:0] f626_clk;
  logic [0:0] f626_rst;
  logic [31:0] f626_rdata;
  sr_buffer_32_1 f626(.wen(f626_wen), .wdata(f626_wdata), .clk(f626_clk), .rst(f626_rst), .rdata(f626_rdata));
  assign f626_clk = clk;
  assign f626_rst = rst;
  // Bindings to f626

  // f628
  logic [0:0] f628_wen;
  logic [31:0] f628_wdata;
  logic [0:0] f628_clk;
  logic [0:0] f628_rst;
  logic [31:0] f628_rdata;
  sr_buffer_32_1 f628(.wen(f628_wen), .wdata(f628_wdata), .clk(f628_clk), .rst(f628_rst), .rdata(f628_rdata));
  assign f628_clk = clk;
  assign f628_rst = rst;
  // Bindings to f628

  // f630
  logic [0:0] f630_wen;
  logic [31:0] f630_wdata;
  logic [0:0] f630_clk;
  logic [0:0] f630_rst;
  logic [31:0] f630_rdata;
  sr_buffer_32_1 f630(.wen(f630_wen), .wdata(f630_wdata), .clk(f630_clk), .rst(f630_rst), .rdata(f630_rdata));
  assign f630_clk = clk;
  assign f630_rst = rst;
  // Bindings to f630

  // f632
  logic [0:0] f632_wen;
  logic [31:0] f632_wdata;
  logic [0:0] f632_clk;
  logic [0:0] f632_rst;
  logic [31:0] f632_rdata;
  sr_buffer_32_1 f632(.wen(f632_wen), .wdata(f632_wdata), .clk(f632_clk), .rst(f632_rst), .rdata(f632_rdata));
  assign f632_clk = clk;
  assign f632_rst = rst;
  // Bindings to f632

  // f634
  logic [0:0] f634_wen;
  logic [31:0] f634_wdata;
  logic [0:0] f634_clk;
  logic [0:0] f634_rst;
  logic [31:0] f634_rdata;
  sr_buffer_32_1 f634(.wen(f634_wen), .wdata(f634_wdata), .clk(f634_clk), .rst(f634_rst), .rdata(f634_rdata));
  assign f634_clk = clk;
  assign f634_rst = rst;
  // Bindings to f634

  // f636
  logic [0:0] f636_wen;
  logic [31:0] f636_wdata;
  logic [0:0] f636_clk;
  logic [0:0] f636_rst;
  logic [31:0] f636_rdata;
  sr_buffer_32_1 f636(.wen(f636_wen), .wdata(f636_wdata), .clk(f636_clk), .rst(f636_rst), .rdata(f636_rdata));
  assign f636_clk = clk;
  assign f636_rst = rst;
  // Bindings to f636

  // f638
  logic [0:0] f638_wen;
  logic [31:0] f638_wdata;
  logic [0:0] f638_clk;
  logic [0:0] f638_rst;
  logic [31:0] f638_rdata;
  sr_buffer_32_1 f638(.wen(f638_wen), .wdata(f638_wdata), .clk(f638_clk), .rst(f638_rst), .rdata(f638_rdata));
  assign f638_clk = clk;
  assign f638_rst = rst;
  // Bindings to f638

  // f640
  logic [0:0] f640_wen;
  logic [31:0] f640_wdata;
  logic [0:0] f640_clk;
  logic [0:0] f640_rst;
  logic [31:0] f640_rdata;
  sr_buffer_32_1 f640(.wen(f640_wen), .wdata(f640_wdata), .clk(f640_clk), .rst(f640_rst), .rdata(f640_rdata));
  assign f640_clk = clk;
  assign f640_rst = rst;
  // Bindings to f640

  // f642
  logic [0:0] f642_wen;
  logic [31:0] f642_wdata;
  logic [0:0] f642_clk;
  logic [0:0] f642_rst;
  logic [31:0] f642_rdata;
  sr_buffer_32_1 f642(.wen(f642_wen), .wdata(f642_wdata), .clk(f642_clk), .rst(f642_rst), .rdata(f642_rdata));
  assign f642_clk = clk;
  assign f642_rst = rst;
  // Bindings to f642

  // f644
  logic [0:0] f644_wen;
  logic [31:0] f644_wdata;
  logic [0:0] f644_clk;
  logic [0:0] f644_rst;
  logic [31:0] f644_rdata;
  sr_buffer_32_1 f644(.wen(f644_wen), .wdata(f644_wdata), .clk(f644_clk), .rst(f644_rst), .rdata(f644_rdata));
  assign f644_clk = clk;
  assign f644_rst = rst;
  // Bindings to f644

  // f646
  logic [0:0] f646_wen;
  logic [31:0] f646_wdata;
  logic [0:0] f646_clk;
  logic [0:0] f646_rst;
  logic [31:0] f646_rdata;
  sr_buffer_32_1 f646(.wen(f646_wen), .wdata(f646_wdata), .clk(f646_clk), .rst(f646_rst), .rdata(f646_rdata));
  assign f646_clk = clk;
  assign f646_rst = rst;
  // Bindings to f646

  // f648
  logic [0:0] f648_wen;
  logic [31:0] f648_wdata;
  logic [0:0] f648_clk;
  logic [0:0] f648_rst;
  logic [31:0] f648_rdata;
  sr_buffer_32_1 f648(.wen(f648_wen), .wdata(f648_wdata), .clk(f648_clk), .rst(f648_rst), .rdata(f648_rdata));
  assign f648_clk = clk;
  assign f648_rst = rst;
  // Bindings to f648

  // f650
  logic [0:0] f650_wen;
  logic [31:0] f650_wdata;
  logic [0:0] f650_clk;
  logic [0:0] f650_rst;
  logic [31:0] f650_rdata;
  sr_buffer_32_1 f650(.wen(f650_wen), .wdata(f650_wdata), .clk(f650_clk), .rst(f650_rst), .rdata(f650_rdata));
  assign f650_clk = clk;
  assign f650_rst = rst;
  // Bindings to f650

  // f652
  logic [0:0] f652_wen;
  logic [31:0] f652_wdata;
  logic [0:0] f652_clk;
  logic [0:0] f652_rst;
  logic [31:0] f652_rdata;
  sr_buffer_32_1 f652(.wen(f652_wen), .wdata(f652_wdata), .clk(f652_clk), .rst(f652_rst), .rdata(f652_rdata));
  assign f652_clk = clk;
  assign f652_rst = rst;
  // Bindings to f652

  // f654
  logic [0:0] f654_wen;
  logic [31:0] f654_wdata;
  logic [0:0] f654_clk;
  logic [0:0] f654_rst;
  logic [31:0] f654_rdata;
  sr_buffer_32_1 f654(.wen(f654_wen), .wdata(f654_wdata), .clk(f654_clk), .rst(f654_rst), .rdata(f654_rdata));
  assign f654_clk = clk;
  assign f654_rst = rst;
  // Bindings to f654

  // f656
  logic [0:0] f656_wen;
  logic [31:0] f656_wdata;
  logic [0:0] f656_clk;
  logic [0:0] f656_rst;
  logic [31:0] f656_rdata;
  sr_buffer_32_1 f656(.wen(f656_wen), .wdata(f656_wdata), .clk(f656_clk), .rst(f656_rst), .rdata(f656_rdata));
  assign f656_clk = clk;
  assign f656_rst = rst;
  // Bindings to f656

  // f658
  logic [0:0] f658_wen;
  logic [31:0] f658_wdata;
  logic [0:0] f658_clk;
  logic [0:0] f658_rst;
  logic [31:0] f658_rdata;
  sr_buffer_32_1 f658(.wen(f658_wen), .wdata(f658_wdata), .clk(f658_clk), .rst(f658_rst), .rdata(f658_rdata));
  assign f658_clk = clk;
  assign f658_rst = rst;
  // Bindings to f658

  // f660
  logic [0:0] f660_wen;
  logic [31:0] f660_wdata;
  logic [0:0] f660_clk;
  logic [0:0] f660_rst;
  logic [31:0] f660_rdata;
  sr_buffer_32_1 f660(.wen(f660_wen), .wdata(f660_wdata), .clk(f660_clk), .rst(f660_rst), .rdata(f660_rdata));
  assign f660_clk = clk;
  assign f660_rst = rst;
  // Bindings to f660

  // f662
  logic [0:0] f662_wen;
  logic [31:0] f662_wdata;
  logic [0:0] f662_clk;
  logic [0:0] f662_rst;
  logic [31:0] f662_rdata;
  sr_buffer_32_1 f662(.wen(f662_wen), .wdata(f662_wdata), .clk(f662_clk), .rst(f662_rst), .rdata(f662_rdata));
  assign f662_clk = clk;
  assign f662_rst = rst;
  // Bindings to f662

  // f664
  logic [0:0] f664_wen;
  logic [31:0] f664_wdata;
  logic [0:0] f664_clk;
  logic [0:0] f664_rst;
  logic [31:0] f664_rdata;
  sr_buffer_32_1 f664(.wen(f664_wen), .wdata(f664_wdata), .clk(f664_clk), .rst(f664_rst), .rdata(f664_rdata));
  assign f664_clk = clk;
  assign f664_rst = rst;
  // Bindings to f664

  // f666
  logic [0:0] f666_wen;
  logic [31:0] f666_wdata;
  logic [0:0] f666_clk;
  logic [0:0] f666_rst;
  logic [31:0] f666_rdata;
  sr_buffer_32_1 f666(.wen(f666_wen), .wdata(f666_wdata), .clk(f666_clk), .rst(f666_rst), .rdata(f666_rdata));
  assign f666_clk = clk;
  assign f666_rst = rst;
  // Bindings to f666

  // f668
  logic [0:0] f668_wen;
  logic [31:0] f668_wdata;
  logic [0:0] f668_clk;
  logic [0:0] f668_rst;
  logic [31:0] f668_rdata;
  sr_buffer_32_1 f668(.wen(f668_wen), .wdata(f668_wdata), .clk(f668_clk), .rst(f668_rst), .rdata(f668_rdata));
  assign f668_clk = clk;
  assign f668_rst = rst;
  // Bindings to f668

  // f670
  logic [0:0] f670_wen;
  logic [31:0] f670_wdata;
  logic [0:0] f670_clk;
  logic [0:0] f670_rst;
  logic [31:0] f670_rdata;
  sr_buffer_32_1 f670(.wen(f670_wen), .wdata(f670_wdata), .clk(f670_clk), .rst(f670_rst), .rdata(f670_rdata));
  assign f670_clk = clk;
  assign f670_rst = rst;
  // Bindings to f670

  // f672
  logic [0:0] f672_wen;
  logic [31:0] f672_wdata;
  logic [0:0] f672_clk;
  logic [0:0] f672_rst;
  logic [31:0] f672_rdata;
  sr_buffer_32_1 f672(.wen(f672_wen), .wdata(f672_wdata), .clk(f672_clk), .rst(f672_rst), .rdata(f672_rdata));
  assign f672_clk = clk;
  assign f672_rst = rst;
  // Bindings to f672

  // f674
  logic [0:0] f674_wen;
  logic [31:0] f674_wdata;
  logic [0:0] f674_clk;
  logic [0:0] f674_rst;
  logic [31:0] f674_rdata;
  sr_buffer_32_1 f674(.wen(f674_wen), .wdata(f674_wdata), .clk(f674_clk), .rst(f674_rst), .rdata(f674_rdata));
  assign f674_clk = clk;
  assign f674_rst = rst;
  // Bindings to f674



endmodule


module fused_level_0_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (-97 + d0 == 0 && 96 - d1 >= 0) ? (1567) : (96 - d1 >= 0 && 96 - d0 >= 0) ? (1568) : (-97 + d1 == 0) ? ((1553 - d0)) : (-98 + d0 >= 0 && 96 - d1 >= 0) ? ((1664 - d0)) : (-98 + d1 >= 0) ? (((12320 - d0) - 111 * d1)) : 0;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 113;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 224;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 223;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (107 - d0 >= 0) ? (222) : (-108 + d0 == 0) ? (222) : 0;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 112;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_update_0_write_wen(output [0:0] dark_weights_normed_update_0_write_wen);

endmodule


module dark_weights_normed_gauss_blur_1_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (107 - d0 >= 0) ? (111) : (-108 + d0 == 0) ? (111) : 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_update_0_write_wdata(output [31:0] dark_weights_normed_update_0_write_wdata);

endmodule


module in_wire_dark_weights_normed_gauss_blur_1_update_0_read_dummy(output [287:0] dark_weights_normed_gauss_blur_1_update_0_read_dummy);

endmodule


module out_wire_dark_weights_normed_gauss_blur_1_update_0_read_rdata(input [287:0] dark_weights_normed_gauss_blur_1_update_0_read_rdata);

endmodule


module dark_weights_normed_gauss_ds_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_weights_normed_gauss_blur_1_update_0_write_wen(output [0:0] dark_weights_normed_gauss_blur_1_update_0_write_wen);

endmodule


module in_wire_dark_weights_normed_gauss_blur_1_update_0_write_wdata(output [31:0] dark_weights_normed_gauss_blur_1_update_0_write_wdata);

endmodule


module dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_weights_normed_gauss_ds_1_update_0_read_dummy(output [31:0] dark_weights_normed_gauss_ds_1_update_0_read_dummy);

endmodule


module out_wire_dark_weights_normed_gauss_ds_1_update_0_read_rdata(input [31:0] dark_weights_normed_gauss_ds_1_update_0_read_rdata);

endmodule


module in_wire_dark_weights_normed_gauss_blur_2_update_0_write_wen(output [0:0] dark_weights_normed_gauss_blur_2_update_0_write_wen);

endmodule


module dark_weights_normed_gauss_ds_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_gauss_blur_2_update_0_write_wdata(output [31:0] dark_weights_normed_gauss_blur_2_update_0_write_wdata);

endmodule


module in_wire_dark_weights_normed_gauss_ds_2_update_0_read_dummy(output [31:0] dark_weights_normed_gauss_ds_2_update_0_read_dummy);

endmodule


module out_wire_dark_weights_normed_gauss_ds_2_update_0_read_rdata(input [31:0] dark_weights_normed_gauss_ds_2_update_0_read_rdata);

endmodule


module dark_weights_normed_gauss_blur_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_weights_normed_gauss_blur_2_update_0_write_wen, input [31:0] dark_weights_normed_gauss_blur_2_update_0_write_wdata, input [31:0] dark_weights_normed_gauss_ds_2_update_0_read_dummy, output [31:0] dark_weights_normed_gauss_ds_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1
  logic [0:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_done;
  dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1 dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1(.clk(dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_clk), .rst(dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_rst), .start(dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_start), .done(dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_done));
  assign dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_clk = clk;
  assign dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1

  // Bindings to dark_weights_normed_gauss_blur_2_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_normed_gauss_blur_2_update_0_write_wen;

  // selector_dark_weights_normed_gauss_ds_2_rd0_select
  logic [0:0] selector_dark_weights_normed_gauss_ds_2_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_ds_2_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_ds_2_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_ds_2_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_ds_2_rd0_select_out;
  dark_weights_normed_gauss_ds_2_rd0_select selector_dark_weights_normed_gauss_ds_2_rd0_select(.clk(selector_dark_weights_normed_gauss_ds_2_rd0_select_clk), .rst(selector_dark_weights_normed_gauss_ds_2_rd0_select_rst), .d0(selector_dark_weights_normed_gauss_ds_2_rd0_select_d0), .d1(selector_dark_weights_normed_gauss_ds_2_rd0_select_d1), .out(selector_dark_weights_normed_gauss_ds_2_rd0_select_out));
  assign selector_dark_weights_normed_gauss_ds_2_rd0_select_clk = clk;
  assign selector_dark_weights_normed_gauss_ds_2_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_ds_2_rd0_select

  // Bindings to dark_weights_normed_gauss_blur_2_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_normed_gauss_blur_2_update_0_write_wdata;

  // Bindings to dark_weights_normed_gauss_ds_2_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_weights_normed_gauss_ds_2_update_0_read_dummy;

  // Bindings to dark_weights_normed_gauss_ds_2_update_0_read_rdata
    // wr_3
  assign dark_weights_normed_gauss_ds_2_update_0_read_rdata = rd_2;



endmodule


module dark_weights_normed_gauss_ds_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] fused_level_2_update_0_read_dummy, input [287:0] dark_weights_normed_gauss_blur_3_update_0_read_dummy, input [0:0] dark_weights_normed_gauss_ds_2_update_0_write_wen, input [31:0] dark_weights_normed_gauss_ds_2_update_0_write_wdata, output [287:0] dark_weights_normed_gauss_blur_3_update_0_read_rdata, output [31:0] fused_level_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // selector_dark_weights_normed_gauss_blur_3_rd2_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd2_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd2_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd2_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd2_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd2_select_out;
  dark_weights_normed_gauss_blur_3_rd2_select selector_dark_weights_normed_gauss_blur_3_rd2_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd2_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd2_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd2_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd2_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd2_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd2_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd2_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd2_select

  // dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10
  logic [0:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_clk;
  logic [0:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_rst;
  logic [0:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_start;
  logic [0:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_done;
  dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10 dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10(.clk(dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_clk), .rst(dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_rst), .start(dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_start), .done(dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_done));
  assign dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_clk = clk;
  assign dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10

  // selector_dark_weights_normed_gauss_blur_3_rd1_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd1_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd1_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd1_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd1_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd1_select_out;
  dark_weights_normed_gauss_blur_3_rd1_select selector_dark_weights_normed_gauss_blur_3_rd1_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd1_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd1_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd1_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd1_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd1_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd1_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd1_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd1_select

  // selector_dark_weights_normed_gauss_blur_3_rd0_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd0_select_out;
  dark_weights_normed_gauss_blur_3_rd0_select selector_dark_weights_normed_gauss_blur_3_rd0_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd0_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd0_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd0_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd0_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd0_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd0_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd0_select

  // selector_dark_weights_normed_gauss_blur_3_rd3_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd3_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd3_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd3_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd3_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd3_select_out;
  dark_weights_normed_gauss_blur_3_rd3_select selector_dark_weights_normed_gauss_blur_3_rd3_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd3_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd3_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd3_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd3_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd3_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd3_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd3_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd3_select

  // selector_dark_weights_normed_gauss_blur_3_rd4_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd4_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd4_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd4_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd4_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd4_select_out;
  dark_weights_normed_gauss_blur_3_rd4_select selector_dark_weights_normed_gauss_blur_3_rd4_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd4_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd4_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd4_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd4_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd4_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd4_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd4_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd4_select

  // selector_dark_weights_normed_gauss_blur_3_rd6_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd6_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd6_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd6_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd6_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd6_select_out;
  dark_weights_normed_gauss_blur_3_rd6_select selector_dark_weights_normed_gauss_blur_3_rd6_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd6_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd6_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd6_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd6_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd6_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd6_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd6_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd6_select

  // selector_dark_weights_normed_gauss_blur_3_rd5_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd5_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd5_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd5_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd5_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd5_select_out;
  dark_weights_normed_gauss_blur_3_rd5_select selector_dark_weights_normed_gauss_blur_3_rd5_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd5_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd5_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd5_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd5_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd5_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd5_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd5_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd5_select

  // selector_fused_level_2_rd0_select
  logic [0:0] selector_fused_level_2_rd0_select_clk;
  logic [0:0] selector_fused_level_2_rd0_select_rst;
  logic [31:0] selector_fused_level_2_rd0_select_d0;
  logic [31:0] selector_fused_level_2_rd0_select_d1;
  logic [31:0] selector_fused_level_2_rd0_select_out;
  fused_level_2_rd0_select selector_fused_level_2_rd0_select(.clk(selector_fused_level_2_rd0_select_clk), .rst(selector_fused_level_2_rd0_select_rst), .d0(selector_fused_level_2_rd0_select_d0), .d1(selector_fused_level_2_rd0_select_d1), .out(selector_fused_level_2_rd0_select_out));
  assign selector_fused_level_2_rd0_select_clk = clk;
  assign selector_fused_level_2_rd0_select_rst = rst;
  // Bindings to selector_fused_level_2_rd0_select

  // Bindings to fused_level_2_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_2_update_0_read_dummy;

  // Bindings to dark_weights_normed_gauss_blur_3_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_weights_normed_gauss_blur_3_update_0_read_dummy;

  // selector_dark_weights_normed_gauss_blur_3_rd7_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd7_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd7_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd7_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd7_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd7_select_out;
  dark_weights_normed_gauss_blur_3_rd7_select selector_dark_weights_normed_gauss_blur_3_rd7_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd7_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd7_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd7_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd7_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd7_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd7_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd7_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd7_select

  // Bindings to dark_weights_normed_gauss_ds_2_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_normed_gauss_ds_2_update_0_write_wen;

  // selector_dark_weights_normed_gauss_blur_3_rd8_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd8_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd8_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd8_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd8_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd8_select_out;
  dark_weights_normed_gauss_blur_3_rd8_select selector_dark_weights_normed_gauss_blur_3_rd8_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd8_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd8_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd8_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd8_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd8_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd8_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd8_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd8_select

  // Bindings to dark_weights_normed_gauss_ds_2_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_normed_gauss_ds_2_update_0_write_wdata;

  // Bindings to dark_weights_normed_gauss_blur_3_update_0_read_rdata
    // wr_3
  assign dark_weights_normed_gauss_blur_3_update_0_read_rdata = rd_2;

  // Bindings to fused_level_2_update_0_read_rdata
    // wr_5
  assign fused_level_2_update_0_read_rdata = rd_4;



endmodule


module dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module final_merged_0_final_merged_0_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_final_merged_0_update_0_write_wen(output [0:0] final_merged_0_update_0_write_wen);

endmodule


module pyramid_synthetic_exposure_fusion_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_final_merged_0_update_0_write_wdata(output [31:0] final_merged_0_update_0_write_wdata);

endmodule


module in_wire_pyramid_synthetic_exposure_fusion_update_0_read_dummy(output [31:0] pyramid_synthetic_exposure_fusion_update_0_read_dummy);

endmodule


module out_wire_pyramid_synthetic_exposure_fusion_update_0_read_rdata(input [31:0] pyramid_synthetic_exposure_fusion_update_0_read_rdata);

endmodule


module final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98



endmodule


module in_wire_final_merged_1_update_0_write_wdata(output [31:0] final_merged_1_update_0_write_wdata);

endmodule


module in_wire_final_merged_1_update_0_write_wen(output [0:0] final_merged_1_update_0_write_wen);

endmodule


module in_wire_final_merged_0_update_0_read_dummy(output [31:0] final_merged_0_update_0_read_dummy);

endmodule


module out_wire_final_merged_0_update_0_read_rdata(input [31:0] final_merged_0_update_0_read_rdata);

endmodule


module final_merged_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_fused_level_1_update_0_write_wen(output [0:0] fused_level_1_update_0_write_wen);

endmodule


module in_wire_fused_level_1_update_0_write_wdata(output [31:0] fused_level_1_update_0_write_wdata);

endmodule


module fused_level_2_fused_level_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_fused_level_2_update_0_write_wen(output [0:0] fused_level_2_update_0_write_wen);

endmodule


module in_wire_fused_level_2_update_0_write_wdata(output [31:0] fused_level_2_update_0_write_wdata);

endmodule


module in_wire_final_merged_2_update_0_read_dummy(output [31:0] final_merged_2_update_0_read_dummy);

endmodule


module out_wire_final_merged_2_update_0_read_rdata(input [31:0] final_merged_2_update_0_read_rdata);

endmodule


module fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24



endmodule


module in_wire_fused_level_3_update_0_write_wen(output [0:0] fused_level_3_update_0_write_wen);

endmodule


module final_merged_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = ((-1 - d1) % 2 == 0 && 23 - d0 >= 0) ? ((12 - floord(2*d0, 4))) : 0;
    end
  end

endmodule


module in_wire_fused_level_3_update_0_write_wdata(output [31:0] fused_level_3_update_0_write_wdata);

endmodule


module bright_bright_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_108 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_108 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6



endmodule


module sr_buffer_32_1231(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 1231;

  reg [31:0] data [1230:0];

  reg [31:0] rdata_d;

  reg [10:0] waddr;

  wire [10:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_diff_1_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_279 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114



endmodule


module sr_buffer_32_278(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 278;

  reg [31:0] data [277:0];

  reg [31:0] rdata_d;

  reg [8:0] waddr;

  wire [8:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module bright_laplace_diff_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] fused_level_2_update_0_read_dummy, input [0:0] bright_laplace_diff_2_update_0_write_wen, input [31:0] bright_laplace_diff_2_update_0_write_wdata, output [31:0] fused_level_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to fused_level_2_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_2_update_0_read_dummy;

  // selector_fused_level_2_rd0_select
  logic [0:0] selector_fused_level_2_rd0_select_clk;
  logic [0:0] selector_fused_level_2_rd0_select_rst;
  logic [31:0] selector_fused_level_2_rd0_select_d0;
  logic [31:0] selector_fused_level_2_rd0_select_d1;
  logic [31:0] selector_fused_level_2_rd0_select_out;
  fused_level_2_rd0_select selector_fused_level_2_rd0_select(.clk(selector_fused_level_2_rd0_select_clk), .rst(selector_fused_level_2_rd0_select_rst), .d0(selector_fused_level_2_rd0_select_d0), .d1(selector_fused_level_2_rd0_select_d1), .out(selector_fused_level_2_rd0_select_out));
  assign selector_fused_level_2_rd0_select_clk = clk;
  assign selector_fused_level_2_rd0_select_rst = rst;
  // Bindings to selector_fused_level_2_rd0_select

  // bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1
  logic [0:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_done;
  bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1 bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1(.clk(bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_clk), .rst(bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_rst), .start(bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_start), .done(bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_done));
  assign bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_clk = clk;
  assign bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1

  // Bindings to bright_laplace_diff_2_update_0_write_wen
    // rd_0
  assign rd_0 = bright_laplace_diff_2_update_0_write_wen;

  // Bindings to bright_laplace_diff_2_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_laplace_diff_2_update_0_write_wdata;

  // Bindings to fused_level_2_update_0_read_rdata
    // wr_3
  assign fused_level_2_update_0_read_rdata = rd_2;



endmodule


module in_wire_bright_laplace_us_0_update_0_write_wdata(output [31:0] bright_laplace_us_0_update_0_write_wdata);

endmodule


module bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_laplace_us_0_update_0_write_wen(output [0:0] bright_laplace_us_0_update_0_write_wen);

endmodule


module bright_laplace_diff_0_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module bright_laplace_us_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_laplace_us_0_update_0_write_wen, input [31:0] bright_laplace_us_0_update_0_write_wdata, input [31:0] bright_laplace_diff_0_update_0_read_dummy, output [31:0] bright_laplace_diff_0_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to bright_laplace_us_0_update_0_write_wen
    // rd_0
  assign rd_0 = bright_laplace_us_0_update_0_write_wen;

  // selector_bright_laplace_diff_0_rd0_select
  logic [0:0] selector_bright_laplace_diff_0_rd0_select_clk;
  logic [0:0] selector_bright_laplace_diff_0_rd0_select_rst;
  logic [31:0] selector_bright_laplace_diff_0_rd0_select_d0;
  logic [31:0] selector_bright_laplace_diff_0_rd0_select_d1;
  logic [31:0] selector_bright_laplace_diff_0_rd0_select_out;
  bright_laplace_diff_0_rd0_select selector_bright_laplace_diff_0_rd0_select(.clk(selector_bright_laplace_diff_0_rd0_select_clk), .rst(selector_bright_laplace_diff_0_rd0_select_rst), .d0(selector_bright_laplace_diff_0_rd0_select_d0), .d1(selector_bright_laplace_diff_0_rd0_select_d1), .out(selector_bright_laplace_diff_0_rd0_select_out));
  assign selector_bright_laplace_diff_0_rd0_select_clk = clk;
  assign selector_bright_laplace_diff_0_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_diff_0_rd0_select

  // bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1
  logic [0:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_done;
  bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1 bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1(.clk(bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_clk), .rst(bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_rst), .start(bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_start), .done(bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_done));
  assign bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_clk = clk;
  assign bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1

  // Bindings to bright_laplace_us_0_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_laplace_us_0_update_0_write_wdata;

  // Bindings to bright_laplace_diff_0_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_laplace_diff_0_update_0_read_dummy;

  // Bindings to bright_laplace_diff_0_update_0_read_rdata
    // wr_3
  assign bright_laplace_diff_0_update_0_read_rdata = rd_2;



endmodule


module in_wire_bright_laplace_us_1_update_0_write_wen(output [0:0] bright_laplace_us_1_update_0_write_wen);

endmodule


module bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module bright_laplace_diff_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_laplace_us_1_update_0_write_wdata(output [31:0] bright_laplace_us_1_update_0_write_wdata);

endmodule


module bright_laplace_us_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_laplace_us_1_update_0_write_wen, output [31:0] bright_laplace_diff_1_update_0_read_rdata, input [31:0] bright_laplace_us_1_update_0_write_wdata, input [31:0] bright_laplace_diff_1_update_0_read_dummy);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to bright_laplace_us_1_update_0_write_wen
    // rd_0
  assign rd_0 = bright_laplace_us_1_update_0_write_wen;

  // Bindings to bright_laplace_diff_1_update_0_read_rdata
    // wr_3
  assign bright_laplace_diff_1_update_0_read_rdata = rd_2;

  // bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1
  logic [0:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_done;
  bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1 bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1(.clk(bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_clk), .rst(bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_rst), .start(bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_start), .done(bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_done));
  assign bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_clk = clk;
  assign bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1

  // selector_bright_laplace_diff_1_rd0_select
  logic [0:0] selector_bright_laplace_diff_1_rd0_select_clk;
  logic [0:0] selector_bright_laplace_diff_1_rd0_select_rst;
  logic [31:0] selector_bright_laplace_diff_1_rd0_select_d0;
  logic [31:0] selector_bright_laplace_diff_1_rd0_select_d1;
  logic [31:0] selector_bright_laplace_diff_1_rd0_select_out;
  bright_laplace_diff_1_rd0_select selector_bright_laplace_diff_1_rd0_select(.clk(selector_bright_laplace_diff_1_rd0_select_clk), .rst(selector_bright_laplace_diff_1_rd0_select_rst), .d0(selector_bright_laplace_diff_1_rd0_select_d0), .d1(selector_bright_laplace_diff_1_rd0_select_d1), .out(selector_bright_laplace_diff_1_rd0_select_out));
  assign selector_bright_laplace_diff_1_rd0_select_clk = clk;
  assign selector_bright_laplace_diff_1_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_diff_1_rd0_select

  // Bindings to bright_laplace_us_1_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_laplace_us_1_update_0_write_wdata;

  // Bindings to bright_laplace_diff_1_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_laplace_diff_1_update_0_read_dummy;



endmodule


module in_wire_bright_laplace_us_2_update_0_write_wen(output [0:0] bright_laplace_us_2_update_0_write_wen);

endmodule


module bright_laplace_diff_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_laplace_us_2_update_0_write_wdata(output [31:0] bright_laplace_us_2_update_0_write_wdata);

endmodule


module bright_laplace_us_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_laplace_us_2_update_0_write_wen, input [31:0] bright_laplace_us_2_update_0_write_wdata, input [31:0] bright_laplace_diff_2_update_0_read_dummy, output [31:0] bright_laplace_diff_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to bright_laplace_us_2_update_0_write_wen
    // rd_0
  assign rd_0 = bright_laplace_us_2_update_0_write_wen;

  // bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1
  logic [0:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_done;
  bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1 bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1(.clk(bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_clk), .rst(bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_rst), .start(bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_start), .done(bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_done));
  assign bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_clk = clk;
  assign bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1

  // selector_bright_laplace_diff_2_rd0_select
  logic [0:0] selector_bright_laplace_diff_2_rd0_select_clk;
  logic [0:0] selector_bright_laplace_diff_2_rd0_select_rst;
  logic [31:0] selector_bright_laplace_diff_2_rd0_select_d0;
  logic [31:0] selector_bright_laplace_diff_2_rd0_select_d1;
  logic [31:0] selector_bright_laplace_diff_2_rd0_select_out;
  bright_laplace_diff_2_rd0_select selector_bright_laplace_diff_2_rd0_select(.clk(selector_bright_laplace_diff_2_rd0_select_clk), .rst(selector_bright_laplace_diff_2_rd0_select_rst), .d0(selector_bright_laplace_diff_2_rd0_select_d0), .d1(selector_bright_laplace_diff_2_rd0_select_d1), .out(selector_bright_laplace_diff_2_rd0_select_out));
  assign selector_bright_laplace_diff_2_rd0_select_clk = clk;
  assign selector_bright_laplace_diff_2_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_diff_2_rd0_select

  // Bindings to bright_laplace_us_2_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_laplace_us_2_update_0_write_wdata;

  // Bindings to bright_laplace_diff_2_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_laplace_diff_2_update_0_read_dummy;

  // Bindings to bright_laplace_diff_2_update_0_read_rdata
    // wr_3
  assign bright_laplace_diff_2_update_0_read_rdata = rd_2;



endmodule


module in_wire_bright_weights_update_0_write_wen(output [0:0] bright_weights_update_0_write_wen);

endmodule


module bright_weights_bright_weights_update_0_write0_merged_banks_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_weights_update_0_write_wdata(output [31:0] bright_weights_update_0_write_wdata);

endmodule


module in_wire_bright_weights_normed_update_0_read_dummy(output [31:0] bright_weights_normed_update_0_read_dummy);

endmodule


module out_wire_bright_weights_normed_update_0_read_rdata(input [31:0] bright_weights_normed_update_0_read_rdata);

endmodule


module in_wire_weight_sums_update_0_read_dummy(output [31:0] weight_sums_update_0_read_dummy);

endmodule


module out_wire_weight_sums_update_0_read_rdata(input [31:0] weight_sums_update_0_read_rdata);

endmodule


module bright_weights(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_weights_update_0_write_wen, input [31:0] weight_sums_update_0_read_dummy, input [31:0] bright_weights_update_0_write_wdata, input [31:0] bright_weights_normed_update_0_read_dummy, output [31:0] bright_weights_normed_update_0_read_rdata, output [31:0] weight_sums_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // Bindings to bright_weights_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_update_0_write_wen;

  // bright_weights_bright_weights_update_0_write0_merged_banks_2
  logic [0:0] bright_weights_bright_weights_update_0_write0_merged_banks_2_clk;
  logic [0:0] bright_weights_bright_weights_update_0_write0_merged_banks_2_rst;
  logic [0:0] bright_weights_bright_weights_update_0_write0_merged_banks_2_start;
  logic [0:0] bright_weights_bright_weights_update_0_write0_merged_banks_2_done;
  bright_weights_bright_weights_update_0_write0_merged_banks_2 bright_weights_bright_weights_update_0_write0_merged_banks_2(.clk(bright_weights_bright_weights_update_0_write0_merged_banks_2_clk), .rst(bright_weights_bright_weights_update_0_write0_merged_banks_2_rst), .start(bright_weights_bright_weights_update_0_write0_merged_banks_2_start), .done(bright_weights_bright_weights_update_0_write0_merged_banks_2_done));
  assign bright_weights_bright_weights_update_0_write0_merged_banks_2_clk = clk;
  assign bright_weights_bright_weights_update_0_write0_merged_banks_2_rst = rst;
  // Bindings to bright_weights_bright_weights_update_0_write0_merged_banks_2

  // selector_weight_sums_rd0_select
  logic [0:0] selector_weight_sums_rd0_select_clk;
  logic [0:0] selector_weight_sums_rd0_select_rst;
  logic [31:0] selector_weight_sums_rd0_select_d0;
  logic [31:0] selector_weight_sums_rd0_select_d1;
  logic [31:0] selector_weight_sums_rd0_select_out;
  weight_sums_rd0_select selector_weight_sums_rd0_select(.clk(selector_weight_sums_rd0_select_clk), .rst(selector_weight_sums_rd0_select_rst), .d0(selector_weight_sums_rd0_select_d0), .d1(selector_weight_sums_rd0_select_d1), .out(selector_weight_sums_rd0_select_out));
  assign selector_weight_sums_rd0_select_clk = clk;
  assign selector_weight_sums_rd0_select_rst = rst;
  // Bindings to selector_weight_sums_rd0_select

  // selector_bright_weights_normed_rd0_select
  logic [0:0] selector_bright_weights_normed_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_rd0_select_out;
  bright_weights_normed_rd0_select selector_bright_weights_normed_rd0_select(.clk(selector_bright_weights_normed_rd0_select_clk), .rst(selector_bright_weights_normed_rd0_select_rst), .d0(selector_bright_weights_normed_rd0_select_d0), .d1(selector_bright_weights_normed_rd0_select_d1), .out(selector_bright_weights_normed_rd0_select_out));
  assign selector_bright_weights_normed_rd0_select_clk = clk;
  assign selector_bright_weights_normed_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_rd0_select

  // Bindings to weight_sums_update_0_read_dummy
    // rd_4
  assign rd_4 = weight_sums_update_0_read_dummy;

  // Bindings to bright_weights_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_update_0_write_wdata;

  // Bindings to bright_weights_normed_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_update_0_read_dummy;

  // Bindings to bright_weights_normed_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_update_0_read_rdata = rd_2;

  // Bindings to weight_sums_update_0_read_rdata
    // wr_5
  assign weight_sums_update_0_read_rdata = rd_4;



endmodule


module bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1231 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f314
  logic [0:0] f314_wen;
  logic [31:0] f314_wdata;
  logic [0:0] f314_clk;
  logic [0:0] f314_rst;
  logic [31:0] f314_rdata;
  sr_buffer_32_1 f314(.wen(f314_wen), .wdata(f314_wdata), .clk(f314_clk), .rst(f314_rst), .rdata(f314_rdata));
  assign f314_clk = clk;
  assign f314_rst = rst;
  // Bindings to f314

  // f316
  logic [0:0] f316_wen;
  logic [31:0] f316_wdata;
  logic [0:0] f316_clk;
  logic [0:0] f316_rst;
  logic [31:0] f316_rdata;
  sr_buffer_32_1 f316(.wen(f316_wen), .wdata(f316_wdata), .clk(f316_clk), .rst(f316_rst), .rdata(f316_rdata));
  assign f316_clk = clk;
  assign f316_rst = rst;
  // Bindings to f316

  // f318
  logic [0:0] f318_wen;
  logic [31:0] f318_wdata;
  logic [0:0] f318_clk;
  logic [0:0] f318_rst;
  logic [31:0] f318_rdata;
  sr_buffer_32_1 f318(.wen(f318_wen), .wdata(f318_wdata), .clk(f318_clk), .rst(f318_rst), .rdata(f318_rdata));
  assign f318_clk = clk;
  assign f318_rst = rst;
  // Bindings to f318

  // f320
  logic [0:0] f320_wen;
  logic [31:0] f320_wdata;
  logic [0:0] f320_clk;
  logic [0:0] f320_rst;
  logic [31:0] f320_rdata;
  sr_buffer_32_1 f320(.wen(f320_wen), .wdata(f320_wdata), .clk(f320_clk), .rst(f320_rst), .rdata(f320_rdata));
  assign f320_clk = clk;
  assign f320_rst = rst;
  // Bindings to f320

  // f322
  logic [0:0] f322_wen;
  logic [31:0] f322_wdata;
  logic [0:0] f322_clk;
  logic [0:0] f322_rst;
  logic [31:0] f322_rdata;
  sr_buffer_32_1 f322(.wen(f322_wen), .wdata(f322_wdata), .clk(f322_clk), .rst(f322_rst), .rdata(f322_rdata));
  assign f322_clk = clk;
  assign f322_rst = rst;
  // Bindings to f322

  // f324
  logic [0:0] f324_wen;
  logic [31:0] f324_wdata;
  logic [0:0] f324_clk;
  logic [0:0] f324_rst;
  logic [31:0] f324_rdata;
  sr_buffer_32_1 f324(.wen(f324_wen), .wdata(f324_wdata), .clk(f324_clk), .rst(f324_rst), .rdata(f324_rdata));
  assign f324_clk = clk;
  assign f324_rst = rst;
  // Bindings to f324

  // f326
  logic [0:0] f326_wen;
  logic [31:0] f326_wdata;
  logic [0:0] f326_clk;
  logic [0:0] f326_rst;
  logic [31:0] f326_rdata;
  sr_buffer_32_1 f326(.wen(f326_wen), .wdata(f326_wdata), .clk(f326_clk), .rst(f326_rst), .rdata(f326_rdata));
  assign f326_clk = clk;
  assign f326_rst = rst;
  // Bindings to f326

  // f328
  logic [0:0] f328_wen;
  logic [31:0] f328_wdata;
  logic [0:0] f328_clk;
  logic [0:0] f328_rst;
  logic [31:0] f328_rdata;
  sr_buffer_32_1 f328(.wen(f328_wen), .wdata(f328_wdata), .clk(f328_clk), .rst(f328_rst), .rdata(f328_rdata));
  assign f328_clk = clk;
  assign f328_rst = rst;
  // Bindings to f328

  // f330
  logic [0:0] f330_wen;
  logic [31:0] f330_wdata;
  logic [0:0] f330_clk;
  logic [0:0] f330_rst;
  logic [31:0] f330_rdata;
  sr_buffer_32_1 f330(.wen(f330_wen), .wdata(f330_wdata), .clk(f330_clk), .rst(f330_rst), .rdata(f330_rdata));
  assign f330_clk = clk;
  assign f330_rst = rst;
  // Bindings to f330

  // f332
  logic [0:0] f332_wen;
  logic [31:0] f332_wdata;
  logic [0:0] f332_clk;
  logic [0:0] f332_rst;
  logic [31:0] f332_rdata;
  sr_buffer_32_1 f332(.wen(f332_wen), .wdata(f332_wdata), .clk(f332_clk), .rst(f332_rst), .rdata(f332_rdata));
  assign f332_clk = clk;
  assign f332_rst = rst;
  // Bindings to f332

  // f334
  logic [0:0] f334_wen;
  logic [31:0] f334_wdata;
  logic [0:0] f334_clk;
  logic [0:0] f334_rst;
  logic [31:0] f334_rdata;
  sr_buffer_32_1 f334(.wen(f334_wen), .wdata(f334_wdata), .clk(f334_clk), .rst(f334_rst), .rdata(f334_rdata));
  assign f334_clk = clk;
  assign f334_rst = rst;
  // Bindings to f334

  // f336
  logic [0:0] f336_wen;
  logic [31:0] f336_wdata;
  logic [0:0] f336_clk;
  logic [0:0] f336_rst;
  logic [31:0] f336_rdata;
  sr_buffer_32_1 f336(.wen(f336_wen), .wdata(f336_wdata), .clk(f336_clk), .rst(f336_rst), .rdata(f336_rdata));
  assign f336_clk = clk;
  assign f336_rst = rst;
  // Bindings to f336

  // f338
  logic [0:0] f338_wen;
  logic [31:0] f338_wdata;
  logic [0:0] f338_clk;
  logic [0:0] f338_rst;
  logic [31:0] f338_rdata;
  sr_buffer_32_1 f338(.wen(f338_wen), .wdata(f338_wdata), .clk(f338_clk), .rst(f338_rst), .rdata(f338_rdata));
  assign f338_clk = clk;
  assign f338_rst = rst;
  // Bindings to f338

  // f340
  logic [0:0] f340_wen;
  logic [31:0] f340_wdata;
  logic [0:0] f340_clk;
  logic [0:0] f340_rst;
  logic [31:0] f340_rdata;
  sr_buffer_32_1 f340(.wen(f340_wen), .wdata(f340_wdata), .clk(f340_clk), .rst(f340_rst), .rdata(f340_rdata));
  assign f340_clk = clk;
  assign f340_rst = rst;
  // Bindings to f340

  // f342
  logic [0:0] f342_wen;
  logic [31:0] f342_wdata;
  logic [0:0] f342_clk;
  logic [0:0] f342_rst;
  logic [31:0] f342_rdata;
  sr_buffer_32_1 f342(.wen(f342_wen), .wdata(f342_wdata), .clk(f342_clk), .rst(f342_rst), .rdata(f342_rdata));
  assign f342_clk = clk;
  assign f342_rst = rst;
  // Bindings to f342

  // f344
  logic [0:0] f344_wen;
  logic [31:0] f344_wdata;
  logic [0:0] f344_clk;
  logic [0:0] f344_rst;
  logic [31:0] f344_rdata;
  sr_buffer_32_1 f344(.wen(f344_wen), .wdata(f344_wdata), .clk(f344_clk), .rst(f344_rst), .rdata(f344_rdata));
  assign f344_clk = clk;
  assign f344_rst = rst;
  // Bindings to f344

  // f346
  logic [0:0] f346_wen;
  logic [31:0] f346_wdata;
  logic [0:0] f346_clk;
  logic [0:0] f346_rst;
  logic [31:0] f346_rdata;
  sr_buffer_32_1 f346(.wen(f346_wen), .wdata(f346_wdata), .clk(f346_clk), .rst(f346_rst), .rdata(f346_rdata));
  assign f346_clk = clk;
  assign f346_rst = rst;
  // Bindings to f346

  // f348
  logic [0:0] f348_wen;
  logic [31:0] f348_wdata;
  logic [0:0] f348_clk;
  logic [0:0] f348_rst;
  logic [31:0] f348_rdata;
  sr_buffer_32_1 f348(.wen(f348_wen), .wdata(f348_wdata), .clk(f348_clk), .rst(f348_rst), .rdata(f348_rdata));
  assign f348_clk = clk;
  assign f348_rst = rst;
  // Bindings to f348

  // f350
  logic [0:0] f350_wen;
  logic [31:0] f350_wdata;
  logic [0:0] f350_clk;
  logic [0:0] f350_rst;
  logic [31:0] f350_rdata;
  sr_buffer_32_1 f350(.wen(f350_wen), .wdata(f350_wdata), .clk(f350_clk), .rst(f350_rst), .rdata(f350_rdata));
  assign f350_clk = clk;
  assign f350_rst = rst;
  // Bindings to f350

  // f352
  logic [0:0] f352_wen;
  logic [31:0] f352_wdata;
  logic [0:0] f352_clk;
  logic [0:0] f352_rst;
  logic [31:0] f352_rdata;
  sr_buffer_32_1 f352(.wen(f352_wen), .wdata(f352_wdata), .clk(f352_clk), .rst(f352_rst), .rdata(f352_rdata));
  assign f352_clk = clk;
  assign f352_rst = rst;
  // Bindings to f352

  // f354
  logic [0:0] f354_wen;
  logic [31:0] f354_wdata;
  logic [0:0] f354_clk;
  logic [0:0] f354_rst;
  logic [31:0] f354_rdata;
  sr_buffer_32_1 f354(.wen(f354_wen), .wdata(f354_wdata), .clk(f354_clk), .rst(f354_rst), .rdata(f354_rdata));
  assign f354_clk = clk;
  assign f354_rst = rst;
  // Bindings to f354

  // f356
  logic [0:0] f356_wen;
  logic [31:0] f356_wdata;
  logic [0:0] f356_clk;
  logic [0:0] f356_rst;
  logic [31:0] f356_rdata;
  sr_buffer_32_1 f356(.wen(f356_wen), .wdata(f356_wdata), .clk(f356_clk), .rst(f356_rst), .rdata(f356_rdata));
  assign f356_clk = clk;
  assign f356_rst = rst;
  // Bindings to f356

  // f358
  logic [0:0] f358_wen;
  logic [31:0] f358_wdata;
  logic [0:0] f358_clk;
  logic [0:0] f358_rst;
  logic [31:0] f358_rdata;
  sr_buffer_32_1 f358(.wen(f358_wen), .wdata(f358_wdata), .clk(f358_clk), .rst(f358_rst), .rdata(f358_rdata));
  assign f358_clk = clk;
  assign f358_rst = rst;
  // Bindings to f358

  // f360
  logic [0:0] f360_wen;
  logic [31:0] f360_wdata;
  logic [0:0] f360_clk;
  logic [0:0] f360_rst;
  logic [31:0] f360_rdata;
  sr_buffer_32_1 f360(.wen(f360_wen), .wdata(f360_wdata), .clk(f360_clk), .rst(f360_rst), .rdata(f360_rdata));
  assign f360_clk = clk;
  assign f360_rst = rst;
  // Bindings to f360

  // f362
  logic [0:0] f362_wen;
  logic [31:0] f362_wdata;
  logic [0:0] f362_clk;
  logic [0:0] f362_rst;
  logic [31:0] f362_rdata;
  sr_buffer_32_1 f362(.wen(f362_wen), .wdata(f362_wdata), .clk(f362_clk), .rst(f362_rst), .rdata(f362_rdata));
  assign f362_clk = clk;
  assign f362_rst = rst;
  // Bindings to f362

  // f364
  logic [0:0] f364_wen;
  logic [31:0] f364_wdata;
  logic [0:0] f364_clk;
  logic [0:0] f364_rst;
  logic [31:0] f364_rdata;
  sr_buffer_32_1 f364(.wen(f364_wen), .wdata(f364_wdata), .clk(f364_clk), .rst(f364_rst), .rdata(f364_rdata));
  assign f364_clk = clk;
  assign f364_rst = rst;
  // Bindings to f364

  // f366
  logic [0:0] f366_wen;
  logic [31:0] f366_wdata;
  logic [0:0] f366_clk;
  logic [0:0] f366_rst;
  logic [31:0] f366_rdata;
  sr_buffer_32_1 f366(.wen(f366_wen), .wdata(f366_wdata), .clk(f366_clk), .rst(f366_rst), .rdata(f366_rdata));
  assign f366_clk = clk;
  assign f366_rst = rst;
  // Bindings to f366

  // f368
  logic [0:0] f368_wen;
  logic [31:0] f368_wdata;
  logic [0:0] f368_clk;
  logic [0:0] f368_rst;
  logic [31:0] f368_rdata;
  sr_buffer_32_1 f368(.wen(f368_wen), .wdata(f368_wdata), .clk(f368_clk), .rst(f368_rst), .rdata(f368_rdata));
  assign f368_clk = clk;
  assign f368_rst = rst;
  // Bindings to f368

  // f370
  logic [0:0] f370_wen;
  logic [31:0] f370_wdata;
  logic [0:0] f370_clk;
  logic [0:0] f370_rst;
  logic [31:0] f370_rdata;
  sr_buffer_32_1 f370(.wen(f370_wen), .wdata(f370_wdata), .clk(f370_clk), .rst(f370_rst), .rdata(f370_rdata));
  assign f370_clk = clk;
  assign f370_rst = rst;
  // Bindings to f370

  // f372
  logic [0:0] f372_wen;
  logic [31:0] f372_wdata;
  logic [0:0] f372_clk;
  logic [0:0] f372_rst;
  logic [31:0] f372_rdata;
  sr_buffer_32_1 f372(.wen(f372_wen), .wdata(f372_wdata), .clk(f372_clk), .rst(f372_rst), .rdata(f372_rdata));
  assign f372_clk = clk;
  assign f372_rst = rst;
  // Bindings to f372

  // f374
  logic [0:0] f374_wen;
  logic [31:0] f374_wdata;
  logic [0:0] f374_clk;
  logic [0:0] f374_rst;
  logic [31:0] f374_rdata;
  sr_buffer_32_1 f374(.wen(f374_wen), .wdata(f374_wdata), .clk(f374_clk), .rst(f374_rst), .rdata(f374_rdata));
  assign f374_clk = clk;
  assign f374_rst = rst;
  // Bindings to f374

  // f376
  logic [0:0] f376_wen;
  logic [31:0] f376_wdata;
  logic [0:0] f376_clk;
  logic [0:0] f376_rst;
  logic [31:0] f376_rdata;
  sr_buffer_32_1 f376(.wen(f376_wen), .wdata(f376_wdata), .clk(f376_clk), .rst(f376_rst), .rdata(f376_rdata));
  assign f376_clk = clk;
  assign f376_rst = rst;
  // Bindings to f376

  // f378
  logic [0:0] f378_wen;
  logic [31:0] f378_wdata;
  logic [0:0] f378_clk;
  logic [0:0] f378_rst;
  logic [31:0] f378_rdata;
  sr_buffer_32_1 f378(.wen(f378_wen), .wdata(f378_wdata), .clk(f378_clk), .rst(f378_rst), .rdata(f378_rdata));
  assign f378_clk = clk;
  assign f378_rst = rst;
  // Bindings to f378

  // f380
  logic [0:0] f380_wen;
  logic [31:0] f380_wdata;
  logic [0:0] f380_clk;
  logic [0:0] f380_rst;
  logic [31:0] f380_rdata;
  sr_buffer_32_1 f380(.wen(f380_wen), .wdata(f380_wdata), .clk(f380_clk), .rst(f380_rst), .rdata(f380_rdata));
  assign f380_clk = clk;
  assign f380_rst = rst;
  // Bindings to f380

  // f382
  logic [0:0] f382_wen;
  logic [31:0] f382_wdata;
  logic [0:0] f382_clk;
  logic [0:0] f382_rst;
  logic [31:0] f382_rdata;
  sr_buffer_32_1 f382(.wen(f382_wen), .wdata(f382_wdata), .clk(f382_clk), .rst(f382_rst), .rdata(f382_rdata));
  assign f382_clk = clk;
  assign f382_rst = rst;
  // Bindings to f382

  // f384
  logic [0:0] f384_wen;
  logic [31:0] f384_wdata;
  logic [0:0] f384_clk;
  logic [0:0] f384_rst;
  logic [31:0] f384_rdata;
  sr_buffer_32_1 f384(.wen(f384_wen), .wdata(f384_wdata), .clk(f384_clk), .rst(f384_rst), .rdata(f384_rdata));
  assign f384_clk = clk;
  assign f384_rst = rst;
  // Bindings to f384

  // f386
  logic [0:0] f386_wen;
  logic [31:0] f386_wdata;
  logic [0:0] f386_clk;
  logic [0:0] f386_rst;
  logic [31:0] f386_rdata;
  sr_buffer_32_1 f386(.wen(f386_wen), .wdata(f386_wdata), .clk(f386_clk), .rst(f386_rst), .rdata(f386_rdata));
  assign f386_clk = clk;
  assign f386_rst = rst;
  // Bindings to f386

  // f388
  logic [0:0] f388_wen;
  logic [31:0] f388_wdata;
  logic [0:0] f388_clk;
  logic [0:0] f388_rst;
  logic [31:0] f388_rdata;
  sr_buffer_32_1 f388(.wen(f388_wen), .wdata(f388_wdata), .clk(f388_clk), .rst(f388_rst), .rdata(f388_rdata));
  assign f388_clk = clk;
  assign f388_rst = rst;
  // Bindings to f388

  // f390
  logic [0:0] f390_wen;
  logic [31:0] f390_wdata;
  logic [0:0] f390_clk;
  logic [0:0] f390_rst;
  logic [31:0] f390_rdata;
  sr_buffer_32_1 f390(.wen(f390_wen), .wdata(f390_wdata), .clk(f390_clk), .rst(f390_rst), .rdata(f390_rdata));
  assign f390_clk = clk;
  assign f390_rst = rst;
  // Bindings to f390

  // f392
  logic [0:0] f392_wen;
  logic [31:0] f392_wdata;
  logic [0:0] f392_clk;
  logic [0:0] f392_rst;
  logic [31:0] f392_rdata;
  sr_buffer_32_1 f392(.wen(f392_wen), .wdata(f392_wdata), .clk(f392_clk), .rst(f392_rst), .rdata(f392_rdata));
  assign f392_clk = clk;
  assign f392_rst = rst;
  // Bindings to f392

  // f394
  logic [0:0] f394_wen;
  logic [31:0] f394_wdata;
  logic [0:0] f394_clk;
  logic [0:0] f394_rst;
  logic [31:0] f394_rdata;
  sr_buffer_32_1 f394(.wen(f394_wen), .wdata(f394_wdata), .clk(f394_clk), .rst(f394_rst), .rdata(f394_rdata));
  assign f394_clk = clk;
  assign f394_rst = rst;
  // Bindings to f394

  // f396
  logic [0:0] f396_wen;
  logic [31:0] f396_wdata;
  logic [0:0] f396_clk;
  logic [0:0] f396_rst;
  logic [31:0] f396_rdata;
  sr_buffer_32_1 f396(.wen(f396_wen), .wdata(f396_wdata), .clk(f396_clk), .rst(f396_rst), .rdata(f396_rdata));
  assign f396_clk = clk;
  assign f396_rst = rst;
  // Bindings to f396

  // f398
  logic [0:0] f398_wen;
  logic [31:0] f398_wdata;
  logic [0:0] f398_clk;
  logic [0:0] f398_rst;
  logic [31:0] f398_rdata;
  sr_buffer_32_1 f398(.wen(f398_wen), .wdata(f398_wdata), .clk(f398_clk), .rst(f398_rst), .rdata(f398_rdata));
  assign f398_clk = clk;
  assign f398_rst = rst;
  // Bindings to f398

  // f400
  logic [0:0] f400_wen;
  logic [31:0] f400_wdata;
  logic [0:0] f400_clk;
  logic [0:0] f400_rst;
  logic [31:0] f400_rdata;
  sr_buffer_32_1 f400(.wen(f400_wen), .wdata(f400_wdata), .clk(f400_clk), .rst(f400_rst), .rdata(f400_rdata));
  assign f400_clk = clk;
  assign f400_rst = rst;
  // Bindings to f400

  // f402
  logic [0:0] f402_wen;
  logic [31:0] f402_wdata;
  logic [0:0] f402_clk;
  logic [0:0] f402_rst;
  logic [31:0] f402_rdata;
  sr_buffer_32_1 f402(.wen(f402_wen), .wdata(f402_wdata), .clk(f402_clk), .rst(f402_rst), .rdata(f402_rdata));
  assign f402_clk = clk;
  assign f402_rst = rst;
  // Bindings to f402

  // f404
  logic [0:0] f404_wen;
  logic [31:0] f404_wdata;
  logic [0:0] f404_clk;
  logic [0:0] f404_rst;
  logic [31:0] f404_rdata;
  sr_buffer_32_1 f404(.wen(f404_wen), .wdata(f404_wdata), .clk(f404_clk), .rst(f404_rst), .rdata(f404_rdata));
  assign f404_clk = clk;
  assign f404_rst = rst;
  // Bindings to f404

  // f406
  logic [0:0] f406_wen;
  logic [31:0] f406_wdata;
  logic [0:0] f406_clk;
  logic [0:0] f406_rst;
  logic [31:0] f406_rdata;
  sr_buffer_32_1 f406(.wen(f406_wen), .wdata(f406_wdata), .clk(f406_clk), .rst(f406_rst), .rdata(f406_rdata));
  assign f406_clk = clk;
  assign f406_rst = rst;
  // Bindings to f406

  // f408
  logic [0:0] f408_wen;
  logic [31:0] f408_wdata;
  logic [0:0] f408_clk;
  logic [0:0] f408_rst;
  logic [31:0] f408_rdata;
  sr_buffer_32_1 f408(.wen(f408_wen), .wdata(f408_wdata), .clk(f408_clk), .rst(f408_rst), .rdata(f408_rdata));
  assign f408_clk = clk;
  assign f408_rst = rst;
  // Bindings to f408

  // f410
  logic [0:0] f410_wen;
  logic [31:0] f410_wdata;
  logic [0:0] f410_clk;
  logic [0:0] f410_rst;
  logic [31:0] f410_rdata;
  sr_buffer_32_1 f410(.wen(f410_wen), .wdata(f410_wdata), .clk(f410_clk), .rst(f410_rst), .rdata(f410_rdata));
  assign f410_clk = clk;
  assign f410_rst = rst;
  // Bindings to f410

  // f412
  logic [0:0] f412_wen;
  logic [31:0] f412_wdata;
  logic [0:0] f412_clk;
  logic [0:0] f412_rst;
  logic [31:0] f412_rdata;
  sr_buffer_32_1 f412(.wen(f412_wen), .wdata(f412_wdata), .clk(f412_clk), .rst(f412_rst), .rdata(f412_rdata));
  assign f412_clk = clk;
  assign f412_rst = rst;
  // Bindings to f412

  // f414
  logic [0:0] f414_wen;
  logic [31:0] f414_wdata;
  logic [0:0] f414_clk;
  logic [0:0] f414_rst;
  logic [31:0] f414_rdata;
  sr_buffer_32_1 f414(.wen(f414_wen), .wdata(f414_wdata), .clk(f414_clk), .rst(f414_rst), .rdata(f414_rdata));
  assign f414_clk = clk;
  assign f414_rst = rst;
  // Bindings to f414

  // f416
  logic [0:0] f416_wen;
  logic [31:0] f416_wdata;
  logic [0:0] f416_clk;
  logic [0:0] f416_rst;
  logic [31:0] f416_rdata;
  sr_buffer_32_1 f416(.wen(f416_wen), .wdata(f416_wdata), .clk(f416_clk), .rst(f416_rst), .rdata(f416_rdata));
  assign f416_clk = clk;
  assign f416_rst = rst;
  // Bindings to f416

  // f418
  logic [0:0] f418_wen;
  logic [31:0] f418_wdata;
  logic [0:0] f418_clk;
  logic [0:0] f418_rst;
  logic [31:0] f418_rdata;
  sr_buffer_32_1 f418(.wen(f418_wen), .wdata(f418_wdata), .clk(f418_clk), .rst(f418_rst), .rdata(f418_rdata));
  assign f418_clk = clk;
  assign f418_rst = rst;
  // Bindings to f418

  // f420
  logic [0:0] f420_wen;
  logic [31:0] f420_wdata;
  logic [0:0] f420_clk;
  logic [0:0] f420_rst;
  logic [31:0] f420_rdata;
  sr_buffer_32_1 f420(.wen(f420_wen), .wdata(f420_wdata), .clk(f420_clk), .rst(f420_rst), .rdata(f420_rdata));
  assign f420_clk = clk;
  assign f420_rst = rst;
  // Bindings to f420

  // f422
  logic [0:0] f422_wen;
  logic [31:0] f422_wdata;
  logic [0:0] f422_clk;
  logic [0:0] f422_rst;
  logic [31:0] f422_rdata;
  sr_buffer_32_1 f422(.wen(f422_wen), .wdata(f422_wdata), .clk(f422_clk), .rst(f422_rst), .rdata(f422_rdata));
  assign f422_clk = clk;
  assign f422_rst = rst;
  // Bindings to f422

  // f424
  logic [0:0] f424_wen;
  logic [31:0] f424_wdata;
  logic [0:0] f424_clk;
  logic [0:0] f424_rst;
  logic [31:0] f424_rdata;
  sr_buffer_32_1 f424(.wen(f424_wen), .wdata(f424_wdata), .clk(f424_clk), .rst(f424_rst), .rdata(f424_rdata));
  assign f424_clk = clk;
  assign f424_rst = rst;
  // Bindings to f424

  // f426
  logic [0:0] f426_wen;
  logic [31:0] f426_wdata;
  logic [0:0] f426_clk;
  logic [0:0] f426_rst;
  logic [31:0] f426_rdata;
  sr_buffer_32_1 f426(.wen(f426_wen), .wdata(f426_wdata), .clk(f426_clk), .rst(f426_rst), .rdata(f426_rdata));
  assign f426_clk = clk;
  assign f426_rst = rst;
  // Bindings to f426

  // f428
  logic [0:0] f428_wen;
  logic [31:0] f428_wdata;
  logic [0:0] f428_clk;
  logic [0:0] f428_rst;
  logic [31:0] f428_rdata;
  sr_buffer_32_1 f428(.wen(f428_wen), .wdata(f428_wdata), .clk(f428_clk), .rst(f428_rst), .rdata(f428_rdata));
  assign f428_clk = clk;
  assign f428_rst = rst;
  // Bindings to f428

  // f430
  logic [0:0] f430_wen;
  logic [31:0] f430_wdata;
  logic [0:0] f430_clk;
  logic [0:0] f430_rst;
  logic [31:0] f430_rdata;
  sr_buffer_32_1 f430(.wen(f430_wen), .wdata(f430_wdata), .clk(f430_clk), .rst(f430_rst), .rdata(f430_rdata));
  assign f430_clk = clk;
  assign f430_rst = rst;
  // Bindings to f430

  // f432
  logic [0:0] f432_wen;
  logic [31:0] f432_wdata;
  logic [0:0] f432_clk;
  logic [0:0] f432_rst;
  logic [31:0] f432_rdata;
  sr_buffer_32_1 f432(.wen(f432_wen), .wdata(f432_wdata), .clk(f432_clk), .rst(f432_rst), .rdata(f432_rdata));
  assign f432_clk = clk;
  assign f432_rst = rst;
  // Bindings to f432

  // f434
  logic [0:0] f434_wen;
  logic [31:0] f434_wdata;
  logic [0:0] f434_clk;
  logic [0:0] f434_rst;
  logic [31:0] f434_rdata;
  sr_buffer_32_1 f434(.wen(f434_wen), .wdata(f434_wdata), .clk(f434_clk), .rst(f434_rst), .rdata(f434_rdata));
  assign f434_clk = clk;
  assign f434_rst = rst;
  // Bindings to f434

  // f436
  logic [0:0] f436_wen;
  logic [31:0] f436_wdata;
  logic [0:0] f436_clk;
  logic [0:0] f436_rst;
  logic [31:0] f436_rdata;
  sr_buffer_32_1 f436(.wen(f436_wen), .wdata(f436_wdata), .clk(f436_clk), .rst(f436_rst), .rdata(f436_rdata));
  assign f436_clk = clk;
  assign f436_rst = rst;
  // Bindings to f436

  // f438
  logic [0:0] f438_wen;
  logic [31:0] f438_wdata;
  logic [0:0] f438_clk;
  logic [0:0] f438_rst;
  logic [31:0] f438_rdata;
  sr_buffer_32_1 f438(.wen(f438_wen), .wdata(f438_wdata), .clk(f438_clk), .rst(f438_rst), .rdata(f438_rdata));
  assign f438_clk = clk;
  assign f438_rst = rst;
  // Bindings to f438

  // f440
  logic [0:0] f440_wen;
  logic [31:0] f440_wdata;
  logic [0:0] f440_clk;
  logic [0:0] f440_rst;
  logic [31:0] f440_rdata;
  sr_buffer_32_1 f440(.wen(f440_wen), .wdata(f440_wdata), .clk(f440_clk), .rst(f440_rst), .rdata(f440_rdata));
  assign f440_clk = clk;
  assign f440_rst = rst;
  // Bindings to f440

  // f442
  logic [0:0] f442_wen;
  logic [31:0] f442_wdata;
  logic [0:0] f442_clk;
  logic [0:0] f442_rst;
  logic [31:0] f442_rdata;
  sr_buffer_32_1 f442(.wen(f442_wen), .wdata(f442_wdata), .clk(f442_clk), .rst(f442_rst), .rdata(f442_rdata));
  assign f442_clk = clk;
  assign f442_rst = rst;
  // Bindings to f442

  // f444
  logic [0:0] f444_wen;
  logic [31:0] f444_wdata;
  logic [0:0] f444_clk;
  logic [0:0] f444_rst;
  logic [31:0] f444_rdata;
  sr_buffer_32_1 f444(.wen(f444_wen), .wdata(f444_wdata), .clk(f444_clk), .rst(f444_rst), .rdata(f444_rdata));
  assign f444_clk = clk;
  assign f444_rst = rst;
  // Bindings to f444

  // f446
  logic [0:0] f446_wen;
  logic [31:0] f446_wdata;
  logic [0:0] f446_clk;
  logic [0:0] f446_rst;
  logic [31:0] f446_rdata;
  sr_buffer_32_1 f446(.wen(f446_wen), .wdata(f446_wdata), .clk(f446_clk), .rst(f446_rst), .rdata(f446_rdata));
  assign f446_clk = clk;
  assign f446_rst = rst;
  // Bindings to f446

  // f448
  logic [0:0] f448_wen;
  logic [31:0] f448_wdata;
  logic [0:0] f448_clk;
  logic [0:0] f448_rst;
  logic [31:0] f448_rdata;
  sr_buffer_32_1 f448(.wen(f448_wen), .wdata(f448_wdata), .clk(f448_clk), .rst(f448_rst), .rdata(f448_rdata));
  assign f448_clk = clk;
  assign f448_rst = rst;
  // Bindings to f448

  // f450
  logic [0:0] f450_wen;
  logic [31:0] f450_wdata;
  logic [0:0] f450_clk;
  logic [0:0] f450_rst;
  logic [31:0] f450_rdata;
  sr_buffer_32_1 f450(.wen(f450_wen), .wdata(f450_wdata), .clk(f450_clk), .rst(f450_rst), .rdata(f450_rdata));
  assign f450_clk = clk;
  assign f450_rst = rst;
  // Bindings to f450

  // f452
  logic [0:0] f452_wen;
  logic [31:0] f452_wdata;
  logic [0:0] f452_clk;
  logic [0:0] f452_rst;
  logic [31:0] f452_rdata;
  sr_buffer_32_1 f452(.wen(f452_wen), .wdata(f452_wdata), .clk(f452_clk), .rst(f452_rst), .rdata(f452_rdata));
  assign f452_clk = clk;
  assign f452_rst = rst;
  // Bindings to f452

  // f454
  logic [0:0] f454_wen;
  logic [31:0] f454_wdata;
  logic [0:0] f454_clk;
  logic [0:0] f454_rst;
  logic [31:0] f454_rdata;
  sr_buffer_32_1 f454(.wen(f454_wen), .wdata(f454_wdata), .clk(f454_clk), .rst(f454_rst), .rdata(f454_rdata));
  assign f454_clk = clk;
  assign f454_rst = rst;
  // Bindings to f454

  // f456
  logic [0:0] f456_wen;
  logic [31:0] f456_wdata;
  logic [0:0] f456_clk;
  logic [0:0] f456_rst;
  logic [31:0] f456_rdata;
  sr_buffer_32_1 f456(.wen(f456_wen), .wdata(f456_wdata), .clk(f456_clk), .rst(f456_rst), .rdata(f456_rdata));
  assign f456_clk = clk;
  assign f456_rst = rst;
  // Bindings to f456

  // f458
  logic [0:0] f458_wen;
  logic [31:0] f458_wdata;
  logic [0:0] f458_clk;
  logic [0:0] f458_rst;
  logic [31:0] f458_rdata;
  sr_buffer_32_1 f458(.wen(f458_wen), .wdata(f458_wdata), .clk(f458_clk), .rst(f458_rst), .rdata(f458_rdata));
  assign f458_clk = clk;
  assign f458_rst = rst;
  // Bindings to f458

  // f460
  logic [0:0] f460_wen;
  logic [31:0] f460_wdata;
  logic [0:0] f460_clk;
  logic [0:0] f460_rst;
  logic [31:0] f460_rdata;
  sr_buffer_32_1 f460(.wen(f460_wen), .wdata(f460_wdata), .clk(f460_clk), .rst(f460_rst), .rdata(f460_rdata));
  assign f460_clk = clk;
  assign f460_rst = rst;
  // Bindings to f460

  // f462
  logic [0:0] f462_wen;
  logic [31:0] f462_wdata;
  logic [0:0] f462_clk;
  logic [0:0] f462_rst;
  logic [31:0] f462_rdata;
  sr_buffer_32_1 f462(.wen(f462_wen), .wdata(f462_wdata), .clk(f462_clk), .rst(f462_rst), .rdata(f462_rdata));
  assign f462_clk = clk;
  assign f462_rst = rst;
  // Bindings to f462

  // f464
  logic [0:0] f464_wen;
  logic [31:0] f464_wdata;
  logic [0:0] f464_clk;
  logic [0:0] f464_rst;
  logic [31:0] f464_rdata;
  sr_buffer_32_1 f464(.wen(f464_wen), .wdata(f464_wdata), .clk(f464_clk), .rst(f464_rst), .rdata(f464_rdata));
  assign f464_clk = clk;
  assign f464_rst = rst;
  // Bindings to f464

  // f466
  logic [0:0] f466_wen;
  logic [31:0] f466_wdata;
  logic [0:0] f466_clk;
  logic [0:0] f466_rst;
  logic [31:0] f466_rdata;
  sr_buffer_32_1 f466(.wen(f466_wen), .wdata(f466_wdata), .clk(f466_clk), .rst(f466_rst), .rdata(f466_rdata));
  assign f466_clk = clk;
  assign f466_rst = rst;
  // Bindings to f466

  // f468
  logic [0:0] f468_wen;
  logic [31:0] f468_wdata;
  logic [0:0] f468_clk;
  logic [0:0] f468_rst;
  logic [31:0] f468_rdata;
  sr_buffer_32_1 f468(.wen(f468_wen), .wdata(f468_wdata), .clk(f468_clk), .rst(f468_rst), .rdata(f468_rdata));
  assign f468_clk = clk;
  assign f468_rst = rst;
  // Bindings to f468

  // f470
  logic [0:0] f470_wen;
  logic [31:0] f470_wdata;
  logic [0:0] f470_clk;
  logic [0:0] f470_rst;
  logic [31:0] f470_rdata;
  sr_buffer_32_1 f470(.wen(f470_wen), .wdata(f470_wdata), .clk(f470_clk), .rst(f470_rst), .rdata(f470_rdata));
  assign f470_clk = clk;
  assign f470_rst = rst;
  // Bindings to f470

  // f472
  logic [0:0] f472_wen;
  logic [31:0] f472_wdata;
  logic [0:0] f472_clk;
  logic [0:0] f472_rst;
  logic [31:0] f472_rdata;
  sr_buffer_32_1 f472(.wen(f472_wen), .wdata(f472_wdata), .clk(f472_clk), .rst(f472_rst), .rdata(f472_rdata));
  assign f472_clk = clk;
  assign f472_rst = rst;
  // Bindings to f472

  // f474
  logic [0:0] f474_wen;
  logic [31:0] f474_wdata;
  logic [0:0] f474_clk;
  logic [0:0] f474_rst;
  logic [31:0] f474_rdata;
  sr_buffer_32_1 f474(.wen(f474_wen), .wdata(f474_wdata), .clk(f474_clk), .rst(f474_rst), .rdata(f474_rdata));
  assign f474_clk = clk;
  assign f474_rst = rst;
  // Bindings to f474

  // f476
  logic [0:0] f476_wen;
  logic [31:0] f476_wdata;
  logic [0:0] f476_clk;
  logic [0:0] f476_rst;
  logic [31:0] f476_rdata;
  sr_buffer_32_1 f476(.wen(f476_wen), .wdata(f476_wdata), .clk(f476_clk), .rst(f476_rst), .rdata(f476_rdata));
  assign f476_clk = clk;
  assign f476_rst = rst;
  // Bindings to f476

  // f478
  logic [0:0] f478_wen;
  logic [31:0] f478_wdata;
  logic [0:0] f478_clk;
  logic [0:0] f478_rst;
  logic [31:0] f478_rdata;
  sr_buffer_32_1 f478(.wen(f478_wen), .wdata(f478_wdata), .clk(f478_clk), .rst(f478_rst), .rdata(f478_rdata));
  assign f478_clk = clk;
  assign f478_rst = rst;
  // Bindings to f478

  // f480
  logic [0:0] f480_wen;
  logic [31:0] f480_wdata;
  logic [0:0] f480_clk;
  logic [0:0] f480_rst;
  logic [31:0] f480_rdata;
  sr_buffer_32_1 f480(.wen(f480_wen), .wdata(f480_wdata), .clk(f480_clk), .rst(f480_rst), .rdata(f480_rdata));
  assign f480_clk = clk;
  assign f480_rst = rst;
  // Bindings to f480

  // f482
  logic [0:0] f482_wen;
  logic [31:0] f482_wdata;
  logic [0:0] f482_clk;
  logic [0:0] f482_rst;
  logic [31:0] f482_rdata;
  sr_buffer_32_1 f482(.wen(f482_wen), .wdata(f482_wdata), .clk(f482_clk), .rst(f482_rst), .rdata(f482_rdata));
  assign f482_clk = clk;
  assign f482_rst = rst;
  // Bindings to f482

  // f484
  logic [0:0] f484_wen;
  logic [31:0] f484_wdata;
  logic [0:0] f484_clk;
  logic [0:0] f484_rst;
  logic [31:0] f484_rdata;
  sr_buffer_32_1 f484(.wen(f484_wen), .wdata(f484_wdata), .clk(f484_clk), .rst(f484_rst), .rdata(f484_rdata));
  assign f484_clk = clk;
  assign f484_rst = rst;
  // Bindings to f484

  // f486
  logic [0:0] f486_wen;
  logic [31:0] f486_wdata;
  logic [0:0] f486_clk;
  logic [0:0] f486_rst;
  logic [31:0] f486_rdata;
  sr_buffer_32_1 f486(.wen(f486_wen), .wdata(f486_wdata), .clk(f486_clk), .rst(f486_rst), .rdata(f486_rdata));
  assign f486_clk = clk;
  assign f486_rst = rst;
  // Bindings to f486

  // f488
  logic [0:0] f488_wen;
  logic [31:0] f488_wdata;
  logic [0:0] f488_clk;
  logic [0:0] f488_rst;
  logic [31:0] f488_rdata;
  sr_buffer_32_1 f488(.wen(f488_wen), .wdata(f488_wdata), .clk(f488_clk), .rst(f488_rst), .rdata(f488_rdata));
  assign f488_clk = clk;
  assign f488_rst = rst;
  // Bindings to f488

  // f490
  logic [0:0] f490_wen;
  logic [31:0] f490_wdata;
  logic [0:0] f490_clk;
  logic [0:0] f490_rst;
  logic [31:0] f490_rdata;
  sr_buffer_32_1 f490(.wen(f490_wen), .wdata(f490_wdata), .clk(f490_clk), .rst(f490_rst), .rdata(f490_rdata));
  assign f490_clk = clk;
  assign f490_rst = rst;
  // Bindings to f490

  // f492
  logic [0:0] f492_wen;
  logic [31:0] f492_wdata;
  logic [0:0] f492_clk;
  logic [0:0] f492_rst;
  logic [31:0] f492_rdata;
  sr_buffer_32_1 f492(.wen(f492_wen), .wdata(f492_wdata), .clk(f492_clk), .rst(f492_rst), .rdata(f492_rdata));
  assign f492_clk = clk;
  assign f492_rst = rst;
  // Bindings to f492

  // f494
  logic [0:0] f494_wen;
  logic [31:0] f494_wdata;
  logic [0:0] f494_clk;
  logic [0:0] f494_rst;
  logic [31:0] f494_rdata;
  sr_buffer_32_1 f494(.wen(f494_wen), .wdata(f494_wdata), .clk(f494_clk), .rst(f494_rst), .rdata(f494_rdata));
  assign f494_clk = clk;
  assign f494_rst = rst;
  // Bindings to f494

  // f496
  logic [0:0] f496_wen;
  logic [31:0] f496_wdata;
  logic [0:0] f496_clk;
  logic [0:0] f496_rst;
  logic [31:0] f496_rdata;
  sr_buffer_32_1 f496(.wen(f496_wen), .wdata(f496_wdata), .clk(f496_clk), .rst(f496_rst), .rdata(f496_rdata));
  assign f496_clk = clk;
  assign f496_rst = rst;
  // Bindings to f496

  // f498
  logic [0:0] f498_wen;
  logic [31:0] f498_wdata;
  logic [0:0] f498_clk;
  logic [0:0] f498_rst;
  logic [31:0] f498_rdata;
  sr_buffer_32_1 f498(.wen(f498_wen), .wdata(f498_wdata), .clk(f498_clk), .rst(f498_rst), .rdata(f498_rdata));
  assign f498_clk = clk;
  assign f498_rst = rst;
  // Bindings to f498

  // f500
  logic [0:0] f500_wen;
  logic [31:0] f500_wdata;
  logic [0:0] f500_clk;
  logic [0:0] f500_rst;
  logic [31:0] f500_rdata;
  sr_buffer_32_1 f500(.wen(f500_wen), .wdata(f500_wdata), .clk(f500_clk), .rst(f500_rst), .rdata(f500_rdata));
  assign f500_clk = clk;
  assign f500_rst = rst;
  // Bindings to f500

  // f502
  logic [0:0] f502_wen;
  logic [31:0] f502_wdata;
  logic [0:0] f502_clk;
  logic [0:0] f502_rst;
  logic [31:0] f502_rdata;
  sr_buffer_32_1 f502(.wen(f502_wen), .wdata(f502_wdata), .clk(f502_clk), .rst(f502_rst), .rdata(f502_rdata));
  assign f502_clk = clk;
  assign f502_rst = rst;
  // Bindings to f502

  // f504
  logic [0:0] f504_wen;
  logic [31:0] f504_wdata;
  logic [0:0] f504_clk;
  logic [0:0] f504_rst;
  logic [31:0] f504_rdata;
  sr_buffer_32_1 f504(.wen(f504_wen), .wdata(f504_wdata), .clk(f504_clk), .rst(f504_rst), .rdata(f504_rdata));
  assign f504_clk = clk;
  assign f504_rst = rst;
  // Bindings to f504

  // f506
  logic [0:0] f506_wen;
  logic [31:0] f506_wdata;
  logic [0:0] f506_clk;
  logic [0:0] f506_rst;
  logic [31:0] f506_rdata;
  sr_buffer_32_1 f506(.wen(f506_wen), .wdata(f506_wdata), .clk(f506_clk), .rst(f506_rst), .rdata(f506_rdata));
  assign f506_clk = clk;
  assign f506_rst = rst;
  // Bindings to f506

  // f508
  logic [0:0] f508_wen;
  logic [31:0] f508_wdata;
  logic [0:0] f508_clk;
  logic [0:0] f508_rst;
  logic [31:0] f508_rdata;
  sr_buffer_32_1 f508(.wen(f508_wen), .wdata(f508_wdata), .clk(f508_clk), .rst(f508_rst), .rdata(f508_rdata));
  assign f508_clk = clk;
  assign f508_rst = rst;
  // Bindings to f508

  // f510
  logic [0:0] f510_wen;
  logic [31:0] f510_wdata;
  logic [0:0] f510_clk;
  logic [0:0] f510_rst;
  logic [31:0] f510_rdata;
  sr_buffer_32_1 f510(.wen(f510_wen), .wdata(f510_wdata), .clk(f510_clk), .rst(f510_rst), .rdata(f510_rdata));
  assign f510_clk = clk;
  assign f510_rst = rst;
  // Bindings to f510

  // f512
  logic [0:0] f512_wen;
  logic [31:0] f512_wdata;
  logic [0:0] f512_clk;
  logic [0:0] f512_rst;
  logic [31:0] f512_rdata;
  sr_buffer_32_1 f512(.wen(f512_wen), .wdata(f512_wdata), .clk(f512_clk), .rst(f512_rst), .rdata(f512_rdata));
  assign f512_clk = clk;
  assign f512_rst = rst;
  // Bindings to f512

  // f514
  logic [0:0] f514_wen;
  logic [31:0] f514_wdata;
  logic [0:0] f514_clk;
  logic [0:0] f514_rst;
  logic [31:0] f514_rdata;
  sr_buffer_32_1 f514(.wen(f514_wen), .wdata(f514_wdata), .clk(f514_clk), .rst(f514_rst), .rdata(f514_rdata));
  assign f514_clk = clk;
  assign f514_rst = rst;
  // Bindings to f514

  // f516
  logic [0:0] f516_wen;
  logic [31:0] f516_wdata;
  logic [0:0] f516_clk;
  logic [0:0] f516_rst;
  logic [31:0] f516_rdata;
  sr_buffer_32_1 f516(.wen(f516_wen), .wdata(f516_wdata), .clk(f516_clk), .rst(f516_rst), .rdata(f516_rdata));
  assign f516_clk = clk;
  assign f516_rst = rst;
  // Bindings to f516

  // f518
  logic [0:0] f518_wen;
  logic [31:0] f518_wdata;
  logic [0:0] f518_clk;
  logic [0:0] f518_rst;
  logic [31:0] f518_rdata;
  sr_buffer_32_1 f518(.wen(f518_wen), .wdata(f518_wdata), .clk(f518_clk), .rst(f518_rst), .rdata(f518_rdata));
  assign f518_clk = clk;
  assign f518_rst = rst;
  // Bindings to f518

  // f520
  logic [0:0] f520_wen;
  logic [31:0] f520_wdata;
  logic [0:0] f520_clk;
  logic [0:0] f520_rst;
  logic [31:0] f520_rdata;
  sr_buffer_32_1 f520(.wen(f520_wen), .wdata(f520_wdata), .clk(f520_clk), .rst(f520_rst), .rdata(f520_rdata));
  assign f520_clk = clk;
  assign f520_rst = rst;
  // Bindings to f520

  // f522
  logic [0:0] f522_wen;
  logic [31:0] f522_wdata;
  logic [0:0] f522_clk;
  logic [0:0] f522_rst;
  logic [31:0] f522_rdata;
  sr_buffer_32_1 f522(.wen(f522_wen), .wdata(f522_wdata), .clk(f522_clk), .rst(f522_rst), .rdata(f522_rdata));
  assign f522_clk = clk;
  assign f522_rst = rst;
  // Bindings to f522

  // f524
  logic [0:0] f524_wen;
  logic [31:0] f524_wdata;
  logic [0:0] f524_clk;
  logic [0:0] f524_rst;
  logic [31:0] f524_rdata;
  sr_buffer_32_1 f524(.wen(f524_wen), .wdata(f524_wdata), .clk(f524_clk), .rst(f524_rst), .rdata(f524_rdata));
  assign f524_clk = clk;
  assign f524_rst = rst;
  // Bindings to f524

  // f526
  logic [0:0] f526_wen;
  logic [31:0] f526_wdata;
  logic [0:0] f526_clk;
  logic [0:0] f526_rst;
  logic [31:0] f526_rdata;
  sr_buffer_32_1 f526(.wen(f526_wen), .wdata(f526_wdata), .clk(f526_clk), .rst(f526_rst), .rdata(f526_rdata));
  assign f526_clk = clk;
  assign f526_rst = rst;
  // Bindings to f526

  // f528
  logic [0:0] f528_wen;
  logic [31:0] f528_wdata;
  logic [0:0] f528_clk;
  logic [0:0] f528_rst;
  logic [31:0] f528_rdata;
  sr_buffer_32_1 f528(.wen(f528_wen), .wdata(f528_wdata), .clk(f528_clk), .rst(f528_rst), .rdata(f528_rdata));
  assign f528_clk = clk;
  assign f528_rst = rst;
  // Bindings to f528

  // f530
  logic [0:0] f530_wen;
  logic [31:0] f530_wdata;
  logic [0:0] f530_clk;
  logic [0:0] f530_rst;
  logic [31:0] f530_rdata;
  sr_buffer_32_1 f530(.wen(f530_wen), .wdata(f530_wdata), .clk(f530_clk), .rst(f530_rst), .rdata(f530_rdata));
  assign f530_clk = clk;
  assign f530_rst = rst;
  // Bindings to f530

  // f532
  logic [0:0] f532_wen;
  logic [31:0] f532_wdata;
  logic [0:0] f532_clk;
  logic [0:0] f532_rst;
  logic [31:0] f532_rdata;
  sr_buffer_32_1 f532(.wen(f532_wen), .wdata(f532_wdata), .clk(f532_clk), .rst(f532_rst), .rdata(f532_rdata));
  assign f532_clk = clk;
  assign f532_rst = rst;
  // Bindings to f532

  // f534
  logic [0:0] f534_wen;
  logic [31:0] f534_wdata;
  logic [0:0] f534_clk;
  logic [0:0] f534_rst;
  logic [31:0] f534_rdata;
  sr_buffer_32_1 f534(.wen(f534_wen), .wdata(f534_wdata), .clk(f534_clk), .rst(f534_rst), .rdata(f534_rdata));
  assign f534_clk = clk;
  assign f534_rst = rst;
  // Bindings to f534

  // f536
  logic [0:0] f536_wen;
  logic [31:0] f536_wdata;
  logic [0:0] f536_clk;
  logic [0:0] f536_rst;
  logic [31:0] f536_rdata;
  sr_buffer_32_1 f536(.wen(f536_wen), .wdata(f536_wdata), .clk(f536_clk), .rst(f536_rst), .rdata(f536_rdata));
  assign f536_clk = clk;
  assign f536_rst = rst;
  // Bindings to f536

  // f538
  logic [0:0] f538_wen;
  logic [31:0] f538_wdata;
  logic [0:0] f538_clk;
  logic [0:0] f538_rst;
  logic [31:0] f538_rdata;
  sr_buffer_32_1 f538(.wen(f538_wen), .wdata(f538_wdata), .clk(f538_clk), .rst(f538_rst), .rdata(f538_rdata));
  assign f538_clk = clk;
  assign f538_rst = rst;
  // Bindings to f538

  // f540
  logic [0:0] f540_wen;
  logic [31:0] f540_wdata;
  logic [0:0] f540_clk;
  logic [0:0] f540_rst;
  logic [31:0] f540_rdata;
  sr_buffer_32_1 f540(.wen(f540_wen), .wdata(f540_wdata), .clk(f540_clk), .rst(f540_rst), .rdata(f540_rdata));
  assign f540_clk = clk;
  assign f540_rst = rst;
  // Bindings to f540

  // f542
  logic [0:0] f542_wen;
  logic [31:0] f542_wdata;
  logic [0:0] f542_clk;
  logic [0:0] f542_rst;
  logic [31:0] f542_rdata;
  sr_buffer_32_1 f542(.wen(f542_wen), .wdata(f542_wdata), .clk(f542_clk), .rst(f542_rst), .rdata(f542_rdata));
  assign f542_clk = clk;
  assign f542_rst = rst;
  // Bindings to f542

  // f544
  logic [0:0] f544_wen;
  logic [31:0] f544_wdata;
  logic [0:0] f544_clk;
  logic [0:0] f544_rst;
  logic [31:0] f544_rdata;
  sr_buffer_32_1 f544(.wen(f544_wen), .wdata(f544_wdata), .clk(f544_clk), .rst(f544_rst), .rdata(f544_rdata));
  assign f544_clk = clk;
  assign f544_rst = rst;
  // Bindings to f544

  // f546
  logic [0:0] f546_wen;
  logic [31:0] f546_wdata;
  logic [0:0] f546_clk;
  logic [0:0] f546_rst;
  logic [31:0] f546_rdata;
  sr_buffer_32_1 f546(.wen(f546_wen), .wdata(f546_wdata), .clk(f546_clk), .rst(f546_rst), .rdata(f546_rdata));
  assign f546_clk = clk;
  assign f546_rst = rst;
  // Bindings to f546

  // f548
  logic [0:0] f548_wen;
  logic [31:0] f548_wdata;
  logic [0:0] f548_clk;
  logic [0:0] f548_rst;
  logic [31:0] f548_rdata;
  sr_buffer_32_1 f548(.wen(f548_wen), .wdata(f548_wdata), .clk(f548_clk), .rst(f548_rst), .rdata(f548_rdata));
  assign f548_clk = clk;
  assign f548_rst = rst;
  // Bindings to f548

  // f550
  logic [0:0] f550_wen;
  logic [31:0] f550_wdata;
  logic [0:0] f550_clk;
  logic [0:0] f550_rst;
  logic [31:0] f550_rdata;
  sr_buffer_32_1 f550(.wen(f550_wen), .wdata(f550_wdata), .clk(f550_clk), .rst(f550_rst), .rdata(f550_rdata));
  assign f550_clk = clk;
  assign f550_rst = rst;
  // Bindings to f550

  // f552
  logic [0:0] f552_wen;
  logic [31:0] f552_wdata;
  logic [0:0] f552_clk;
  logic [0:0] f552_rst;
  logic [31:0] f552_rdata;
  sr_buffer_32_1 f552(.wen(f552_wen), .wdata(f552_wdata), .clk(f552_clk), .rst(f552_rst), .rdata(f552_rdata));
  assign f552_clk = clk;
  assign f552_rst = rst;
  // Bindings to f552

  // f554
  logic [0:0] f554_wen;
  logic [31:0] f554_wdata;
  logic [0:0] f554_clk;
  logic [0:0] f554_rst;
  logic [31:0] f554_rdata;
  sr_buffer_32_1 f554(.wen(f554_wen), .wdata(f554_wdata), .clk(f554_clk), .rst(f554_rst), .rdata(f554_rdata));
  assign f554_clk = clk;
  assign f554_rst = rst;
  // Bindings to f554

  // f556
  logic [0:0] f556_wen;
  logic [31:0] f556_wdata;
  logic [0:0] f556_clk;
  logic [0:0] f556_rst;
  logic [31:0] f556_rdata;
  sr_buffer_32_1 f556(.wen(f556_wen), .wdata(f556_wdata), .clk(f556_clk), .rst(f556_rst), .rdata(f556_rdata));
  assign f556_clk = clk;
  assign f556_rst = rst;
  // Bindings to f556

  // f558
  logic [0:0] f558_wen;
  logic [31:0] f558_wdata;
  logic [0:0] f558_clk;
  logic [0:0] f558_rst;
  logic [31:0] f558_rdata;
  sr_buffer_32_1 f558(.wen(f558_wen), .wdata(f558_wdata), .clk(f558_clk), .rst(f558_rst), .rdata(f558_rdata));
  assign f558_clk = clk;
  assign f558_rst = rst;
  // Bindings to f558

  // f560
  logic [0:0] f560_wen;
  logic [31:0] f560_wdata;
  logic [0:0] f560_clk;
  logic [0:0] f560_rst;
  logic [31:0] f560_rdata;
  sr_buffer_32_1 f560(.wen(f560_wen), .wdata(f560_wdata), .clk(f560_clk), .rst(f560_rst), .rdata(f560_rdata));
  assign f560_clk = clk;
  assign f560_rst = rst;
  // Bindings to f560

  // f562
  logic [0:0] f562_wen;
  logic [31:0] f562_wdata;
  logic [0:0] f562_clk;
  logic [0:0] f562_rst;
  logic [31:0] f562_rdata;
  sr_buffer_32_1 f562(.wen(f562_wen), .wdata(f562_wdata), .clk(f562_clk), .rst(f562_rst), .rdata(f562_rdata));
  assign f562_clk = clk;
  assign f562_rst = rst;
  // Bindings to f562

  // f564
  logic [0:0] f564_wen;
  logic [31:0] f564_wdata;
  logic [0:0] f564_clk;
  logic [0:0] f564_rst;
  logic [31:0] f564_rdata;
  sr_buffer_32_1 f564(.wen(f564_wen), .wdata(f564_wdata), .clk(f564_clk), .rst(f564_rst), .rdata(f564_rdata));
  assign f564_clk = clk;
  assign f564_rst = rst;
  // Bindings to f564

  // f566
  logic [0:0] f566_wen;
  logic [31:0] f566_wdata;
  logic [0:0] f566_clk;
  logic [0:0] f566_rst;
  logic [31:0] f566_rdata;
  sr_buffer_32_1 f566(.wen(f566_wen), .wdata(f566_wdata), .clk(f566_clk), .rst(f566_rst), .rdata(f566_rdata));
  assign f566_clk = clk;
  assign f566_rst = rst;
  // Bindings to f566

  // f568
  logic [0:0] f568_wen;
  logic [31:0] f568_wdata;
  logic [0:0] f568_clk;
  logic [0:0] f568_rst;
  logic [31:0] f568_rdata;
  sr_buffer_32_1 f568(.wen(f568_wen), .wdata(f568_wdata), .clk(f568_clk), .rst(f568_rst), .rdata(f568_rdata));
  assign f568_clk = clk;
  assign f568_rst = rst;
  // Bindings to f568

  // f570
  logic [0:0] f570_wen;
  logic [31:0] f570_wdata;
  logic [0:0] f570_clk;
  logic [0:0] f570_rst;
  logic [31:0] f570_rdata;
  sr_buffer_32_1 f570(.wen(f570_wen), .wdata(f570_wdata), .clk(f570_clk), .rst(f570_rst), .rdata(f570_rdata));
  assign f570_clk = clk;
  assign f570_rst = rst;
  // Bindings to f570

  // f572
  logic [0:0] f572_wen;
  logic [31:0] f572_wdata;
  logic [0:0] f572_clk;
  logic [0:0] f572_rst;
  logic [31:0] f572_rdata;
  sr_buffer_32_1 f572(.wen(f572_wen), .wdata(f572_wdata), .clk(f572_clk), .rst(f572_rst), .rdata(f572_rdata));
  assign f572_clk = clk;
  assign f572_rst = rst;
  // Bindings to f572

  // f574
  logic [0:0] f574_wen;
  logic [31:0] f574_wdata;
  logic [0:0] f574_clk;
  logic [0:0] f574_rst;
  logic [31:0] f574_rdata;
  sr_buffer_32_1 f574(.wen(f574_wen), .wdata(f574_wdata), .clk(f574_clk), .rst(f574_rst), .rdata(f574_rdata));
  assign f574_clk = clk;
  assign f574_rst = rst;
  // Bindings to f574

  // f576
  logic [0:0] f576_wen;
  logic [31:0] f576_wdata;
  logic [0:0] f576_clk;
  logic [0:0] f576_rst;
  logic [31:0] f576_rdata;
  sr_buffer_32_1 f576(.wen(f576_wen), .wdata(f576_wdata), .clk(f576_clk), .rst(f576_rst), .rdata(f576_rdata));
  assign f576_clk = clk;
  assign f576_rst = rst;
  // Bindings to f576

  // f578
  logic [0:0] f578_wen;
  logic [31:0] f578_wdata;
  logic [0:0] f578_clk;
  logic [0:0] f578_rst;
  logic [31:0] f578_rdata;
  sr_buffer_32_1 f578(.wen(f578_wen), .wdata(f578_wdata), .clk(f578_clk), .rst(f578_rst), .rdata(f578_rdata));
  assign f578_clk = clk;
  assign f578_rst = rst;
  // Bindings to f578

  // f580
  logic [0:0] f580_wen;
  logic [31:0] f580_wdata;
  logic [0:0] f580_clk;
  logic [0:0] f580_rst;
  logic [31:0] f580_rdata;
  sr_buffer_32_1 f580(.wen(f580_wen), .wdata(f580_wdata), .clk(f580_clk), .rst(f580_rst), .rdata(f580_rdata));
  assign f580_clk = clk;
  assign f580_rst = rst;
  // Bindings to f580

  // f582
  logic [0:0] f582_wen;
  logic [31:0] f582_wdata;
  logic [0:0] f582_clk;
  logic [0:0] f582_rst;
  logic [31:0] f582_rdata;
  sr_buffer_32_1 f582(.wen(f582_wen), .wdata(f582_wdata), .clk(f582_clk), .rst(f582_rst), .rdata(f582_rdata));
  assign f582_clk = clk;
  assign f582_rst = rst;
  // Bindings to f582

  // f584
  logic [0:0] f584_wen;
  logic [31:0] f584_wdata;
  logic [0:0] f584_clk;
  logic [0:0] f584_rst;
  logic [31:0] f584_rdata;
  sr_buffer_32_1 f584(.wen(f584_wen), .wdata(f584_wdata), .clk(f584_clk), .rst(f584_rst), .rdata(f584_rdata));
  assign f584_clk = clk;
  assign f584_rst = rst;
  // Bindings to f584

  // f586
  logic [0:0] f586_wen;
  logic [31:0] f586_wdata;
  logic [0:0] f586_clk;
  logic [0:0] f586_rst;
  logic [31:0] f586_rdata;
  sr_buffer_32_1 f586(.wen(f586_wen), .wdata(f586_wdata), .clk(f586_clk), .rst(f586_rst), .rdata(f586_rdata));
  assign f586_clk = clk;
  assign f586_rst = rst;
  // Bindings to f586

  // f588
  logic [0:0] f588_wen;
  logic [31:0] f588_wdata;
  logic [0:0] f588_clk;
  logic [0:0] f588_rst;
  logic [31:0] f588_rdata;
  sr_buffer_32_1 f588(.wen(f588_wen), .wdata(f588_wdata), .clk(f588_clk), .rst(f588_rst), .rdata(f588_rdata));
  assign f588_clk = clk;
  assign f588_rst = rst;
  // Bindings to f588

  // f590
  logic [0:0] f590_wen;
  logic [31:0] f590_wdata;
  logic [0:0] f590_clk;
  logic [0:0] f590_rst;
  logic [31:0] f590_rdata;
  sr_buffer_32_1 f590(.wen(f590_wen), .wdata(f590_wdata), .clk(f590_clk), .rst(f590_rst), .rdata(f590_rdata));
  assign f590_clk = clk;
  assign f590_rst = rst;
  // Bindings to f590

  // f592
  logic [0:0] f592_wen;
  logic [31:0] f592_wdata;
  logic [0:0] f592_clk;
  logic [0:0] f592_rst;
  logic [31:0] f592_rdata;
  sr_buffer_32_1 f592(.wen(f592_wen), .wdata(f592_wdata), .clk(f592_clk), .rst(f592_rst), .rdata(f592_rdata));
  assign f592_clk = clk;
  assign f592_rst = rst;
  // Bindings to f592

  // f594
  logic [0:0] f594_wen;
  logic [31:0] f594_wdata;
  logic [0:0] f594_clk;
  logic [0:0] f594_rst;
  logic [31:0] f594_rdata;
  sr_buffer_32_1 f594(.wen(f594_wen), .wdata(f594_wdata), .clk(f594_clk), .rst(f594_rst), .rdata(f594_rdata));
  assign f594_clk = clk;
  assign f594_rst = rst;
  // Bindings to f594

  // f596
  logic [0:0] f596_wen;
  logic [31:0] f596_wdata;
  logic [0:0] f596_clk;
  logic [0:0] f596_rst;
  logic [31:0] f596_rdata;
  sr_buffer_32_1 f596(.wen(f596_wen), .wdata(f596_wdata), .clk(f596_clk), .rst(f596_rst), .rdata(f596_rdata));
  assign f596_clk = clk;
  assign f596_rst = rst;
  // Bindings to f596

  // f598
  logic [0:0] f598_wen;
  logic [31:0] f598_wdata;
  logic [0:0] f598_clk;
  logic [0:0] f598_rst;
  logic [31:0] f598_rdata;
  sr_buffer_32_1 f598(.wen(f598_wen), .wdata(f598_wdata), .clk(f598_clk), .rst(f598_rst), .rdata(f598_rdata));
  assign f598_clk = clk;
  assign f598_rst = rst;
  // Bindings to f598

  // f600
  logic [0:0] f600_wen;
  logic [31:0] f600_wdata;
  logic [0:0] f600_clk;
  logic [0:0] f600_rst;
  logic [31:0] f600_rdata;
  sr_buffer_32_1 f600(.wen(f600_wen), .wdata(f600_wdata), .clk(f600_clk), .rst(f600_rst), .rdata(f600_rdata));
  assign f600_clk = clk;
  assign f600_rst = rst;
  // Bindings to f600

  // f602
  logic [0:0] f602_wen;
  logic [31:0] f602_wdata;
  logic [0:0] f602_clk;
  logic [0:0] f602_rst;
  logic [31:0] f602_rdata;
  sr_buffer_32_1 f602(.wen(f602_wen), .wdata(f602_wdata), .clk(f602_clk), .rst(f602_rst), .rdata(f602_rdata));
  assign f602_clk = clk;
  assign f602_rst = rst;
  // Bindings to f602

  // f604
  logic [0:0] f604_wen;
  logic [31:0] f604_wdata;
  logic [0:0] f604_clk;
  logic [0:0] f604_rst;
  logic [31:0] f604_rdata;
  sr_buffer_32_1 f604(.wen(f604_wen), .wdata(f604_wdata), .clk(f604_clk), .rst(f604_rst), .rdata(f604_rdata));
  assign f604_clk = clk;
  assign f604_rst = rst;
  // Bindings to f604

  // f606
  logic [0:0] f606_wen;
  logic [31:0] f606_wdata;
  logic [0:0] f606_clk;
  logic [0:0] f606_rst;
  logic [31:0] f606_rdata;
  sr_buffer_32_1 f606(.wen(f606_wen), .wdata(f606_wdata), .clk(f606_clk), .rst(f606_rst), .rdata(f606_rdata));
  assign f606_clk = clk;
  assign f606_rst = rst;
  // Bindings to f606

  // f608
  logic [0:0] f608_wen;
  logic [31:0] f608_wdata;
  logic [0:0] f608_clk;
  logic [0:0] f608_rst;
  logic [31:0] f608_rdata;
  sr_buffer_32_1 f608(.wen(f608_wen), .wdata(f608_wdata), .clk(f608_clk), .rst(f608_rst), .rdata(f608_rdata));
  assign f608_clk = clk;
  assign f608_rst = rst;
  // Bindings to f608

  // f610
  logic [0:0] f610_wen;
  logic [31:0] f610_wdata;
  logic [0:0] f610_clk;
  logic [0:0] f610_rst;
  logic [31:0] f610_rdata;
  sr_buffer_32_1 f610(.wen(f610_wen), .wdata(f610_wdata), .clk(f610_clk), .rst(f610_rst), .rdata(f610_rdata));
  assign f610_clk = clk;
  assign f610_rst = rst;
  // Bindings to f610

  // f612
  logic [0:0] f612_wen;
  logic [31:0] f612_wdata;
  logic [0:0] f612_clk;
  logic [0:0] f612_rst;
  logic [31:0] f612_rdata;
  sr_buffer_32_1 f612(.wen(f612_wen), .wdata(f612_wdata), .clk(f612_clk), .rst(f612_rst), .rdata(f612_rdata));
  assign f612_clk = clk;
  assign f612_rst = rst;
  // Bindings to f612

  // f614
  logic [0:0] f614_wen;
  logic [31:0] f614_wdata;
  logic [0:0] f614_clk;
  logic [0:0] f614_rst;
  logic [31:0] f614_rdata;
  sr_buffer_32_1 f614(.wen(f614_wen), .wdata(f614_wdata), .clk(f614_clk), .rst(f614_rst), .rdata(f614_rdata));
  assign f614_clk = clk;
  assign f614_rst = rst;
  // Bindings to f614

  // f616
  logic [0:0] f616_wen;
  logic [31:0] f616_wdata;
  logic [0:0] f616_clk;
  logic [0:0] f616_rst;
  logic [31:0] f616_rdata;
  sr_buffer_32_1 f616(.wen(f616_wen), .wdata(f616_wdata), .clk(f616_clk), .rst(f616_rst), .rdata(f616_rdata));
  assign f616_clk = clk;
  assign f616_rst = rst;
  // Bindings to f616

  // f618
  logic [0:0] f618_wen;
  logic [31:0] f618_wdata;
  logic [0:0] f618_clk;
  logic [0:0] f618_rst;
  logic [31:0] f618_rdata;
  sr_buffer_32_1 f618(.wen(f618_wen), .wdata(f618_wdata), .clk(f618_clk), .rst(f618_rst), .rdata(f618_rdata));
  assign f618_clk = clk;
  assign f618_rst = rst;
  // Bindings to f618

  // f620
  logic [0:0] f620_wen;
  logic [31:0] f620_wdata;
  logic [0:0] f620_clk;
  logic [0:0] f620_rst;
  logic [31:0] f620_rdata;
  sr_buffer_32_1 f620(.wen(f620_wen), .wdata(f620_wdata), .clk(f620_clk), .rst(f620_rst), .rdata(f620_rdata));
  assign f620_clk = clk;
  assign f620_rst = rst;
  // Bindings to f620

  // f622
  logic [0:0] f622_wen;
  logic [31:0] f622_wdata;
  logic [0:0] f622_clk;
  logic [0:0] f622_rst;
  logic [31:0] f622_rdata;
  sr_buffer_32_1 f622(.wen(f622_wen), .wdata(f622_wdata), .clk(f622_clk), .rst(f622_rst), .rdata(f622_rdata));
  assign f622_clk = clk;
  assign f622_rst = rst;
  // Bindings to f622

  // f624
  logic [0:0] f624_wen;
  logic [31:0] f624_wdata;
  logic [0:0] f624_clk;
  logic [0:0] f624_rst;
  logic [31:0] f624_rdata;
  sr_buffer_32_1 f624(.wen(f624_wen), .wdata(f624_wdata), .clk(f624_clk), .rst(f624_rst), .rdata(f624_rdata));
  assign f624_clk = clk;
  assign f624_rst = rst;
  // Bindings to f624

  // f626
  logic [0:0] f626_wen;
  logic [31:0] f626_wdata;
  logic [0:0] f626_clk;
  logic [0:0] f626_rst;
  logic [31:0] f626_rdata;
  sr_buffer_32_1 f626(.wen(f626_wen), .wdata(f626_wdata), .clk(f626_clk), .rst(f626_rst), .rdata(f626_rdata));
  assign f626_clk = clk;
  assign f626_rst = rst;
  // Bindings to f626

  // f628
  logic [0:0] f628_wen;
  logic [31:0] f628_wdata;
  logic [0:0] f628_clk;
  logic [0:0] f628_rst;
  logic [31:0] f628_rdata;
  sr_buffer_32_1 f628(.wen(f628_wen), .wdata(f628_wdata), .clk(f628_clk), .rst(f628_rst), .rdata(f628_rdata));
  assign f628_clk = clk;
  assign f628_rst = rst;
  // Bindings to f628

  // f630
  logic [0:0] f630_wen;
  logic [31:0] f630_wdata;
  logic [0:0] f630_clk;
  logic [0:0] f630_rst;
  logic [31:0] f630_rdata;
  sr_buffer_32_1 f630(.wen(f630_wen), .wdata(f630_wdata), .clk(f630_clk), .rst(f630_rst), .rdata(f630_rdata));
  assign f630_clk = clk;
  assign f630_rst = rst;
  // Bindings to f630

  // f632
  logic [0:0] f632_wen;
  logic [31:0] f632_wdata;
  logic [0:0] f632_clk;
  logic [0:0] f632_rst;
  logic [31:0] f632_rdata;
  sr_buffer_32_1 f632(.wen(f632_wen), .wdata(f632_wdata), .clk(f632_clk), .rst(f632_rst), .rdata(f632_rdata));
  assign f632_clk = clk;
  assign f632_rst = rst;
  // Bindings to f632

  // f634
  logic [0:0] f634_wen;
  logic [31:0] f634_wdata;
  logic [0:0] f634_clk;
  logic [0:0] f634_rst;
  logic [31:0] f634_rdata;
  sr_buffer_32_1 f634(.wen(f634_wen), .wdata(f634_wdata), .clk(f634_clk), .rst(f634_rst), .rdata(f634_rdata));
  assign f634_clk = clk;
  assign f634_rst = rst;
  // Bindings to f634

  // f636
  logic [0:0] f636_wen;
  logic [31:0] f636_wdata;
  logic [0:0] f636_clk;
  logic [0:0] f636_rst;
  logic [31:0] f636_rdata;
  sr_buffer_32_1 f636(.wen(f636_wen), .wdata(f636_wdata), .clk(f636_clk), .rst(f636_rst), .rdata(f636_rdata));
  assign f636_clk = clk;
  assign f636_rst = rst;
  // Bindings to f636

  // f638
  logic [0:0] f638_wen;
  logic [31:0] f638_wdata;
  logic [0:0] f638_clk;
  logic [0:0] f638_rst;
  logic [31:0] f638_rdata;
  sr_buffer_32_1 f638(.wen(f638_wen), .wdata(f638_wdata), .clk(f638_clk), .rst(f638_rst), .rdata(f638_rdata));
  assign f638_clk = clk;
  assign f638_rst = rst;
  // Bindings to f638

  // f640
  logic [0:0] f640_wen;
  logic [31:0] f640_wdata;
  logic [0:0] f640_clk;
  logic [0:0] f640_rst;
  logic [31:0] f640_rdata;
  sr_buffer_32_1 f640(.wen(f640_wen), .wdata(f640_wdata), .clk(f640_clk), .rst(f640_rst), .rdata(f640_rdata));
  assign f640_clk = clk;
  assign f640_rst = rst;
  // Bindings to f640

  // f642
  logic [0:0] f642_wen;
  logic [31:0] f642_wdata;
  logic [0:0] f642_clk;
  logic [0:0] f642_rst;
  logic [31:0] f642_rdata;
  sr_buffer_32_1 f642(.wen(f642_wen), .wdata(f642_wdata), .clk(f642_clk), .rst(f642_rst), .rdata(f642_rdata));
  assign f642_clk = clk;
  assign f642_rst = rst;
  // Bindings to f642

  // f644
  logic [0:0] f644_wen;
  logic [31:0] f644_wdata;
  logic [0:0] f644_clk;
  logic [0:0] f644_rst;
  logic [31:0] f644_rdata;
  sr_buffer_32_1 f644(.wen(f644_wen), .wdata(f644_wdata), .clk(f644_clk), .rst(f644_rst), .rdata(f644_rdata));
  assign f644_clk = clk;
  assign f644_rst = rst;
  // Bindings to f644

  // f646
  logic [0:0] f646_wen;
  logic [31:0] f646_wdata;
  logic [0:0] f646_clk;
  logic [0:0] f646_rst;
  logic [31:0] f646_rdata;
  sr_buffer_32_1 f646(.wen(f646_wen), .wdata(f646_wdata), .clk(f646_clk), .rst(f646_rst), .rdata(f646_rdata));
  assign f646_clk = clk;
  assign f646_rst = rst;
  // Bindings to f646

  // f648
  logic [0:0] f648_wen;
  logic [31:0] f648_wdata;
  logic [0:0] f648_clk;
  logic [0:0] f648_rst;
  logic [31:0] f648_rdata;
  sr_buffer_32_1 f648(.wen(f648_wen), .wdata(f648_wdata), .clk(f648_clk), .rst(f648_rst), .rdata(f648_rdata));
  assign f648_clk = clk;
  assign f648_rst = rst;
  // Bindings to f648

  // f650
  logic [0:0] f650_wen;
  logic [31:0] f650_wdata;
  logic [0:0] f650_clk;
  logic [0:0] f650_rst;
  logic [31:0] f650_rdata;
  sr_buffer_32_1 f650(.wen(f650_wen), .wdata(f650_wdata), .clk(f650_clk), .rst(f650_rst), .rdata(f650_rdata));
  assign f650_clk = clk;
  assign f650_rst = rst;
  // Bindings to f650

  // f652
  logic [0:0] f652_wen;
  logic [31:0] f652_wdata;
  logic [0:0] f652_clk;
  logic [0:0] f652_rst;
  logic [31:0] f652_rdata;
  sr_buffer_32_1 f652(.wen(f652_wen), .wdata(f652_wdata), .clk(f652_clk), .rst(f652_rst), .rdata(f652_rdata));
  assign f652_clk = clk;
  assign f652_rst = rst;
  // Bindings to f652

  // f654
  logic [0:0] f654_wen;
  logic [31:0] f654_wdata;
  logic [0:0] f654_clk;
  logic [0:0] f654_rst;
  logic [31:0] f654_rdata;
  sr_buffer_32_1 f654(.wen(f654_wen), .wdata(f654_wdata), .clk(f654_clk), .rst(f654_rst), .rdata(f654_rdata));
  assign f654_clk = clk;
  assign f654_rst = rst;
  // Bindings to f654

  // f656
  logic [0:0] f656_wen;
  logic [31:0] f656_wdata;
  logic [0:0] f656_clk;
  logic [0:0] f656_rst;
  logic [31:0] f656_rdata;
  sr_buffer_32_1 f656(.wen(f656_wen), .wdata(f656_wdata), .clk(f656_clk), .rst(f656_rst), .rdata(f656_rdata));
  assign f656_clk = clk;
  assign f656_rst = rst;
  // Bindings to f656

  // f658
  logic [0:0] f658_wen;
  logic [31:0] f658_wdata;
  logic [0:0] f658_clk;
  logic [0:0] f658_rst;
  logic [31:0] f658_rdata;
  sr_buffer_32_1 f658(.wen(f658_wen), .wdata(f658_wdata), .clk(f658_clk), .rst(f658_rst), .rdata(f658_rdata));
  assign f658_clk = clk;
  assign f658_rst = rst;
  // Bindings to f658

  // f660
  logic [0:0] f660_wen;
  logic [31:0] f660_wdata;
  logic [0:0] f660_clk;
  logic [0:0] f660_rst;
  logic [31:0] f660_rdata;
  sr_buffer_32_1 f660(.wen(f660_wen), .wdata(f660_wdata), .clk(f660_clk), .rst(f660_rst), .rdata(f660_rdata));
  assign f660_clk = clk;
  assign f660_rst = rst;
  // Bindings to f660

  // f662
  logic [0:0] f662_wen;
  logic [31:0] f662_wdata;
  logic [0:0] f662_clk;
  logic [0:0] f662_rst;
  logic [31:0] f662_rdata;
  sr_buffer_32_1 f662(.wen(f662_wen), .wdata(f662_wdata), .clk(f662_clk), .rst(f662_rst), .rdata(f662_rdata));
  assign f662_clk = clk;
  assign f662_rst = rst;
  // Bindings to f662

  // f664
  logic [0:0] f664_wen;
  logic [31:0] f664_wdata;
  logic [0:0] f664_clk;
  logic [0:0] f664_rst;
  logic [31:0] f664_rdata;
  sr_buffer_32_1 f664(.wen(f664_wen), .wdata(f664_wdata), .clk(f664_clk), .rst(f664_rst), .rdata(f664_rdata));
  assign f664_clk = clk;
  assign f664_rst = rst;
  // Bindings to f664

  // f666
  logic [0:0] f666_wen;
  logic [31:0] f666_wdata;
  logic [0:0] f666_clk;
  logic [0:0] f666_rst;
  logic [31:0] f666_rdata;
  sr_buffer_32_1 f666(.wen(f666_wen), .wdata(f666_wdata), .clk(f666_clk), .rst(f666_rst), .rdata(f666_rdata));
  assign f666_clk = clk;
  assign f666_rst = rst;
  // Bindings to f666

  // f668
  logic [0:0] f668_wen;
  logic [31:0] f668_wdata;
  logic [0:0] f668_clk;
  logic [0:0] f668_rst;
  logic [31:0] f668_rdata;
  sr_buffer_32_1 f668(.wen(f668_wen), .wdata(f668_wdata), .clk(f668_clk), .rst(f668_rst), .rdata(f668_rdata));
  assign f668_clk = clk;
  assign f668_rst = rst;
  // Bindings to f668

  // f670
  logic [0:0] f670_wen;
  logic [31:0] f670_wdata;
  logic [0:0] f670_clk;
  logic [0:0] f670_rst;
  logic [31:0] f670_rdata;
  sr_buffer_32_1 f670(.wen(f670_wen), .wdata(f670_wdata), .clk(f670_clk), .rst(f670_rst), .rdata(f670_rdata));
  assign f670_clk = clk;
  assign f670_rst = rst;
  // Bindings to f670

  // f672
  logic [0:0] f672_wen;
  logic [31:0] f672_wdata;
  logic [0:0] f672_clk;
  logic [0:0] f672_rst;
  logic [31:0] f672_rdata;
  sr_buffer_32_1 f672(.wen(f672_wen), .wdata(f672_wdata), .clk(f672_clk), .rst(f672_rst), .rdata(f672_rdata));
  assign f672_clk = clk;
  assign f672_rst = rst;
  // Bindings to f672

  // f674
  logic [0:0] f674_wen;
  logic [31:0] f674_wdata;
  logic [0:0] f674_clk;
  logic [0:0] f674_rst;
  logic [31:0] f674_rdata;
  sr_buffer_32_1 f674(.wen(f674_wen), .wdata(f674_wdata), .clk(f674_clk), .rst(f674_rst), .rdata(f674_rdata));
  assign f674_clk = clk;
  assign f674_rst = rst;
  // Bindings to f674



endmodule


module bright_weights_normed_gauss_blur_1_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 113;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 224;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_1_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (107 - d0 >= 0) ? (222) : (-108 + d0 == 0) ? (222) : 0;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_1_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_1_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 223;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_1_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 112;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_1_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_1_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_weights_normed_update_0_write_wen(output [0:0] bright_weights_normed_update_0_write_wen);

endmodule


module bright_weights_normed_gauss_blur_1_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (107 - d0 >= 0) ? (111) : (-108 + d0 == 0) ? (111) : 0;
    end
  end

endmodule


module in_wire_bright_weights_normed_update_0_write_wdata(output [31:0] bright_weights_normed_update_0_write_wdata);

endmodule


module in_wire_bright_weights_normed_gauss_blur_1_update_0_read_dummy(output [287:0] bright_weights_normed_gauss_blur_1_update_0_read_dummy);

endmodule


module out_wire_bright_weights_normed_gauss_blur_1_update_0_read_rdata(input [287:0] bright_weights_normed_gauss_blur_1_update_0_read_rdata);

endmodule


module bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_279 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114



endmodule


module bright_weights_normed_gauss_blur_2_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 111;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_2_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 112;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_2_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 57;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_2_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (51 - d0 >= 0) ? (110) : (-52 + d0 == 0) ? (110) : 0;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_2_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 56;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_2_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_2_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_weights_normed_gauss_ds_1_update_0_write_wen(output [0:0] bright_weights_normed_gauss_ds_1_update_0_write_wen);

endmodule


module bright_weights_normed_gauss_blur_2_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (51 - d0 >= 0) ? (55) : (-52 + d0 == 0) ? (55) : 0;
    end
  end

endmodule


module in_wire_bright_weights_normed_gauss_ds_1_update_0_write_wdata(output [31:0] bright_weights_normed_gauss_ds_1_update_0_write_wdata);

endmodule


module in_wire_bright_weights_normed_gauss_blur_2_update_0_read_dummy(output [287:0] bright_weights_normed_gauss_blur_2_update_0_read_dummy);

endmodule


module out_wire_bright_weights_normed_gauss_blur_2_update_0_read_rdata(input [287:0] bright_weights_normed_gauss_blur_2_update_0_read_rdata);

endmodule


module dark_gauss_blur_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_gauss_blur_3_update_0_write_wen, input [31:0] dark_gauss_ds_3_update_0_read_dummy, input [31:0] dark_gauss_blur_3_update_0_write_wdata, output [31:0] dark_gauss_ds_3_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_gauss_blur_3_update_0_write_wen
    // rd_0
  assign rd_0 = dark_gauss_blur_3_update_0_write_wen;

  // dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1
  logic [0:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_done;
  dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1 dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1(.clk(dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_clk), .rst(dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_rst), .start(dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_start), .done(dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_done));
  assign dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_clk = clk;
  assign dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1

  // selector_dark_gauss_ds_3_rd0_select
  logic [0:0] selector_dark_gauss_ds_3_rd0_select_clk;
  logic [0:0] selector_dark_gauss_ds_3_rd0_select_rst;
  logic [31:0] selector_dark_gauss_ds_3_rd0_select_d0;
  logic [31:0] selector_dark_gauss_ds_3_rd0_select_d1;
  logic [31:0] selector_dark_gauss_ds_3_rd0_select_out;
  dark_gauss_ds_3_rd0_select selector_dark_gauss_ds_3_rd0_select(.clk(selector_dark_gauss_ds_3_rd0_select_clk), .rst(selector_dark_gauss_ds_3_rd0_select_rst), .d0(selector_dark_gauss_ds_3_rd0_select_d0), .d1(selector_dark_gauss_ds_3_rd0_select_d1), .out(selector_dark_gauss_ds_3_rd0_select_out));
  assign selector_dark_gauss_ds_3_rd0_select_clk = clk;
  assign selector_dark_gauss_ds_3_rd0_select_rst = rst;
  // Bindings to selector_dark_gauss_ds_3_rd0_select

  // Bindings to dark_gauss_ds_3_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_gauss_ds_3_update_0_read_dummy;

  // Bindings to dark_gauss_blur_3_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_gauss_blur_3_update_0_write_wdata;

  // Bindings to dark_gauss_ds_3_update_0_read_rdata
    // wr_3
  assign dark_gauss_ds_3_update_0_read_rdata = rd_2;



endmodule


module dark_weights_normed_gauss_blur_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_weights_normed_gauss_blur_3_update_0_write_wen, input [31:0] dark_weights_normed_gauss_blur_3_update_0_write_wdata, input [31:0] dark_weights_normed_gauss_ds_3_update_0_read_dummy, output [31:0] dark_weights_normed_gauss_ds_3_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1
  logic [0:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_done;
  dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1 dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1(.clk(dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_clk), .rst(dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_rst), .start(dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_start), .done(dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_done));
  assign dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_clk = clk;
  assign dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1

  // Bindings to dark_weights_normed_gauss_blur_3_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_normed_gauss_blur_3_update_0_write_wen;

  // selector_dark_weights_normed_gauss_ds_3_rd0_select
  logic [0:0] selector_dark_weights_normed_gauss_ds_3_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_ds_3_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_ds_3_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_ds_3_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_ds_3_rd0_select_out;
  dark_weights_normed_gauss_ds_3_rd0_select selector_dark_weights_normed_gauss_ds_3_rd0_select(.clk(selector_dark_weights_normed_gauss_ds_3_rd0_select_clk), .rst(selector_dark_weights_normed_gauss_ds_3_rd0_select_rst), .d0(selector_dark_weights_normed_gauss_ds_3_rd0_select_d0), .d1(selector_dark_weights_normed_gauss_ds_3_rd0_select_d1), .out(selector_dark_weights_normed_gauss_ds_3_rd0_select_out));
  assign selector_dark_weights_normed_gauss_ds_3_rd0_select_clk = clk;
  assign selector_dark_weights_normed_gauss_ds_3_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_ds_3_rd0_select

  // Bindings to dark_weights_normed_gauss_blur_3_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_normed_gauss_blur_3_update_0_write_wdata;

  // Bindings to dark_weights_normed_gauss_ds_3_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_weights_normed_gauss_ds_3_update_0_read_dummy;

  // Bindings to dark_weights_normed_gauss_ds_3_update_0_read_rdata
    // wr_3
  assign dark_weights_normed_gauss_ds_3_update_0_read_rdata = rd_2;



endmodule


module dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_108 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_108 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16



endmodule


module dark_weights_normed_gauss_blur_2_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 112;
    end
  end

endmodule


module dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_to_fused_level_1_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_279 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module dark_weights_normed_gauss_blur_2_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (51 - d0 >= 0) ? (110) : (-52 + d0 == 0) ? (110) : 0;
    end
  end

endmodule


module dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_9(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_52 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_52 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0



endmodule


module dark_weights_normed_gauss_blur_2_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 57;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_2_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 111;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_2_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 56;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_2_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_2_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module in_wire_dark_weights_normed_gauss_ds_1_update_0_write_wen(output [0:0] dark_weights_normed_gauss_ds_1_update_0_write_wen);

endmodule


module fused_level_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (-49 + d0 == 0 && 48 - d1 >= 0) ? (335) : (48 - d1 >= 0 && 48 - d0 >= 0) ? (336) : (-49 + d1 == 0) ? ((329 - d0)) : 0;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_2_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (51 - d0 >= 0) ? (55) : (-52 + d0 == 0) ? (55) : 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_gauss_ds_1_update_0_write_wdata(output [31:0] dark_weights_normed_gauss_ds_1_update_0_write_wdata);

endmodule


module in_wire_dark_weights_normed_gauss_blur_2_update_0_read_dummy(output [287:0] dark_weights_normed_gauss_blur_2_update_0_read_dummy);

endmodule


module out_wire_dark_weights_normed_gauss_blur_2_update_0_read_rdata(input [287:0] dark_weights_normed_gauss_blur_2_update_0_read_rdata);

endmodule


module dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_24 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_24 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16



endmodule


module dark_weights_normed_gauss_blur_3_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 28;
    end
  end

endmodule


module in_wire_dark_weights_normed_gauss_ds_2_update_0_write_wen(output [0:0] dark_weights_normed_gauss_ds_2_update_0_write_wen);

endmodule


module dark_weights_normed_gauss_blur_3_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 29;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 56;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_3_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_3_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 55;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_3_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_3_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (23 - d0 >= 0) ? (54) : (-24 + d0 == 0) ? (54) : 0;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_3_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module fused_level_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 56;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_3_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (23 - d0 >= 0) ? (27) : (-24 + d0 == 0) ? (27) : 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_gauss_ds_2_update_0_write_wdata(output [31:0] dark_weights_normed_gauss_ds_2_update_0_write_wdata);

endmodule


module in_wire_dark_weights_normed_gauss_blur_3_update_0_read_dummy(output [287:0] dark_weights_normed_gauss_blur_3_update_0_read_dummy);

endmodule


module out_wire_dark_weights_normed_gauss_blur_3_update_0_read_rdata(input [287:0] dark_weights_normed_gauss_blur_3_update_0_read_rdata);

endmodule


module final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48



endmodule


module in_wire_final_merged_2_update_0_write_wen(output [0:0] final_merged_2_update_0_write_wen);

endmodule


module in_wire_final_merged_2_update_0_write_wdata(output [31:0] final_merged_2_update_0_write_wdata);

endmodule


module in_wire_final_merged_1_update_0_read_dummy(output [31:0] final_merged_1_update_0_read_dummy);

endmodule


module out_wire_final_merged_1_update_0_read_rdata(input [31:0] final_merged_1_update_0_read_rdata);

endmodule


module dark_laplace_diff_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module in_wire_fused_level_0_update_0_write_wen(output [0:0] fused_level_0_update_0_write_wen);

endmodule


module final_merged_0_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_fused_level_0_update_0_write_wdata(output [31:0] fused_level_0_update_0_write_wdata);

endmodule


module bright_weights_normed_gauss_blur_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_weights_normed_gauss_ds_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module fused_level_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1231 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f314
  logic [0:0] f314_wen;
  logic [31:0] f314_wdata;
  logic [0:0] f314_clk;
  logic [0:0] f314_rst;
  logic [31:0] f314_rdata;
  sr_buffer_32_1 f314(.wen(f314_wen), .wdata(f314_wdata), .clk(f314_clk), .rst(f314_rst), .rdata(f314_rdata));
  assign f314_clk = clk;
  assign f314_rst = rst;
  // Bindings to f314

  // f316
  logic [0:0] f316_wen;
  logic [31:0] f316_wdata;
  logic [0:0] f316_clk;
  logic [0:0] f316_rst;
  logic [31:0] f316_rdata;
  sr_buffer_32_1 f316(.wen(f316_wen), .wdata(f316_wdata), .clk(f316_clk), .rst(f316_rst), .rdata(f316_rdata));
  assign f316_clk = clk;
  assign f316_rst = rst;
  // Bindings to f316

  // f318
  logic [0:0] f318_wen;
  logic [31:0] f318_wdata;
  logic [0:0] f318_clk;
  logic [0:0] f318_rst;
  logic [31:0] f318_rdata;
  sr_buffer_32_1 f318(.wen(f318_wen), .wdata(f318_wdata), .clk(f318_clk), .rst(f318_rst), .rdata(f318_rdata));
  assign f318_clk = clk;
  assign f318_rst = rst;
  // Bindings to f318

  // f320
  logic [0:0] f320_wen;
  logic [31:0] f320_wdata;
  logic [0:0] f320_clk;
  logic [0:0] f320_rst;
  logic [31:0] f320_rdata;
  sr_buffer_32_1 f320(.wen(f320_wen), .wdata(f320_wdata), .clk(f320_clk), .rst(f320_rst), .rdata(f320_rdata));
  assign f320_clk = clk;
  assign f320_rst = rst;
  // Bindings to f320

  // f322
  logic [0:0] f322_wen;
  logic [31:0] f322_wdata;
  logic [0:0] f322_clk;
  logic [0:0] f322_rst;
  logic [31:0] f322_rdata;
  sr_buffer_32_1 f322(.wen(f322_wen), .wdata(f322_wdata), .clk(f322_clk), .rst(f322_rst), .rdata(f322_rdata));
  assign f322_clk = clk;
  assign f322_rst = rst;
  // Bindings to f322

  // f324
  logic [0:0] f324_wen;
  logic [31:0] f324_wdata;
  logic [0:0] f324_clk;
  logic [0:0] f324_rst;
  logic [31:0] f324_rdata;
  sr_buffer_32_1 f324(.wen(f324_wen), .wdata(f324_wdata), .clk(f324_clk), .rst(f324_rst), .rdata(f324_rdata));
  assign f324_clk = clk;
  assign f324_rst = rst;
  // Bindings to f324

  // f326
  logic [0:0] f326_wen;
  logic [31:0] f326_wdata;
  logic [0:0] f326_clk;
  logic [0:0] f326_rst;
  logic [31:0] f326_rdata;
  sr_buffer_32_1 f326(.wen(f326_wen), .wdata(f326_wdata), .clk(f326_clk), .rst(f326_rst), .rdata(f326_rdata));
  assign f326_clk = clk;
  assign f326_rst = rst;
  // Bindings to f326

  // f328
  logic [0:0] f328_wen;
  logic [31:0] f328_wdata;
  logic [0:0] f328_clk;
  logic [0:0] f328_rst;
  logic [31:0] f328_rdata;
  sr_buffer_32_1 f328(.wen(f328_wen), .wdata(f328_wdata), .clk(f328_clk), .rst(f328_rst), .rdata(f328_rdata));
  assign f328_clk = clk;
  assign f328_rst = rst;
  // Bindings to f328

  // f330
  logic [0:0] f330_wen;
  logic [31:0] f330_wdata;
  logic [0:0] f330_clk;
  logic [0:0] f330_rst;
  logic [31:0] f330_rdata;
  sr_buffer_32_1 f330(.wen(f330_wen), .wdata(f330_wdata), .clk(f330_clk), .rst(f330_rst), .rdata(f330_rdata));
  assign f330_clk = clk;
  assign f330_rst = rst;
  // Bindings to f330

  // f332
  logic [0:0] f332_wen;
  logic [31:0] f332_wdata;
  logic [0:0] f332_clk;
  logic [0:0] f332_rst;
  logic [31:0] f332_rdata;
  sr_buffer_32_1 f332(.wen(f332_wen), .wdata(f332_wdata), .clk(f332_clk), .rst(f332_rst), .rdata(f332_rdata));
  assign f332_clk = clk;
  assign f332_rst = rst;
  // Bindings to f332

  // f334
  logic [0:0] f334_wen;
  logic [31:0] f334_wdata;
  logic [0:0] f334_clk;
  logic [0:0] f334_rst;
  logic [31:0] f334_rdata;
  sr_buffer_32_1 f334(.wen(f334_wen), .wdata(f334_wdata), .clk(f334_clk), .rst(f334_rst), .rdata(f334_rdata));
  assign f334_clk = clk;
  assign f334_rst = rst;
  // Bindings to f334

  // f336
  logic [0:0] f336_wen;
  logic [31:0] f336_wdata;
  logic [0:0] f336_clk;
  logic [0:0] f336_rst;
  logic [31:0] f336_rdata;
  sr_buffer_32_1 f336(.wen(f336_wen), .wdata(f336_wdata), .clk(f336_clk), .rst(f336_rst), .rdata(f336_rdata));
  assign f336_clk = clk;
  assign f336_rst = rst;
  // Bindings to f336

  // f338
  logic [0:0] f338_wen;
  logic [31:0] f338_wdata;
  logic [0:0] f338_clk;
  logic [0:0] f338_rst;
  logic [31:0] f338_rdata;
  sr_buffer_32_1 f338(.wen(f338_wen), .wdata(f338_wdata), .clk(f338_clk), .rst(f338_rst), .rdata(f338_rdata));
  assign f338_clk = clk;
  assign f338_rst = rst;
  // Bindings to f338

  // f340
  logic [0:0] f340_wen;
  logic [31:0] f340_wdata;
  logic [0:0] f340_clk;
  logic [0:0] f340_rst;
  logic [31:0] f340_rdata;
  sr_buffer_32_1 f340(.wen(f340_wen), .wdata(f340_wdata), .clk(f340_clk), .rst(f340_rst), .rdata(f340_rdata));
  assign f340_clk = clk;
  assign f340_rst = rst;
  // Bindings to f340

  // f342
  logic [0:0] f342_wen;
  logic [31:0] f342_wdata;
  logic [0:0] f342_clk;
  logic [0:0] f342_rst;
  logic [31:0] f342_rdata;
  sr_buffer_32_1 f342(.wen(f342_wen), .wdata(f342_wdata), .clk(f342_clk), .rst(f342_rst), .rdata(f342_rdata));
  assign f342_clk = clk;
  assign f342_rst = rst;
  // Bindings to f342

  // f344
  logic [0:0] f344_wen;
  logic [31:0] f344_wdata;
  logic [0:0] f344_clk;
  logic [0:0] f344_rst;
  logic [31:0] f344_rdata;
  sr_buffer_32_1 f344(.wen(f344_wen), .wdata(f344_wdata), .clk(f344_clk), .rst(f344_rst), .rdata(f344_rdata));
  assign f344_clk = clk;
  assign f344_rst = rst;
  // Bindings to f344

  // f346
  logic [0:0] f346_wen;
  logic [31:0] f346_wdata;
  logic [0:0] f346_clk;
  logic [0:0] f346_rst;
  logic [31:0] f346_rdata;
  sr_buffer_32_1 f346(.wen(f346_wen), .wdata(f346_wdata), .clk(f346_clk), .rst(f346_rst), .rdata(f346_rdata));
  assign f346_clk = clk;
  assign f346_rst = rst;
  // Bindings to f346

  // f348
  logic [0:0] f348_wen;
  logic [31:0] f348_wdata;
  logic [0:0] f348_clk;
  logic [0:0] f348_rst;
  logic [31:0] f348_rdata;
  sr_buffer_32_1 f348(.wen(f348_wen), .wdata(f348_wdata), .clk(f348_clk), .rst(f348_rst), .rdata(f348_rdata));
  assign f348_clk = clk;
  assign f348_rst = rst;
  // Bindings to f348

  // f350
  logic [0:0] f350_wen;
  logic [31:0] f350_wdata;
  logic [0:0] f350_clk;
  logic [0:0] f350_rst;
  logic [31:0] f350_rdata;
  sr_buffer_32_1 f350(.wen(f350_wen), .wdata(f350_wdata), .clk(f350_clk), .rst(f350_rst), .rdata(f350_rdata));
  assign f350_clk = clk;
  assign f350_rst = rst;
  // Bindings to f350

  // f352
  logic [0:0] f352_wen;
  logic [31:0] f352_wdata;
  logic [0:0] f352_clk;
  logic [0:0] f352_rst;
  logic [31:0] f352_rdata;
  sr_buffer_32_1 f352(.wen(f352_wen), .wdata(f352_wdata), .clk(f352_clk), .rst(f352_rst), .rdata(f352_rdata));
  assign f352_clk = clk;
  assign f352_rst = rst;
  // Bindings to f352

  // f354
  logic [0:0] f354_wen;
  logic [31:0] f354_wdata;
  logic [0:0] f354_clk;
  logic [0:0] f354_rst;
  logic [31:0] f354_rdata;
  sr_buffer_32_1 f354(.wen(f354_wen), .wdata(f354_wdata), .clk(f354_clk), .rst(f354_rst), .rdata(f354_rdata));
  assign f354_clk = clk;
  assign f354_rst = rst;
  // Bindings to f354

  // f356
  logic [0:0] f356_wen;
  logic [31:0] f356_wdata;
  logic [0:0] f356_clk;
  logic [0:0] f356_rst;
  logic [31:0] f356_rdata;
  sr_buffer_32_1 f356(.wen(f356_wen), .wdata(f356_wdata), .clk(f356_clk), .rst(f356_rst), .rdata(f356_rdata));
  assign f356_clk = clk;
  assign f356_rst = rst;
  // Bindings to f356

  // f358
  logic [0:0] f358_wen;
  logic [31:0] f358_wdata;
  logic [0:0] f358_clk;
  logic [0:0] f358_rst;
  logic [31:0] f358_rdata;
  sr_buffer_32_1 f358(.wen(f358_wen), .wdata(f358_wdata), .clk(f358_clk), .rst(f358_rst), .rdata(f358_rdata));
  assign f358_clk = clk;
  assign f358_rst = rst;
  // Bindings to f358

  // f360
  logic [0:0] f360_wen;
  logic [31:0] f360_wdata;
  logic [0:0] f360_clk;
  logic [0:0] f360_rst;
  logic [31:0] f360_rdata;
  sr_buffer_32_1 f360(.wen(f360_wen), .wdata(f360_wdata), .clk(f360_clk), .rst(f360_rst), .rdata(f360_rdata));
  assign f360_clk = clk;
  assign f360_rst = rst;
  // Bindings to f360

  // f362
  logic [0:0] f362_wen;
  logic [31:0] f362_wdata;
  logic [0:0] f362_clk;
  logic [0:0] f362_rst;
  logic [31:0] f362_rdata;
  sr_buffer_32_1 f362(.wen(f362_wen), .wdata(f362_wdata), .clk(f362_clk), .rst(f362_rst), .rdata(f362_rdata));
  assign f362_clk = clk;
  assign f362_rst = rst;
  // Bindings to f362

  // f364
  logic [0:0] f364_wen;
  logic [31:0] f364_wdata;
  logic [0:0] f364_clk;
  logic [0:0] f364_rst;
  logic [31:0] f364_rdata;
  sr_buffer_32_1 f364(.wen(f364_wen), .wdata(f364_wdata), .clk(f364_clk), .rst(f364_rst), .rdata(f364_rdata));
  assign f364_clk = clk;
  assign f364_rst = rst;
  // Bindings to f364

  // f366
  logic [0:0] f366_wen;
  logic [31:0] f366_wdata;
  logic [0:0] f366_clk;
  logic [0:0] f366_rst;
  logic [31:0] f366_rdata;
  sr_buffer_32_1 f366(.wen(f366_wen), .wdata(f366_wdata), .clk(f366_clk), .rst(f366_rst), .rdata(f366_rdata));
  assign f366_clk = clk;
  assign f366_rst = rst;
  // Bindings to f366

  // f368
  logic [0:0] f368_wen;
  logic [31:0] f368_wdata;
  logic [0:0] f368_clk;
  logic [0:0] f368_rst;
  logic [31:0] f368_rdata;
  sr_buffer_32_1 f368(.wen(f368_wen), .wdata(f368_wdata), .clk(f368_clk), .rst(f368_rst), .rdata(f368_rdata));
  assign f368_clk = clk;
  assign f368_rst = rst;
  // Bindings to f368

  // f370
  logic [0:0] f370_wen;
  logic [31:0] f370_wdata;
  logic [0:0] f370_clk;
  logic [0:0] f370_rst;
  logic [31:0] f370_rdata;
  sr_buffer_32_1 f370(.wen(f370_wen), .wdata(f370_wdata), .clk(f370_clk), .rst(f370_rst), .rdata(f370_rdata));
  assign f370_clk = clk;
  assign f370_rst = rst;
  // Bindings to f370

  // f372
  logic [0:0] f372_wen;
  logic [31:0] f372_wdata;
  logic [0:0] f372_clk;
  logic [0:0] f372_rst;
  logic [31:0] f372_rdata;
  sr_buffer_32_1 f372(.wen(f372_wen), .wdata(f372_wdata), .clk(f372_clk), .rst(f372_rst), .rdata(f372_rdata));
  assign f372_clk = clk;
  assign f372_rst = rst;
  // Bindings to f372

  // f374
  logic [0:0] f374_wen;
  logic [31:0] f374_wdata;
  logic [0:0] f374_clk;
  logic [0:0] f374_rst;
  logic [31:0] f374_rdata;
  sr_buffer_32_1 f374(.wen(f374_wen), .wdata(f374_wdata), .clk(f374_clk), .rst(f374_rst), .rdata(f374_rdata));
  assign f374_clk = clk;
  assign f374_rst = rst;
  // Bindings to f374

  // f376
  logic [0:0] f376_wen;
  logic [31:0] f376_wdata;
  logic [0:0] f376_clk;
  logic [0:0] f376_rst;
  logic [31:0] f376_rdata;
  sr_buffer_32_1 f376(.wen(f376_wen), .wdata(f376_wdata), .clk(f376_clk), .rst(f376_rst), .rdata(f376_rdata));
  assign f376_clk = clk;
  assign f376_rst = rst;
  // Bindings to f376

  // f378
  logic [0:0] f378_wen;
  logic [31:0] f378_wdata;
  logic [0:0] f378_clk;
  logic [0:0] f378_rst;
  logic [31:0] f378_rdata;
  sr_buffer_32_1 f378(.wen(f378_wen), .wdata(f378_wdata), .clk(f378_clk), .rst(f378_rst), .rdata(f378_rdata));
  assign f378_clk = clk;
  assign f378_rst = rst;
  // Bindings to f378

  // f380
  logic [0:0] f380_wen;
  logic [31:0] f380_wdata;
  logic [0:0] f380_clk;
  logic [0:0] f380_rst;
  logic [31:0] f380_rdata;
  sr_buffer_32_1 f380(.wen(f380_wen), .wdata(f380_wdata), .clk(f380_clk), .rst(f380_rst), .rdata(f380_rdata));
  assign f380_clk = clk;
  assign f380_rst = rst;
  // Bindings to f380

  // f382
  logic [0:0] f382_wen;
  logic [31:0] f382_wdata;
  logic [0:0] f382_clk;
  logic [0:0] f382_rst;
  logic [31:0] f382_rdata;
  sr_buffer_32_1 f382(.wen(f382_wen), .wdata(f382_wdata), .clk(f382_clk), .rst(f382_rst), .rdata(f382_rdata));
  assign f382_clk = clk;
  assign f382_rst = rst;
  // Bindings to f382

  // f384
  logic [0:0] f384_wen;
  logic [31:0] f384_wdata;
  logic [0:0] f384_clk;
  logic [0:0] f384_rst;
  logic [31:0] f384_rdata;
  sr_buffer_32_1 f384(.wen(f384_wen), .wdata(f384_wdata), .clk(f384_clk), .rst(f384_rst), .rdata(f384_rdata));
  assign f384_clk = clk;
  assign f384_rst = rst;
  // Bindings to f384

  // f386
  logic [0:0] f386_wen;
  logic [31:0] f386_wdata;
  logic [0:0] f386_clk;
  logic [0:0] f386_rst;
  logic [31:0] f386_rdata;
  sr_buffer_32_1 f386(.wen(f386_wen), .wdata(f386_wdata), .clk(f386_clk), .rst(f386_rst), .rdata(f386_rdata));
  assign f386_clk = clk;
  assign f386_rst = rst;
  // Bindings to f386

  // f388
  logic [0:0] f388_wen;
  logic [31:0] f388_wdata;
  logic [0:0] f388_clk;
  logic [0:0] f388_rst;
  logic [31:0] f388_rdata;
  sr_buffer_32_1 f388(.wen(f388_wen), .wdata(f388_wdata), .clk(f388_clk), .rst(f388_rst), .rdata(f388_rdata));
  assign f388_clk = clk;
  assign f388_rst = rst;
  // Bindings to f388

  // f390
  logic [0:0] f390_wen;
  logic [31:0] f390_wdata;
  logic [0:0] f390_clk;
  logic [0:0] f390_rst;
  logic [31:0] f390_rdata;
  sr_buffer_32_1 f390(.wen(f390_wen), .wdata(f390_wdata), .clk(f390_clk), .rst(f390_rst), .rdata(f390_rdata));
  assign f390_clk = clk;
  assign f390_rst = rst;
  // Bindings to f390

  // f392
  logic [0:0] f392_wen;
  logic [31:0] f392_wdata;
  logic [0:0] f392_clk;
  logic [0:0] f392_rst;
  logic [31:0] f392_rdata;
  sr_buffer_32_1 f392(.wen(f392_wen), .wdata(f392_wdata), .clk(f392_clk), .rst(f392_rst), .rdata(f392_rdata));
  assign f392_clk = clk;
  assign f392_rst = rst;
  // Bindings to f392

  // f394
  logic [0:0] f394_wen;
  logic [31:0] f394_wdata;
  logic [0:0] f394_clk;
  logic [0:0] f394_rst;
  logic [31:0] f394_rdata;
  sr_buffer_32_1 f394(.wen(f394_wen), .wdata(f394_wdata), .clk(f394_clk), .rst(f394_rst), .rdata(f394_rdata));
  assign f394_clk = clk;
  assign f394_rst = rst;
  // Bindings to f394

  // f396
  logic [0:0] f396_wen;
  logic [31:0] f396_wdata;
  logic [0:0] f396_clk;
  logic [0:0] f396_rst;
  logic [31:0] f396_rdata;
  sr_buffer_32_1 f396(.wen(f396_wen), .wdata(f396_wdata), .clk(f396_clk), .rst(f396_rst), .rdata(f396_rdata));
  assign f396_clk = clk;
  assign f396_rst = rst;
  // Bindings to f396

  // f398
  logic [0:0] f398_wen;
  logic [31:0] f398_wdata;
  logic [0:0] f398_clk;
  logic [0:0] f398_rst;
  logic [31:0] f398_rdata;
  sr_buffer_32_1 f398(.wen(f398_wen), .wdata(f398_wdata), .clk(f398_clk), .rst(f398_rst), .rdata(f398_rdata));
  assign f398_clk = clk;
  assign f398_rst = rst;
  // Bindings to f398

  // f400
  logic [0:0] f400_wen;
  logic [31:0] f400_wdata;
  logic [0:0] f400_clk;
  logic [0:0] f400_rst;
  logic [31:0] f400_rdata;
  sr_buffer_32_1 f400(.wen(f400_wen), .wdata(f400_wdata), .clk(f400_clk), .rst(f400_rst), .rdata(f400_rdata));
  assign f400_clk = clk;
  assign f400_rst = rst;
  // Bindings to f400

  // f402
  logic [0:0] f402_wen;
  logic [31:0] f402_wdata;
  logic [0:0] f402_clk;
  logic [0:0] f402_rst;
  logic [31:0] f402_rdata;
  sr_buffer_32_1 f402(.wen(f402_wen), .wdata(f402_wdata), .clk(f402_clk), .rst(f402_rst), .rdata(f402_rdata));
  assign f402_clk = clk;
  assign f402_rst = rst;
  // Bindings to f402

  // f404
  logic [0:0] f404_wen;
  logic [31:0] f404_wdata;
  logic [0:0] f404_clk;
  logic [0:0] f404_rst;
  logic [31:0] f404_rdata;
  sr_buffer_32_1 f404(.wen(f404_wen), .wdata(f404_wdata), .clk(f404_clk), .rst(f404_rst), .rdata(f404_rdata));
  assign f404_clk = clk;
  assign f404_rst = rst;
  // Bindings to f404

  // f406
  logic [0:0] f406_wen;
  logic [31:0] f406_wdata;
  logic [0:0] f406_clk;
  logic [0:0] f406_rst;
  logic [31:0] f406_rdata;
  sr_buffer_32_1 f406(.wen(f406_wen), .wdata(f406_wdata), .clk(f406_clk), .rst(f406_rst), .rdata(f406_rdata));
  assign f406_clk = clk;
  assign f406_rst = rst;
  // Bindings to f406

  // f408
  logic [0:0] f408_wen;
  logic [31:0] f408_wdata;
  logic [0:0] f408_clk;
  logic [0:0] f408_rst;
  logic [31:0] f408_rdata;
  sr_buffer_32_1 f408(.wen(f408_wen), .wdata(f408_wdata), .clk(f408_clk), .rst(f408_rst), .rdata(f408_rdata));
  assign f408_clk = clk;
  assign f408_rst = rst;
  // Bindings to f408

  // f410
  logic [0:0] f410_wen;
  logic [31:0] f410_wdata;
  logic [0:0] f410_clk;
  logic [0:0] f410_rst;
  logic [31:0] f410_rdata;
  sr_buffer_32_1 f410(.wen(f410_wen), .wdata(f410_wdata), .clk(f410_clk), .rst(f410_rst), .rdata(f410_rdata));
  assign f410_clk = clk;
  assign f410_rst = rst;
  // Bindings to f410

  // f412
  logic [0:0] f412_wen;
  logic [31:0] f412_wdata;
  logic [0:0] f412_clk;
  logic [0:0] f412_rst;
  logic [31:0] f412_rdata;
  sr_buffer_32_1 f412(.wen(f412_wen), .wdata(f412_wdata), .clk(f412_clk), .rst(f412_rst), .rdata(f412_rdata));
  assign f412_clk = clk;
  assign f412_rst = rst;
  // Bindings to f412

  // f414
  logic [0:0] f414_wen;
  logic [31:0] f414_wdata;
  logic [0:0] f414_clk;
  logic [0:0] f414_rst;
  logic [31:0] f414_rdata;
  sr_buffer_32_1 f414(.wen(f414_wen), .wdata(f414_wdata), .clk(f414_clk), .rst(f414_rst), .rdata(f414_rdata));
  assign f414_clk = clk;
  assign f414_rst = rst;
  // Bindings to f414

  // f416
  logic [0:0] f416_wen;
  logic [31:0] f416_wdata;
  logic [0:0] f416_clk;
  logic [0:0] f416_rst;
  logic [31:0] f416_rdata;
  sr_buffer_32_1 f416(.wen(f416_wen), .wdata(f416_wdata), .clk(f416_clk), .rst(f416_rst), .rdata(f416_rdata));
  assign f416_clk = clk;
  assign f416_rst = rst;
  // Bindings to f416

  // f418
  logic [0:0] f418_wen;
  logic [31:0] f418_wdata;
  logic [0:0] f418_clk;
  logic [0:0] f418_rst;
  logic [31:0] f418_rdata;
  sr_buffer_32_1 f418(.wen(f418_wen), .wdata(f418_wdata), .clk(f418_clk), .rst(f418_rst), .rdata(f418_rdata));
  assign f418_clk = clk;
  assign f418_rst = rst;
  // Bindings to f418

  // f420
  logic [0:0] f420_wen;
  logic [31:0] f420_wdata;
  logic [0:0] f420_clk;
  logic [0:0] f420_rst;
  logic [31:0] f420_rdata;
  sr_buffer_32_1 f420(.wen(f420_wen), .wdata(f420_wdata), .clk(f420_clk), .rst(f420_rst), .rdata(f420_rdata));
  assign f420_clk = clk;
  assign f420_rst = rst;
  // Bindings to f420

  // f422
  logic [0:0] f422_wen;
  logic [31:0] f422_wdata;
  logic [0:0] f422_clk;
  logic [0:0] f422_rst;
  logic [31:0] f422_rdata;
  sr_buffer_32_1 f422(.wen(f422_wen), .wdata(f422_wdata), .clk(f422_clk), .rst(f422_rst), .rdata(f422_rdata));
  assign f422_clk = clk;
  assign f422_rst = rst;
  // Bindings to f422

  // f424
  logic [0:0] f424_wen;
  logic [31:0] f424_wdata;
  logic [0:0] f424_clk;
  logic [0:0] f424_rst;
  logic [31:0] f424_rdata;
  sr_buffer_32_1 f424(.wen(f424_wen), .wdata(f424_wdata), .clk(f424_clk), .rst(f424_rst), .rdata(f424_rdata));
  assign f424_clk = clk;
  assign f424_rst = rst;
  // Bindings to f424

  // f426
  logic [0:0] f426_wen;
  logic [31:0] f426_wdata;
  logic [0:0] f426_clk;
  logic [0:0] f426_rst;
  logic [31:0] f426_rdata;
  sr_buffer_32_1 f426(.wen(f426_wen), .wdata(f426_wdata), .clk(f426_clk), .rst(f426_rst), .rdata(f426_rdata));
  assign f426_clk = clk;
  assign f426_rst = rst;
  // Bindings to f426

  // f428
  logic [0:0] f428_wen;
  logic [31:0] f428_wdata;
  logic [0:0] f428_clk;
  logic [0:0] f428_rst;
  logic [31:0] f428_rdata;
  sr_buffer_32_1 f428(.wen(f428_wen), .wdata(f428_wdata), .clk(f428_clk), .rst(f428_rst), .rdata(f428_rdata));
  assign f428_clk = clk;
  assign f428_rst = rst;
  // Bindings to f428

  // f430
  logic [0:0] f430_wen;
  logic [31:0] f430_wdata;
  logic [0:0] f430_clk;
  logic [0:0] f430_rst;
  logic [31:0] f430_rdata;
  sr_buffer_32_1 f430(.wen(f430_wen), .wdata(f430_wdata), .clk(f430_clk), .rst(f430_rst), .rdata(f430_rdata));
  assign f430_clk = clk;
  assign f430_rst = rst;
  // Bindings to f430

  // f432
  logic [0:0] f432_wen;
  logic [31:0] f432_wdata;
  logic [0:0] f432_clk;
  logic [0:0] f432_rst;
  logic [31:0] f432_rdata;
  sr_buffer_32_1 f432(.wen(f432_wen), .wdata(f432_wdata), .clk(f432_clk), .rst(f432_rst), .rdata(f432_rdata));
  assign f432_clk = clk;
  assign f432_rst = rst;
  // Bindings to f432

  // f434
  logic [0:0] f434_wen;
  logic [31:0] f434_wdata;
  logic [0:0] f434_clk;
  logic [0:0] f434_rst;
  logic [31:0] f434_rdata;
  sr_buffer_32_1 f434(.wen(f434_wen), .wdata(f434_wdata), .clk(f434_clk), .rst(f434_rst), .rdata(f434_rdata));
  assign f434_clk = clk;
  assign f434_rst = rst;
  // Bindings to f434

  // f436
  logic [0:0] f436_wen;
  logic [31:0] f436_wdata;
  logic [0:0] f436_clk;
  logic [0:0] f436_rst;
  logic [31:0] f436_rdata;
  sr_buffer_32_1 f436(.wen(f436_wen), .wdata(f436_wdata), .clk(f436_clk), .rst(f436_rst), .rdata(f436_rdata));
  assign f436_clk = clk;
  assign f436_rst = rst;
  // Bindings to f436

  // f438
  logic [0:0] f438_wen;
  logic [31:0] f438_wdata;
  logic [0:0] f438_clk;
  logic [0:0] f438_rst;
  logic [31:0] f438_rdata;
  sr_buffer_32_1 f438(.wen(f438_wen), .wdata(f438_wdata), .clk(f438_clk), .rst(f438_rst), .rdata(f438_rdata));
  assign f438_clk = clk;
  assign f438_rst = rst;
  // Bindings to f438

  // f440
  logic [0:0] f440_wen;
  logic [31:0] f440_wdata;
  logic [0:0] f440_clk;
  logic [0:0] f440_rst;
  logic [31:0] f440_rdata;
  sr_buffer_32_1 f440(.wen(f440_wen), .wdata(f440_wdata), .clk(f440_clk), .rst(f440_rst), .rdata(f440_rdata));
  assign f440_clk = clk;
  assign f440_rst = rst;
  // Bindings to f440

  // f442
  logic [0:0] f442_wen;
  logic [31:0] f442_wdata;
  logic [0:0] f442_clk;
  logic [0:0] f442_rst;
  logic [31:0] f442_rdata;
  sr_buffer_32_1 f442(.wen(f442_wen), .wdata(f442_wdata), .clk(f442_clk), .rst(f442_rst), .rdata(f442_rdata));
  assign f442_clk = clk;
  assign f442_rst = rst;
  // Bindings to f442

  // f444
  logic [0:0] f444_wen;
  logic [31:0] f444_wdata;
  logic [0:0] f444_clk;
  logic [0:0] f444_rst;
  logic [31:0] f444_rdata;
  sr_buffer_32_1 f444(.wen(f444_wen), .wdata(f444_wdata), .clk(f444_clk), .rst(f444_rst), .rdata(f444_rdata));
  assign f444_clk = clk;
  assign f444_rst = rst;
  // Bindings to f444

  // f446
  logic [0:0] f446_wen;
  logic [31:0] f446_wdata;
  logic [0:0] f446_clk;
  logic [0:0] f446_rst;
  logic [31:0] f446_rdata;
  sr_buffer_32_1 f446(.wen(f446_wen), .wdata(f446_wdata), .clk(f446_clk), .rst(f446_rst), .rdata(f446_rdata));
  assign f446_clk = clk;
  assign f446_rst = rst;
  // Bindings to f446

  // f448
  logic [0:0] f448_wen;
  logic [31:0] f448_wdata;
  logic [0:0] f448_clk;
  logic [0:0] f448_rst;
  logic [31:0] f448_rdata;
  sr_buffer_32_1 f448(.wen(f448_wen), .wdata(f448_wdata), .clk(f448_clk), .rst(f448_rst), .rdata(f448_rdata));
  assign f448_clk = clk;
  assign f448_rst = rst;
  // Bindings to f448

  // f450
  logic [0:0] f450_wen;
  logic [31:0] f450_wdata;
  logic [0:0] f450_clk;
  logic [0:0] f450_rst;
  logic [31:0] f450_rdata;
  sr_buffer_32_1 f450(.wen(f450_wen), .wdata(f450_wdata), .clk(f450_clk), .rst(f450_rst), .rdata(f450_rdata));
  assign f450_clk = clk;
  assign f450_rst = rst;
  // Bindings to f450

  // f452
  logic [0:0] f452_wen;
  logic [31:0] f452_wdata;
  logic [0:0] f452_clk;
  logic [0:0] f452_rst;
  logic [31:0] f452_rdata;
  sr_buffer_32_1 f452(.wen(f452_wen), .wdata(f452_wdata), .clk(f452_clk), .rst(f452_rst), .rdata(f452_rdata));
  assign f452_clk = clk;
  assign f452_rst = rst;
  // Bindings to f452

  // f454
  logic [0:0] f454_wen;
  logic [31:0] f454_wdata;
  logic [0:0] f454_clk;
  logic [0:0] f454_rst;
  logic [31:0] f454_rdata;
  sr_buffer_32_1 f454(.wen(f454_wen), .wdata(f454_wdata), .clk(f454_clk), .rst(f454_rst), .rdata(f454_rdata));
  assign f454_clk = clk;
  assign f454_rst = rst;
  // Bindings to f454

  // f456
  logic [0:0] f456_wen;
  logic [31:0] f456_wdata;
  logic [0:0] f456_clk;
  logic [0:0] f456_rst;
  logic [31:0] f456_rdata;
  sr_buffer_32_1 f456(.wen(f456_wen), .wdata(f456_wdata), .clk(f456_clk), .rst(f456_rst), .rdata(f456_rdata));
  assign f456_clk = clk;
  assign f456_rst = rst;
  // Bindings to f456

  // f458
  logic [0:0] f458_wen;
  logic [31:0] f458_wdata;
  logic [0:0] f458_clk;
  logic [0:0] f458_rst;
  logic [31:0] f458_rdata;
  sr_buffer_32_1 f458(.wen(f458_wen), .wdata(f458_wdata), .clk(f458_clk), .rst(f458_rst), .rdata(f458_rdata));
  assign f458_clk = clk;
  assign f458_rst = rst;
  // Bindings to f458

  // f460
  logic [0:0] f460_wen;
  logic [31:0] f460_wdata;
  logic [0:0] f460_clk;
  logic [0:0] f460_rst;
  logic [31:0] f460_rdata;
  sr_buffer_32_1 f460(.wen(f460_wen), .wdata(f460_wdata), .clk(f460_clk), .rst(f460_rst), .rdata(f460_rdata));
  assign f460_clk = clk;
  assign f460_rst = rst;
  // Bindings to f460

  // f462
  logic [0:0] f462_wen;
  logic [31:0] f462_wdata;
  logic [0:0] f462_clk;
  logic [0:0] f462_rst;
  logic [31:0] f462_rdata;
  sr_buffer_32_1 f462(.wen(f462_wen), .wdata(f462_wdata), .clk(f462_clk), .rst(f462_rst), .rdata(f462_rdata));
  assign f462_clk = clk;
  assign f462_rst = rst;
  // Bindings to f462

  // f464
  logic [0:0] f464_wen;
  logic [31:0] f464_wdata;
  logic [0:0] f464_clk;
  logic [0:0] f464_rst;
  logic [31:0] f464_rdata;
  sr_buffer_32_1 f464(.wen(f464_wen), .wdata(f464_wdata), .clk(f464_clk), .rst(f464_rst), .rdata(f464_rdata));
  assign f464_clk = clk;
  assign f464_rst = rst;
  // Bindings to f464

  // f466
  logic [0:0] f466_wen;
  logic [31:0] f466_wdata;
  logic [0:0] f466_clk;
  logic [0:0] f466_rst;
  logic [31:0] f466_rdata;
  sr_buffer_32_1 f466(.wen(f466_wen), .wdata(f466_wdata), .clk(f466_clk), .rst(f466_rst), .rdata(f466_rdata));
  assign f466_clk = clk;
  assign f466_rst = rst;
  // Bindings to f466

  // f468
  logic [0:0] f468_wen;
  logic [31:0] f468_wdata;
  logic [0:0] f468_clk;
  logic [0:0] f468_rst;
  logic [31:0] f468_rdata;
  sr_buffer_32_1 f468(.wen(f468_wen), .wdata(f468_wdata), .clk(f468_clk), .rst(f468_rst), .rdata(f468_rdata));
  assign f468_clk = clk;
  assign f468_rst = rst;
  // Bindings to f468

  // f470
  logic [0:0] f470_wen;
  logic [31:0] f470_wdata;
  logic [0:0] f470_clk;
  logic [0:0] f470_rst;
  logic [31:0] f470_rdata;
  sr_buffer_32_1 f470(.wen(f470_wen), .wdata(f470_wdata), .clk(f470_clk), .rst(f470_rst), .rdata(f470_rdata));
  assign f470_clk = clk;
  assign f470_rst = rst;
  // Bindings to f470

  // f472
  logic [0:0] f472_wen;
  logic [31:0] f472_wdata;
  logic [0:0] f472_clk;
  logic [0:0] f472_rst;
  logic [31:0] f472_rdata;
  sr_buffer_32_1 f472(.wen(f472_wen), .wdata(f472_wdata), .clk(f472_clk), .rst(f472_rst), .rdata(f472_rdata));
  assign f472_clk = clk;
  assign f472_rst = rst;
  // Bindings to f472

  // f474
  logic [0:0] f474_wen;
  logic [31:0] f474_wdata;
  logic [0:0] f474_clk;
  logic [0:0] f474_rst;
  logic [31:0] f474_rdata;
  sr_buffer_32_1 f474(.wen(f474_wen), .wdata(f474_wdata), .clk(f474_clk), .rst(f474_rst), .rdata(f474_rdata));
  assign f474_clk = clk;
  assign f474_rst = rst;
  // Bindings to f474

  // f476
  logic [0:0] f476_wen;
  logic [31:0] f476_wdata;
  logic [0:0] f476_clk;
  logic [0:0] f476_rst;
  logic [31:0] f476_rdata;
  sr_buffer_32_1 f476(.wen(f476_wen), .wdata(f476_wdata), .clk(f476_clk), .rst(f476_rst), .rdata(f476_rdata));
  assign f476_clk = clk;
  assign f476_rst = rst;
  // Bindings to f476

  // f478
  logic [0:0] f478_wen;
  logic [31:0] f478_wdata;
  logic [0:0] f478_clk;
  logic [0:0] f478_rst;
  logic [31:0] f478_rdata;
  sr_buffer_32_1 f478(.wen(f478_wen), .wdata(f478_wdata), .clk(f478_clk), .rst(f478_rst), .rdata(f478_rdata));
  assign f478_clk = clk;
  assign f478_rst = rst;
  // Bindings to f478

  // f480
  logic [0:0] f480_wen;
  logic [31:0] f480_wdata;
  logic [0:0] f480_clk;
  logic [0:0] f480_rst;
  logic [31:0] f480_rdata;
  sr_buffer_32_1 f480(.wen(f480_wen), .wdata(f480_wdata), .clk(f480_clk), .rst(f480_rst), .rdata(f480_rdata));
  assign f480_clk = clk;
  assign f480_rst = rst;
  // Bindings to f480

  // f482
  logic [0:0] f482_wen;
  logic [31:0] f482_wdata;
  logic [0:0] f482_clk;
  logic [0:0] f482_rst;
  logic [31:0] f482_rdata;
  sr_buffer_32_1 f482(.wen(f482_wen), .wdata(f482_wdata), .clk(f482_clk), .rst(f482_rst), .rdata(f482_rdata));
  assign f482_clk = clk;
  assign f482_rst = rst;
  // Bindings to f482

  // f484
  logic [0:0] f484_wen;
  logic [31:0] f484_wdata;
  logic [0:0] f484_clk;
  logic [0:0] f484_rst;
  logic [31:0] f484_rdata;
  sr_buffer_32_1 f484(.wen(f484_wen), .wdata(f484_wdata), .clk(f484_clk), .rst(f484_rst), .rdata(f484_rdata));
  assign f484_clk = clk;
  assign f484_rst = rst;
  // Bindings to f484

  // f486
  logic [0:0] f486_wen;
  logic [31:0] f486_wdata;
  logic [0:0] f486_clk;
  logic [0:0] f486_rst;
  logic [31:0] f486_rdata;
  sr_buffer_32_1 f486(.wen(f486_wen), .wdata(f486_wdata), .clk(f486_clk), .rst(f486_rst), .rdata(f486_rdata));
  assign f486_clk = clk;
  assign f486_rst = rst;
  // Bindings to f486

  // f488
  logic [0:0] f488_wen;
  logic [31:0] f488_wdata;
  logic [0:0] f488_clk;
  logic [0:0] f488_rst;
  logic [31:0] f488_rdata;
  sr_buffer_32_1 f488(.wen(f488_wen), .wdata(f488_wdata), .clk(f488_clk), .rst(f488_rst), .rdata(f488_rdata));
  assign f488_clk = clk;
  assign f488_rst = rst;
  // Bindings to f488

  // f490
  logic [0:0] f490_wen;
  logic [31:0] f490_wdata;
  logic [0:0] f490_clk;
  logic [0:0] f490_rst;
  logic [31:0] f490_rdata;
  sr_buffer_32_1 f490(.wen(f490_wen), .wdata(f490_wdata), .clk(f490_clk), .rst(f490_rst), .rdata(f490_rdata));
  assign f490_clk = clk;
  assign f490_rst = rst;
  // Bindings to f490

  // f492
  logic [0:0] f492_wen;
  logic [31:0] f492_wdata;
  logic [0:0] f492_clk;
  logic [0:0] f492_rst;
  logic [31:0] f492_rdata;
  sr_buffer_32_1 f492(.wen(f492_wen), .wdata(f492_wdata), .clk(f492_clk), .rst(f492_rst), .rdata(f492_rdata));
  assign f492_clk = clk;
  assign f492_rst = rst;
  // Bindings to f492

  // f494
  logic [0:0] f494_wen;
  logic [31:0] f494_wdata;
  logic [0:0] f494_clk;
  logic [0:0] f494_rst;
  logic [31:0] f494_rdata;
  sr_buffer_32_1 f494(.wen(f494_wen), .wdata(f494_wdata), .clk(f494_clk), .rst(f494_rst), .rdata(f494_rdata));
  assign f494_clk = clk;
  assign f494_rst = rst;
  // Bindings to f494

  // f496
  logic [0:0] f496_wen;
  logic [31:0] f496_wdata;
  logic [0:0] f496_clk;
  logic [0:0] f496_rst;
  logic [31:0] f496_rdata;
  sr_buffer_32_1 f496(.wen(f496_wen), .wdata(f496_wdata), .clk(f496_clk), .rst(f496_rst), .rdata(f496_rdata));
  assign f496_clk = clk;
  assign f496_rst = rst;
  // Bindings to f496

  // f498
  logic [0:0] f498_wen;
  logic [31:0] f498_wdata;
  logic [0:0] f498_clk;
  logic [0:0] f498_rst;
  logic [31:0] f498_rdata;
  sr_buffer_32_1 f498(.wen(f498_wen), .wdata(f498_wdata), .clk(f498_clk), .rst(f498_rst), .rdata(f498_rdata));
  assign f498_clk = clk;
  assign f498_rst = rst;
  // Bindings to f498

  // f500
  logic [0:0] f500_wen;
  logic [31:0] f500_wdata;
  logic [0:0] f500_clk;
  logic [0:0] f500_rst;
  logic [31:0] f500_rdata;
  sr_buffer_32_1 f500(.wen(f500_wen), .wdata(f500_wdata), .clk(f500_clk), .rst(f500_rst), .rdata(f500_rdata));
  assign f500_clk = clk;
  assign f500_rst = rst;
  // Bindings to f500

  // f502
  logic [0:0] f502_wen;
  logic [31:0] f502_wdata;
  logic [0:0] f502_clk;
  logic [0:0] f502_rst;
  logic [31:0] f502_rdata;
  sr_buffer_32_1 f502(.wen(f502_wen), .wdata(f502_wdata), .clk(f502_clk), .rst(f502_rst), .rdata(f502_rdata));
  assign f502_clk = clk;
  assign f502_rst = rst;
  // Bindings to f502

  // f504
  logic [0:0] f504_wen;
  logic [31:0] f504_wdata;
  logic [0:0] f504_clk;
  logic [0:0] f504_rst;
  logic [31:0] f504_rdata;
  sr_buffer_32_1 f504(.wen(f504_wen), .wdata(f504_wdata), .clk(f504_clk), .rst(f504_rst), .rdata(f504_rdata));
  assign f504_clk = clk;
  assign f504_rst = rst;
  // Bindings to f504

  // f506
  logic [0:0] f506_wen;
  logic [31:0] f506_wdata;
  logic [0:0] f506_clk;
  logic [0:0] f506_rst;
  logic [31:0] f506_rdata;
  sr_buffer_32_1 f506(.wen(f506_wen), .wdata(f506_wdata), .clk(f506_clk), .rst(f506_rst), .rdata(f506_rdata));
  assign f506_clk = clk;
  assign f506_rst = rst;
  // Bindings to f506

  // f508
  logic [0:0] f508_wen;
  logic [31:0] f508_wdata;
  logic [0:0] f508_clk;
  logic [0:0] f508_rst;
  logic [31:0] f508_rdata;
  sr_buffer_32_1 f508(.wen(f508_wen), .wdata(f508_wdata), .clk(f508_clk), .rst(f508_rst), .rdata(f508_rdata));
  assign f508_clk = clk;
  assign f508_rst = rst;
  // Bindings to f508

  // f510
  logic [0:0] f510_wen;
  logic [31:0] f510_wdata;
  logic [0:0] f510_clk;
  logic [0:0] f510_rst;
  logic [31:0] f510_rdata;
  sr_buffer_32_1 f510(.wen(f510_wen), .wdata(f510_wdata), .clk(f510_clk), .rst(f510_rst), .rdata(f510_rdata));
  assign f510_clk = clk;
  assign f510_rst = rst;
  // Bindings to f510

  // f512
  logic [0:0] f512_wen;
  logic [31:0] f512_wdata;
  logic [0:0] f512_clk;
  logic [0:0] f512_rst;
  logic [31:0] f512_rdata;
  sr_buffer_32_1 f512(.wen(f512_wen), .wdata(f512_wdata), .clk(f512_clk), .rst(f512_rst), .rdata(f512_rdata));
  assign f512_clk = clk;
  assign f512_rst = rst;
  // Bindings to f512

  // f514
  logic [0:0] f514_wen;
  logic [31:0] f514_wdata;
  logic [0:0] f514_clk;
  logic [0:0] f514_rst;
  logic [31:0] f514_rdata;
  sr_buffer_32_1 f514(.wen(f514_wen), .wdata(f514_wdata), .clk(f514_clk), .rst(f514_rst), .rdata(f514_rdata));
  assign f514_clk = clk;
  assign f514_rst = rst;
  // Bindings to f514

  // f516
  logic [0:0] f516_wen;
  logic [31:0] f516_wdata;
  logic [0:0] f516_clk;
  logic [0:0] f516_rst;
  logic [31:0] f516_rdata;
  sr_buffer_32_1 f516(.wen(f516_wen), .wdata(f516_wdata), .clk(f516_clk), .rst(f516_rst), .rdata(f516_rdata));
  assign f516_clk = clk;
  assign f516_rst = rst;
  // Bindings to f516

  // f518
  logic [0:0] f518_wen;
  logic [31:0] f518_wdata;
  logic [0:0] f518_clk;
  logic [0:0] f518_rst;
  logic [31:0] f518_rdata;
  sr_buffer_32_1 f518(.wen(f518_wen), .wdata(f518_wdata), .clk(f518_clk), .rst(f518_rst), .rdata(f518_rdata));
  assign f518_clk = clk;
  assign f518_rst = rst;
  // Bindings to f518

  // f520
  logic [0:0] f520_wen;
  logic [31:0] f520_wdata;
  logic [0:0] f520_clk;
  logic [0:0] f520_rst;
  logic [31:0] f520_rdata;
  sr_buffer_32_1 f520(.wen(f520_wen), .wdata(f520_wdata), .clk(f520_clk), .rst(f520_rst), .rdata(f520_rdata));
  assign f520_clk = clk;
  assign f520_rst = rst;
  // Bindings to f520

  // f522
  logic [0:0] f522_wen;
  logic [31:0] f522_wdata;
  logic [0:0] f522_clk;
  logic [0:0] f522_rst;
  logic [31:0] f522_rdata;
  sr_buffer_32_1 f522(.wen(f522_wen), .wdata(f522_wdata), .clk(f522_clk), .rst(f522_rst), .rdata(f522_rdata));
  assign f522_clk = clk;
  assign f522_rst = rst;
  // Bindings to f522

  // f524
  logic [0:0] f524_wen;
  logic [31:0] f524_wdata;
  logic [0:0] f524_clk;
  logic [0:0] f524_rst;
  logic [31:0] f524_rdata;
  sr_buffer_32_1 f524(.wen(f524_wen), .wdata(f524_wdata), .clk(f524_clk), .rst(f524_rst), .rdata(f524_rdata));
  assign f524_clk = clk;
  assign f524_rst = rst;
  // Bindings to f524

  // f526
  logic [0:0] f526_wen;
  logic [31:0] f526_wdata;
  logic [0:0] f526_clk;
  logic [0:0] f526_rst;
  logic [31:0] f526_rdata;
  sr_buffer_32_1 f526(.wen(f526_wen), .wdata(f526_wdata), .clk(f526_clk), .rst(f526_rst), .rdata(f526_rdata));
  assign f526_clk = clk;
  assign f526_rst = rst;
  // Bindings to f526

  // f528
  logic [0:0] f528_wen;
  logic [31:0] f528_wdata;
  logic [0:0] f528_clk;
  logic [0:0] f528_rst;
  logic [31:0] f528_rdata;
  sr_buffer_32_1 f528(.wen(f528_wen), .wdata(f528_wdata), .clk(f528_clk), .rst(f528_rst), .rdata(f528_rdata));
  assign f528_clk = clk;
  assign f528_rst = rst;
  // Bindings to f528

  // f530
  logic [0:0] f530_wen;
  logic [31:0] f530_wdata;
  logic [0:0] f530_clk;
  logic [0:0] f530_rst;
  logic [31:0] f530_rdata;
  sr_buffer_32_1 f530(.wen(f530_wen), .wdata(f530_wdata), .clk(f530_clk), .rst(f530_rst), .rdata(f530_rdata));
  assign f530_clk = clk;
  assign f530_rst = rst;
  // Bindings to f530

  // f532
  logic [0:0] f532_wen;
  logic [31:0] f532_wdata;
  logic [0:0] f532_clk;
  logic [0:0] f532_rst;
  logic [31:0] f532_rdata;
  sr_buffer_32_1 f532(.wen(f532_wen), .wdata(f532_wdata), .clk(f532_clk), .rst(f532_rst), .rdata(f532_rdata));
  assign f532_clk = clk;
  assign f532_rst = rst;
  // Bindings to f532

  // f534
  logic [0:0] f534_wen;
  logic [31:0] f534_wdata;
  logic [0:0] f534_clk;
  logic [0:0] f534_rst;
  logic [31:0] f534_rdata;
  sr_buffer_32_1 f534(.wen(f534_wen), .wdata(f534_wdata), .clk(f534_clk), .rst(f534_rst), .rdata(f534_rdata));
  assign f534_clk = clk;
  assign f534_rst = rst;
  // Bindings to f534

  // f536
  logic [0:0] f536_wen;
  logic [31:0] f536_wdata;
  logic [0:0] f536_clk;
  logic [0:0] f536_rst;
  logic [31:0] f536_rdata;
  sr_buffer_32_1 f536(.wen(f536_wen), .wdata(f536_wdata), .clk(f536_clk), .rst(f536_rst), .rdata(f536_rdata));
  assign f536_clk = clk;
  assign f536_rst = rst;
  // Bindings to f536

  // f538
  logic [0:0] f538_wen;
  logic [31:0] f538_wdata;
  logic [0:0] f538_clk;
  logic [0:0] f538_rst;
  logic [31:0] f538_rdata;
  sr_buffer_32_1 f538(.wen(f538_wen), .wdata(f538_wdata), .clk(f538_clk), .rst(f538_rst), .rdata(f538_rdata));
  assign f538_clk = clk;
  assign f538_rst = rst;
  // Bindings to f538

  // f540
  logic [0:0] f540_wen;
  logic [31:0] f540_wdata;
  logic [0:0] f540_clk;
  logic [0:0] f540_rst;
  logic [31:0] f540_rdata;
  sr_buffer_32_1 f540(.wen(f540_wen), .wdata(f540_wdata), .clk(f540_clk), .rst(f540_rst), .rdata(f540_rdata));
  assign f540_clk = clk;
  assign f540_rst = rst;
  // Bindings to f540

  // f542
  logic [0:0] f542_wen;
  logic [31:0] f542_wdata;
  logic [0:0] f542_clk;
  logic [0:0] f542_rst;
  logic [31:0] f542_rdata;
  sr_buffer_32_1 f542(.wen(f542_wen), .wdata(f542_wdata), .clk(f542_clk), .rst(f542_rst), .rdata(f542_rdata));
  assign f542_clk = clk;
  assign f542_rst = rst;
  // Bindings to f542

  // f544
  logic [0:0] f544_wen;
  logic [31:0] f544_wdata;
  logic [0:0] f544_clk;
  logic [0:0] f544_rst;
  logic [31:0] f544_rdata;
  sr_buffer_32_1 f544(.wen(f544_wen), .wdata(f544_wdata), .clk(f544_clk), .rst(f544_rst), .rdata(f544_rdata));
  assign f544_clk = clk;
  assign f544_rst = rst;
  // Bindings to f544

  // f546
  logic [0:0] f546_wen;
  logic [31:0] f546_wdata;
  logic [0:0] f546_clk;
  logic [0:0] f546_rst;
  logic [31:0] f546_rdata;
  sr_buffer_32_1 f546(.wen(f546_wen), .wdata(f546_wdata), .clk(f546_clk), .rst(f546_rst), .rdata(f546_rdata));
  assign f546_clk = clk;
  assign f546_rst = rst;
  // Bindings to f546

  // f548
  logic [0:0] f548_wen;
  logic [31:0] f548_wdata;
  logic [0:0] f548_clk;
  logic [0:0] f548_rst;
  logic [31:0] f548_rdata;
  sr_buffer_32_1 f548(.wen(f548_wen), .wdata(f548_wdata), .clk(f548_clk), .rst(f548_rst), .rdata(f548_rdata));
  assign f548_clk = clk;
  assign f548_rst = rst;
  // Bindings to f548

  // f550
  logic [0:0] f550_wen;
  logic [31:0] f550_wdata;
  logic [0:0] f550_clk;
  logic [0:0] f550_rst;
  logic [31:0] f550_rdata;
  sr_buffer_32_1 f550(.wen(f550_wen), .wdata(f550_wdata), .clk(f550_clk), .rst(f550_rst), .rdata(f550_rdata));
  assign f550_clk = clk;
  assign f550_rst = rst;
  // Bindings to f550

  // f552
  logic [0:0] f552_wen;
  logic [31:0] f552_wdata;
  logic [0:0] f552_clk;
  logic [0:0] f552_rst;
  logic [31:0] f552_rdata;
  sr_buffer_32_1 f552(.wen(f552_wen), .wdata(f552_wdata), .clk(f552_clk), .rst(f552_rst), .rdata(f552_rdata));
  assign f552_clk = clk;
  assign f552_rst = rst;
  // Bindings to f552

  // f554
  logic [0:0] f554_wen;
  logic [31:0] f554_wdata;
  logic [0:0] f554_clk;
  logic [0:0] f554_rst;
  logic [31:0] f554_rdata;
  sr_buffer_32_1 f554(.wen(f554_wen), .wdata(f554_wdata), .clk(f554_clk), .rst(f554_rst), .rdata(f554_rdata));
  assign f554_clk = clk;
  assign f554_rst = rst;
  // Bindings to f554

  // f556
  logic [0:0] f556_wen;
  logic [31:0] f556_wdata;
  logic [0:0] f556_clk;
  logic [0:0] f556_rst;
  logic [31:0] f556_rdata;
  sr_buffer_32_1 f556(.wen(f556_wen), .wdata(f556_wdata), .clk(f556_clk), .rst(f556_rst), .rdata(f556_rdata));
  assign f556_clk = clk;
  assign f556_rst = rst;
  // Bindings to f556

  // f558
  logic [0:0] f558_wen;
  logic [31:0] f558_wdata;
  logic [0:0] f558_clk;
  logic [0:0] f558_rst;
  logic [31:0] f558_rdata;
  sr_buffer_32_1 f558(.wen(f558_wen), .wdata(f558_wdata), .clk(f558_clk), .rst(f558_rst), .rdata(f558_rdata));
  assign f558_clk = clk;
  assign f558_rst = rst;
  // Bindings to f558

  // f560
  logic [0:0] f560_wen;
  logic [31:0] f560_wdata;
  logic [0:0] f560_clk;
  logic [0:0] f560_rst;
  logic [31:0] f560_rdata;
  sr_buffer_32_1 f560(.wen(f560_wen), .wdata(f560_wdata), .clk(f560_clk), .rst(f560_rst), .rdata(f560_rdata));
  assign f560_clk = clk;
  assign f560_rst = rst;
  // Bindings to f560

  // f562
  logic [0:0] f562_wen;
  logic [31:0] f562_wdata;
  logic [0:0] f562_clk;
  logic [0:0] f562_rst;
  logic [31:0] f562_rdata;
  sr_buffer_32_1 f562(.wen(f562_wen), .wdata(f562_wdata), .clk(f562_clk), .rst(f562_rst), .rdata(f562_rdata));
  assign f562_clk = clk;
  assign f562_rst = rst;
  // Bindings to f562

  // f564
  logic [0:0] f564_wen;
  logic [31:0] f564_wdata;
  logic [0:0] f564_clk;
  logic [0:0] f564_rst;
  logic [31:0] f564_rdata;
  sr_buffer_32_1 f564(.wen(f564_wen), .wdata(f564_wdata), .clk(f564_clk), .rst(f564_rst), .rdata(f564_rdata));
  assign f564_clk = clk;
  assign f564_rst = rst;
  // Bindings to f564

  // f566
  logic [0:0] f566_wen;
  logic [31:0] f566_wdata;
  logic [0:0] f566_clk;
  logic [0:0] f566_rst;
  logic [31:0] f566_rdata;
  sr_buffer_32_1 f566(.wen(f566_wen), .wdata(f566_wdata), .clk(f566_clk), .rst(f566_rst), .rdata(f566_rdata));
  assign f566_clk = clk;
  assign f566_rst = rst;
  // Bindings to f566

  // f568
  logic [0:0] f568_wen;
  logic [31:0] f568_wdata;
  logic [0:0] f568_clk;
  logic [0:0] f568_rst;
  logic [31:0] f568_rdata;
  sr_buffer_32_1 f568(.wen(f568_wen), .wdata(f568_wdata), .clk(f568_clk), .rst(f568_rst), .rdata(f568_rdata));
  assign f568_clk = clk;
  assign f568_rst = rst;
  // Bindings to f568

  // f570
  logic [0:0] f570_wen;
  logic [31:0] f570_wdata;
  logic [0:0] f570_clk;
  logic [0:0] f570_rst;
  logic [31:0] f570_rdata;
  sr_buffer_32_1 f570(.wen(f570_wen), .wdata(f570_wdata), .clk(f570_clk), .rst(f570_rst), .rdata(f570_rdata));
  assign f570_clk = clk;
  assign f570_rst = rst;
  // Bindings to f570

  // f572
  logic [0:0] f572_wen;
  logic [31:0] f572_wdata;
  logic [0:0] f572_clk;
  logic [0:0] f572_rst;
  logic [31:0] f572_rdata;
  sr_buffer_32_1 f572(.wen(f572_wen), .wdata(f572_wdata), .clk(f572_clk), .rst(f572_rst), .rdata(f572_rdata));
  assign f572_clk = clk;
  assign f572_rst = rst;
  // Bindings to f572

  // f574
  logic [0:0] f574_wen;
  logic [31:0] f574_wdata;
  logic [0:0] f574_clk;
  logic [0:0] f574_rst;
  logic [31:0] f574_rdata;
  sr_buffer_32_1 f574(.wen(f574_wen), .wdata(f574_wdata), .clk(f574_clk), .rst(f574_rst), .rdata(f574_rdata));
  assign f574_clk = clk;
  assign f574_rst = rst;
  // Bindings to f574

  // f576
  logic [0:0] f576_wen;
  logic [31:0] f576_wdata;
  logic [0:0] f576_clk;
  logic [0:0] f576_rst;
  logic [31:0] f576_rdata;
  sr_buffer_32_1 f576(.wen(f576_wen), .wdata(f576_wdata), .clk(f576_clk), .rst(f576_rst), .rdata(f576_rdata));
  assign f576_clk = clk;
  assign f576_rst = rst;
  // Bindings to f576

  // f578
  logic [0:0] f578_wen;
  logic [31:0] f578_wdata;
  logic [0:0] f578_clk;
  logic [0:0] f578_rst;
  logic [31:0] f578_rdata;
  sr_buffer_32_1 f578(.wen(f578_wen), .wdata(f578_wdata), .clk(f578_clk), .rst(f578_rst), .rdata(f578_rdata));
  assign f578_clk = clk;
  assign f578_rst = rst;
  // Bindings to f578

  // f580
  logic [0:0] f580_wen;
  logic [31:0] f580_wdata;
  logic [0:0] f580_clk;
  logic [0:0] f580_rst;
  logic [31:0] f580_rdata;
  sr_buffer_32_1 f580(.wen(f580_wen), .wdata(f580_wdata), .clk(f580_clk), .rst(f580_rst), .rdata(f580_rdata));
  assign f580_clk = clk;
  assign f580_rst = rst;
  // Bindings to f580

  // f582
  logic [0:0] f582_wen;
  logic [31:0] f582_wdata;
  logic [0:0] f582_clk;
  logic [0:0] f582_rst;
  logic [31:0] f582_rdata;
  sr_buffer_32_1 f582(.wen(f582_wen), .wdata(f582_wdata), .clk(f582_clk), .rst(f582_rst), .rdata(f582_rdata));
  assign f582_clk = clk;
  assign f582_rst = rst;
  // Bindings to f582

  // f584
  logic [0:0] f584_wen;
  logic [31:0] f584_wdata;
  logic [0:0] f584_clk;
  logic [0:0] f584_rst;
  logic [31:0] f584_rdata;
  sr_buffer_32_1 f584(.wen(f584_wen), .wdata(f584_wdata), .clk(f584_clk), .rst(f584_rst), .rdata(f584_rdata));
  assign f584_clk = clk;
  assign f584_rst = rst;
  // Bindings to f584

  // f586
  logic [0:0] f586_wen;
  logic [31:0] f586_wdata;
  logic [0:0] f586_clk;
  logic [0:0] f586_rst;
  logic [31:0] f586_rdata;
  sr_buffer_32_1 f586(.wen(f586_wen), .wdata(f586_wdata), .clk(f586_clk), .rst(f586_rst), .rdata(f586_rdata));
  assign f586_clk = clk;
  assign f586_rst = rst;
  // Bindings to f586

  // f588
  logic [0:0] f588_wen;
  logic [31:0] f588_wdata;
  logic [0:0] f588_clk;
  logic [0:0] f588_rst;
  logic [31:0] f588_rdata;
  sr_buffer_32_1 f588(.wen(f588_wen), .wdata(f588_wdata), .clk(f588_clk), .rst(f588_rst), .rdata(f588_rdata));
  assign f588_clk = clk;
  assign f588_rst = rst;
  // Bindings to f588

  // f590
  logic [0:0] f590_wen;
  logic [31:0] f590_wdata;
  logic [0:0] f590_clk;
  logic [0:0] f590_rst;
  logic [31:0] f590_rdata;
  sr_buffer_32_1 f590(.wen(f590_wen), .wdata(f590_wdata), .clk(f590_clk), .rst(f590_rst), .rdata(f590_rdata));
  assign f590_clk = clk;
  assign f590_rst = rst;
  // Bindings to f590

  // f592
  logic [0:0] f592_wen;
  logic [31:0] f592_wdata;
  logic [0:0] f592_clk;
  logic [0:0] f592_rst;
  logic [31:0] f592_rdata;
  sr_buffer_32_1 f592(.wen(f592_wen), .wdata(f592_wdata), .clk(f592_clk), .rst(f592_rst), .rdata(f592_rdata));
  assign f592_clk = clk;
  assign f592_rst = rst;
  // Bindings to f592

  // f594
  logic [0:0] f594_wen;
  logic [31:0] f594_wdata;
  logic [0:0] f594_clk;
  logic [0:0] f594_rst;
  logic [31:0] f594_rdata;
  sr_buffer_32_1 f594(.wen(f594_wen), .wdata(f594_wdata), .clk(f594_clk), .rst(f594_rst), .rdata(f594_rdata));
  assign f594_clk = clk;
  assign f594_rst = rst;
  // Bindings to f594

  // f596
  logic [0:0] f596_wen;
  logic [31:0] f596_wdata;
  logic [0:0] f596_clk;
  logic [0:0] f596_rst;
  logic [31:0] f596_rdata;
  sr_buffer_32_1 f596(.wen(f596_wen), .wdata(f596_wdata), .clk(f596_clk), .rst(f596_rst), .rdata(f596_rdata));
  assign f596_clk = clk;
  assign f596_rst = rst;
  // Bindings to f596

  // f598
  logic [0:0] f598_wen;
  logic [31:0] f598_wdata;
  logic [0:0] f598_clk;
  logic [0:0] f598_rst;
  logic [31:0] f598_rdata;
  sr_buffer_32_1 f598(.wen(f598_wen), .wdata(f598_wdata), .clk(f598_clk), .rst(f598_rst), .rdata(f598_rdata));
  assign f598_clk = clk;
  assign f598_rst = rst;
  // Bindings to f598

  // f600
  logic [0:0] f600_wen;
  logic [31:0] f600_wdata;
  logic [0:0] f600_clk;
  logic [0:0] f600_rst;
  logic [31:0] f600_rdata;
  sr_buffer_32_1 f600(.wen(f600_wen), .wdata(f600_wdata), .clk(f600_clk), .rst(f600_rst), .rdata(f600_rdata));
  assign f600_clk = clk;
  assign f600_rst = rst;
  // Bindings to f600

  // f602
  logic [0:0] f602_wen;
  logic [31:0] f602_wdata;
  logic [0:0] f602_clk;
  logic [0:0] f602_rst;
  logic [31:0] f602_rdata;
  sr_buffer_32_1 f602(.wen(f602_wen), .wdata(f602_wdata), .clk(f602_clk), .rst(f602_rst), .rdata(f602_rdata));
  assign f602_clk = clk;
  assign f602_rst = rst;
  // Bindings to f602

  // f604
  logic [0:0] f604_wen;
  logic [31:0] f604_wdata;
  logic [0:0] f604_clk;
  logic [0:0] f604_rst;
  logic [31:0] f604_rdata;
  sr_buffer_32_1 f604(.wen(f604_wen), .wdata(f604_wdata), .clk(f604_clk), .rst(f604_rst), .rdata(f604_rdata));
  assign f604_clk = clk;
  assign f604_rst = rst;
  // Bindings to f604

  // f606
  logic [0:0] f606_wen;
  logic [31:0] f606_wdata;
  logic [0:0] f606_clk;
  logic [0:0] f606_rst;
  logic [31:0] f606_rdata;
  sr_buffer_32_1 f606(.wen(f606_wen), .wdata(f606_wdata), .clk(f606_clk), .rst(f606_rst), .rdata(f606_rdata));
  assign f606_clk = clk;
  assign f606_rst = rst;
  // Bindings to f606

  // f608
  logic [0:0] f608_wen;
  logic [31:0] f608_wdata;
  logic [0:0] f608_clk;
  logic [0:0] f608_rst;
  logic [31:0] f608_rdata;
  sr_buffer_32_1 f608(.wen(f608_wen), .wdata(f608_wdata), .clk(f608_clk), .rst(f608_rst), .rdata(f608_rdata));
  assign f608_clk = clk;
  assign f608_rst = rst;
  // Bindings to f608

  // f610
  logic [0:0] f610_wen;
  logic [31:0] f610_wdata;
  logic [0:0] f610_clk;
  logic [0:0] f610_rst;
  logic [31:0] f610_rdata;
  sr_buffer_32_1 f610(.wen(f610_wen), .wdata(f610_wdata), .clk(f610_clk), .rst(f610_rst), .rdata(f610_rdata));
  assign f610_clk = clk;
  assign f610_rst = rst;
  // Bindings to f610

  // f612
  logic [0:0] f612_wen;
  logic [31:0] f612_wdata;
  logic [0:0] f612_clk;
  logic [0:0] f612_rst;
  logic [31:0] f612_rdata;
  sr_buffer_32_1 f612(.wen(f612_wen), .wdata(f612_wdata), .clk(f612_clk), .rst(f612_rst), .rdata(f612_rdata));
  assign f612_clk = clk;
  assign f612_rst = rst;
  // Bindings to f612

  // f614
  logic [0:0] f614_wen;
  logic [31:0] f614_wdata;
  logic [0:0] f614_clk;
  logic [0:0] f614_rst;
  logic [31:0] f614_rdata;
  sr_buffer_32_1 f614(.wen(f614_wen), .wdata(f614_wdata), .clk(f614_clk), .rst(f614_rst), .rdata(f614_rdata));
  assign f614_clk = clk;
  assign f614_rst = rst;
  // Bindings to f614

  // f616
  logic [0:0] f616_wen;
  logic [31:0] f616_wdata;
  logic [0:0] f616_clk;
  logic [0:0] f616_rst;
  logic [31:0] f616_rdata;
  sr_buffer_32_1 f616(.wen(f616_wen), .wdata(f616_wdata), .clk(f616_clk), .rst(f616_rst), .rdata(f616_rdata));
  assign f616_clk = clk;
  assign f616_rst = rst;
  // Bindings to f616

  // f618
  logic [0:0] f618_wen;
  logic [31:0] f618_wdata;
  logic [0:0] f618_clk;
  logic [0:0] f618_rst;
  logic [31:0] f618_rdata;
  sr_buffer_32_1 f618(.wen(f618_wen), .wdata(f618_wdata), .clk(f618_clk), .rst(f618_rst), .rdata(f618_rdata));
  assign f618_clk = clk;
  assign f618_rst = rst;
  // Bindings to f618

  // f620
  logic [0:0] f620_wen;
  logic [31:0] f620_wdata;
  logic [0:0] f620_clk;
  logic [0:0] f620_rst;
  logic [31:0] f620_rdata;
  sr_buffer_32_1 f620(.wen(f620_wen), .wdata(f620_wdata), .clk(f620_clk), .rst(f620_rst), .rdata(f620_rdata));
  assign f620_clk = clk;
  assign f620_rst = rst;
  // Bindings to f620

  // f622
  logic [0:0] f622_wen;
  logic [31:0] f622_wdata;
  logic [0:0] f622_clk;
  logic [0:0] f622_rst;
  logic [31:0] f622_rdata;
  sr_buffer_32_1 f622(.wen(f622_wen), .wdata(f622_wdata), .clk(f622_clk), .rst(f622_rst), .rdata(f622_rdata));
  assign f622_clk = clk;
  assign f622_rst = rst;
  // Bindings to f622

  // f624
  logic [0:0] f624_wen;
  logic [31:0] f624_wdata;
  logic [0:0] f624_clk;
  logic [0:0] f624_rst;
  logic [31:0] f624_rdata;
  sr_buffer_32_1 f624(.wen(f624_wen), .wdata(f624_wdata), .clk(f624_clk), .rst(f624_rst), .rdata(f624_rdata));
  assign f624_clk = clk;
  assign f624_rst = rst;
  // Bindings to f624

  // f626
  logic [0:0] f626_wen;
  logic [31:0] f626_wdata;
  logic [0:0] f626_clk;
  logic [0:0] f626_rst;
  logic [31:0] f626_rdata;
  sr_buffer_32_1 f626(.wen(f626_wen), .wdata(f626_wdata), .clk(f626_clk), .rst(f626_rst), .rdata(f626_rdata));
  assign f626_clk = clk;
  assign f626_rst = rst;
  // Bindings to f626

  // f628
  logic [0:0] f628_wen;
  logic [31:0] f628_wdata;
  logic [0:0] f628_clk;
  logic [0:0] f628_rst;
  logic [31:0] f628_rdata;
  sr_buffer_32_1 f628(.wen(f628_wen), .wdata(f628_wdata), .clk(f628_clk), .rst(f628_rst), .rdata(f628_rdata));
  assign f628_clk = clk;
  assign f628_rst = rst;
  // Bindings to f628

  // f630
  logic [0:0] f630_wen;
  logic [31:0] f630_wdata;
  logic [0:0] f630_clk;
  logic [0:0] f630_rst;
  logic [31:0] f630_rdata;
  sr_buffer_32_1 f630(.wen(f630_wen), .wdata(f630_wdata), .clk(f630_clk), .rst(f630_rst), .rdata(f630_rdata));
  assign f630_clk = clk;
  assign f630_rst = rst;
  // Bindings to f630

  // f632
  logic [0:0] f632_wen;
  logic [31:0] f632_wdata;
  logic [0:0] f632_clk;
  logic [0:0] f632_rst;
  logic [31:0] f632_rdata;
  sr_buffer_32_1 f632(.wen(f632_wen), .wdata(f632_wdata), .clk(f632_clk), .rst(f632_rst), .rdata(f632_rdata));
  assign f632_clk = clk;
  assign f632_rst = rst;
  // Bindings to f632

  // f634
  logic [0:0] f634_wen;
  logic [31:0] f634_wdata;
  logic [0:0] f634_clk;
  logic [0:0] f634_rst;
  logic [31:0] f634_rdata;
  sr_buffer_32_1 f634(.wen(f634_wen), .wdata(f634_wdata), .clk(f634_clk), .rst(f634_rst), .rdata(f634_rdata));
  assign f634_clk = clk;
  assign f634_rst = rst;
  // Bindings to f634

  // f636
  logic [0:0] f636_wen;
  logic [31:0] f636_wdata;
  logic [0:0] f636_clk;
  logic [0:0] f636_rst;
  logic [31:0] f636_rdata;
  sr_buffer_32_1 f636(.wen(f636_wen), .wdata(f636_wdata), .clk(f636_clk), .rst(f636_rst), .rdata(f636_rdata));
  assign f636_clk = clk;
  assign f636_rst = rst;
  // Bindings to f636

  // f638
  logic [0:0] f638_wen;
  logic [31:0] f638_wdata;
  logic [0:0] f638_clk;
  logic [0:0] f638_rst;
  logic [31:0] f638_rdata;
  sr_buffer_32_1 f638(.wen(f638_wen), .wdata(f638_wdata), .clk(f638_clk), .rst(f638_rst), .rdata(f638_rdata));
  assign f638_clk = clk;
  assign f638_rst = rst;
  // Bindings to f638

  // f640
  logic [0:0] f640_wen;
  logic [31:0] f640_wdata;
  logic [0:0] f640_clk;
  logic [0:0] f640_rst;
  logic [31:0] f640_rdata;
  sr_buffer_32_1 f640(.wen(f640_wen), .wdata(f640_wdata), .clk(f640_clk), .rst(f640_rst), .rdata(f640_rdata));
  assign f640_clk = clk;
  assign f640_rst = rst;
  // Bindings to f640

  // f642
  logic [0:0] f642_wen;
  logic [31:0] f642_wdata;
  logic [0:0] f642_clk;
  logic [0:0] f642_rst;
  logic [31:0] f642_rdata;
  sr_buffer_32_1 f642(.wen(f642_wen), .wdata(f642_wdata), .clk(f642_clk), .rst(f642_rst), .rdata(f642_rdata));
  assign f642_clk = clk;
  assign f642_rst = rst;
  // Bindings to f642

  // f644
  logic [0:0] f644_wen;
  logic [31:0] f644_wdata;
  logic [0:0] f644_clk;
  logic [0:0] f644_rst;
  logic [31:0] f644_rdata;
  sr_buffer_32_1 f644(.wen(f644_wen), .wdata(f644_wdata), .clk(f644_clk), .rst(f644_rst), .rdata(f644_rdata));
  assign f644_clk = clk;
  assign f644_rst = rst;
  // Bindings to f644

  // f646
  logic [0:0] f646_wen;
  logic [31:0] f646_wdata;
  logic [0:0] f646_clk;
  logic [0:0] f646_rst;
  logic [31:0] f646_rdata;
  sr_buffer_32_1 f646(.wen(f646_wen), .wdata(f646_wdata), .clk(f646_clk), .rst(f646_rst), .rdata(f646_rdata));
  assign f646_clk = clk;
  assign f646_rst = rst;
  // Bindings to f646

  // f648
  logic [0:0] f648_wen;
  logic [31:0] f648_wdata;
  logic [0:0] f648_clk;
  logic [0:0] f648_rst;
  logic [31:0] f648_rdata;
  sr_buffer_32_1 f648(.wen(f648_wen), .wdata(f648_wdata), .clk(f648_clk), .rst(f648_rst), .rdata(f648_rdata));
  assign f648_clk = clk;
  assign f648_rst = rst;
  // Bindings to f648

  // f650
  logic [0:0] f650_wen;
  logic [31:0] f650_wdata;
  logic [0:0] f650_clk;
  logic [0:0] f650_rst;
  logic [31:0] f650_rdata;
  sr_buffer_32_1 f650(.wen(f650_wen), .wdata(f650_wdata), .clk(f650_clk), .rst(f650_rst), .rdata(f650_rdata));
  assign f650_clk = clk;
  assign f650_rst = rst;
  // Bindings to f650

  // f652
  logic [0:0] f652_wen;
  logic [31:0] f652_wdata;
  logic [0:0] f652_clk;
  logic [0:0] f652_rst;
  logic [31:0] f652_rdata;
  sr_buffer_32_1 f652(.wen(f652_wen), .wdata(f652_wdata), .clk(f652_clk), .rst(f652_rst), .rdata(f652_rdata));
  assign f652_clk = clk;
  assign f652_rst = rst;
  // Bindings to f652

  // f654
  logic [0:0] f654_wen;
  logic [31:0] f654_wdata;
  logic [0:0] f654_clk;
  logic [0:0] f654_rst;
  logic [31:0] f654_rdata;
  sr_buffer_32_1 f654(.wen(f654_wen), .wdata(f654_wdata), .clk(f654_clk), .rst(f654_rst), .rdata(f654_rdata));
  assign f654_clk = clk;
  assign f654_rst = rst;
  // Bindings to f654

  // f656
  logic [0:0] f656_wen;
  logic [31:0] f656_wdata;
  logic [0:0] f656_clk;
  logic [0:0] f656_rst;
  logic [31:0] f656_rdata;
  sr_buffer_32_1 f656(.wen(f656_wen), .wdata(f656_wdata), .clk(f656_clk), .rst(f656_rst), .rdata(f656_rdata));
  assign f656_clk = clk;
  assign f656_rst = rst;
  // Bindings to f656

  // f658
  logic [0:0] f658_wen;
  logic [31:0] f658_wdata;
  logic [0:0] f658_clk;
  logic [0:0] f658_rst;
  logic [31:0] f658_rdata;
  sr_buffer_32_1 f658(.wen(f658_wen), .wdata(f658_wdata), .clk(f658_clk), .rst(f658_rst), .rdata(f658_rdata));
  assign f658_clk = clk;
  assign f658_rst = rst;
  // Bindings to f658

  // f660
  logic [0:0] f660_wen;
  logic [31:0] f660_wdata;
  logic [0:0] f660_clk;
  logic [0:0] f660_rst;
  logic [31:0] f660_rdata;
  sr_buffer_32_1 f660(.wen(f660_wen), .wdata(f660_wdata), .clk(f660_clk), .rst(f660_rst), .rdata(f660_rdata));
  assign f660_clk = clk;
  assign f660_rst = rst;
  // Bindings to f660

  // f662
  logic [0:0] f662_wen;
  logic [31:0] f662_wdata;
  logic [0:0] f662_clk;
  logic [0:0] f662_rst;
  logic [31:0] f662_rdata;
  sr_buffer_32_1 f662(.wen(f662_wen), .wdata(f662_wdata), .clk(f662_clk), .rst(f662_rst), .rdata(f662_rdata));
  assign f662_clk = clk;
  assign f662_rst = rst;
  // Bindings to f662

  // f664
  logic [0:0] f664_wen;
  logic [31:0] f664_wdata;
  logic [0:0] f664_clk;
  logic [0:0] f664_rst;
  logic [31:0] f664_rdata;
  sr_buffer_32_1 f664(.wen(f664_wen), .wdata(f664_wdata), .clk(f664_clk), .rst(f664_rst), .rdata(f664_rdata));
  assign f664_clk = clk;
  assign f664_rst = rst;
  // Bindings to f664

  // f666
  logic [0:0] f666_wen;
  logic [31:0] f666_wdata;
  logic [0:0] f666_clk;
  logic [0:0] f666_rst;
  logic [31:0] f666_rdata;
  sr_buffer_32_1 f666(.wen(f666_wen), .wdata(f666_wdata), .clk(f666_clk), .rst(f666_rst), .rdata(f666_rdata));
  assign f666_clk = clk;
  assign f666_rst = rst;
  // Bindings to f666

  // f668
  logic [0:0] f668_wen;
  logic [31:0] f668_wdata;
  logic [0:0] f668_clk;
  logic [0:0] f668_rst;
  logic [31:0] f668_rdata;
  sr_buffer_32_1 f668(.wen(f668_wen), .wdata(f668_wdata), .clk(f668_clk), .rst(f668_rst), .rdata(f668_rdata));
  assign f668_clk = clk;
  assign f668_rst = rst;
  // Bindings to f668

  // f670
  logic [0:0] f670_wen;
  logic [31:0] f670_wdata;
  logic [0:0] f670_clk;
  logic [0:0] f670_rst;
  logic [31:0] f670_rdata;
  sr_buffer_32_1 f670(.wen(f670_wen), .wdata(f670_wdata), .clk(f670_clk), .rst(f670_rst), .rdata(f670_rdata));
  assign f670_clk = clk;
  assign f670_rst = rst;
  // Bindings to f670

  // f672
  logic [0:0] f672_wen;
  logic [31:0] f672_wdata;
  logic [0:0] f672_clk;
  logic [0:0] f672_rst;
  logic [31:0] f672_rdata;
  sr_buffer_32_1 f672(.wen(f672_wen), .wdata(f672_wdata), .clk(f672_clk), .rst(f672_rst), .rdata(f672_rdata));
  assign f672_clk = clk;
  assign f672_rst = rst;
  // Bindings to f672

  // f674
  logic [0:0] f674_wen;
  logic [31:0] f674_wdata;
  logic [0:0] f674_clk;
  logic [0:0] f674_rst;
  logic [31:0] f674_rdata;
  sr_buffer_32_1 f674(.wen(f674_wen), .wdata(f674_wdata), .clk(f674_clk), .rst(f674_rst), .rdata(f674_rdata));
  assign f674_clk = clk;
  assign f674_rst = rst;
  // Bindings to f674



endmodule


module in_wire_dark_update_0_write_wdata(output [31:0] dark_update_0_write_wdata);

endmodule


module dark_weights_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_gauss_blur_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_gauss_blur_1_update_0_write_wen, input [31:0] dark_gauss_ds_1_update_0_read_dummy, input [31:0] dark_gauss_blur_1_update_0_write_wdata, output [31:0] dark_gauss_ds_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // selector_dark_gauss_ds_1_rd0_select
  logic [0:0] selector_dark_gauss_ds_1_rd0_select_clk;
  logic [0:0] selector_dark_gauss_ds_1_rd0_select_rst;
  logic [31:0] selector_dark_gauss_ds_1_rd0_select_d0;
  logic [31:0] selector_dark_gauss_ds_1_rd0_select_d1;
  logic [31:0] selector_dark_gauss_ds_1_rd0_select_out;
  dark_gauss_ds_1_rd0_select selector_dark_gauss_ds_1_rd0_select(.clk(selector_dark_gauss_ds_1_rd0_select_clk), .rst(selector_dark_gauss_ds_1_rd0_select_rst), .d0(selector_dark_gauss_ds_1_rd0_select_d0), .d1(selector_dark_gauss_ds_1_rd0_select_d1), .out(selector_dark_gauss_ds_1_rd0_select_out));
  assign selector_dark_gauss_ds_1_rd0_select_clk = clk;
  assign selector_dark_gauss_ds_1_rd0_select_rst = rst;
  // Bindings to selector_dark_gauss_ds_1_rd0_select

  // Bindings to dark_gauss_blur_1_update_0_write_wen
    // rd_0
  assign rd_0 = dark_gauss_blur_1_update_0_write_wen;

  // Bindings to dark_gauss_ds_1_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_gauss_ds_1_update_0_read_dummy;

  // dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1
  logic [0:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_done;
  dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1 dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1(.clk(dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_clk), .rst(dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_rst), .start(dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_start), .done(dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_done));
  assign dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_clk = clk;
  assign dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1

  // Bindings to dark_gauss_blur_1_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_gauss_blur_1_update_0_write_wdata;

  // Bindings to dark_gauss_ds_1_update_0_read_rdata
    // wr_3
  assign dark_gauss_ds_1_update_0_read_rdata = rd_2;



endmodule


module in_wire_dark_gauss_blur_1_update_0_read_dummy(output [287:0] dark_gauss_blur_1_update_0_read_dummy);

endmodule


module out_wire_dark_gauss_blur_1_update_0_read_rdata(input [287:0] dark_gauss_blur_1_update_0_read_rdata);

endmodule


module in_wire_dark_laplace_diff_0_update_0_read_dummy(output [31:0] dark_laplace_diff_0_update_0_read_dummy);

endmodule


module out_wire_dark_laplace_diff_0_update_0_read_rdata(input [31:0] dark_laplace_diff_0_update_0_read_rdata);

endmodule


module in_wire_dark_weights_update_0_read_dummy(output [31:0] dark_weights_update_0_read_dummy);

endmodule


module out_wire_dark_weights_update_0_read_rdata(input [31:0] dark_weights_update_0_read_rdata);

endmodule


module in_wire_dark_gauss_blur_2_update_0_write_wen(output [0:0] dark_gauss_blur_2_update_0_write_wen);

endmodule


module dark_gauss_ds_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_gauss_blur_2_update_0_write_wdata(output [31:0] dark_gauss_blur_2_update_0_write_wdata);

endmodule


module in_wire_dark_gauss_ds_2_update_0_read_dummy(output [31:0] dark_gauss_ds_2_update_0_read_dummy);

endmodule


module out_wire_dark_gauss_ds_2_update_0_read_rdata(input [31:0] dark_gauss_ds_2_update_0_read_rdata);

endmodule


module in_wire_dark_gauss_blur_3_update_0_write_wen(output [0:0] dark_gauss_blur_3_update_0_write_wen);

endmodule


module dark_gauss_blur_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] dark_gauss_ds_2_update_0_read_rdata, input [31:0] dark_gauss_blur_2_update_0_write_wdata, input [0:0] dark_gauss_blur_2_update_0_write_wen, input [31:0] dark_gauss_ds_2_update_0_read_dummy);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_gauss_ds_2_update_0_read_rdata
    // wr_3
  assign dark_gauss_ds_2_update_0_read_rdata = rd_2;

  // Bindings to dark_gauss_blur_2_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_gauss_blur_2_update_0_write_wdata;

  // Bindings to dark_gauss_blur_2_update_0_write_wen
    // rd_0
  assign rd_0 = dark_gauss_blur_2_update_0_write_wen;

  // selector_dark_gauss_ds_2_rd0_select
  logic [0:0] selector_dark_gauss_ds_2_rd0_select_clk;
  logic [0:0] selector_dark_gauss_ds_2_rd0_select_rst;
  logic [31:0] selector_dark_gauss_ds_2_rd0_select_d0;
  logic [31:0] selector_dark_gauss_ds_2_rd0_select_d1;
  logic [31:0] selector_dark_gauss_ds_2_rd0_select_out;
  dark_gauss_ds_2_rd0_select selector_dark_gauss_ds_2_rd0_select(.clk(selector_dark_gauss_ds_2_rd0_select_clk), .rst(selector_dark_gauss_ds_2_rd0_select_rst), .d0(selector_dark_gauss_ds_2_rd0_select_d0), .d1(selector_dark_gauss_ds_2_rd0_select_d1), .out(selector_dark_gauss_ds_2_rd0_select_out));
  assign selector_dark_gauss_ds_2_rd0_select_clk = clk;
  assign selector_dark_gauss_ds_2_rd0_select_rst = rst;
  // Bindings to selector_dark_gauss_ds_2_rd0_select

  // Bindings to dark_gauss_ds_2_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_gauss_ds_2_update_0_read_dummy;

  // dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1
  logic [0:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_done;
  dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1 dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1(.clk(dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_clk), .rst(dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_rst), .start(dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_start), .done(dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_done));
  assign dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_clk = clk;
  assign dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1



endmodule


module dark_gauss_ds_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_gauss_blur_3_update_0_write_wdata(output [31:0] dark_gauss_blur_3_update_0_write_wdata);

endmodule


module in_wire_dark_gauss_ds_3_update_0_read_dummy(output [31:0] dark_gauss_ds_3_update_0_read_dummy);

endmodule


module out_wire_dark_gauss_ds_3_update_0_read_rdata(input [31:0] dark_gauss_ds_3_update_0_read_rdata);

endmodule


module dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_52 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_52 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16



endmodule


module dark_gauss_ds_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [287:0] dark_gauss_blur_2_update_0_read_rdata, output [31:0] dark_laplace_us_0_update_0_read_rdata, input [31:0] dark_laplace_us_0_update_0_read_dummy, output [31:0] dark_laplace_diff_1_update_0_read_rdata, input [31:0] dark_laplace_diff_1_update_0_read_dummy, input [287:0] dark_gauss_blur_2_update_0_read_dummy, input [0:0] dark_gauss_ds_1_update_0_write_wen, input [31:0] dark_gauss_ds_1_update_0_write_wdata);

  logic [287:0] rd_2;
  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_4;
  logic [31:0] rd_6;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [287:0] rd_2_stage_1;
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_4_stage_1;
  reg [31:0] rd_6_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_2_stage_1 <= rd_2;
      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_4_stage_1 <= rd_4;
      rd_6_stage_1 <= rd_6;


    end

  end


  // Data processing units...
  // Bindings to dark_gauss_blur_2_update_0_read_rdata
    // wr_3
  assign dark_gauss_blur_2_update_0_read_rdata = rd_2;

  // selector_dark_gauss_blur_2_rd3_select
  logic [0:0] selector_dark_gauss_blur_2_rd3_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd3_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd3_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd3_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd3_select_out;
  dark_gauss_blur_2_rd3_select selector_dark_gauss_blur_2_rd3_select(.clk(selector_dark_gauss_blur_2_rd3_select_clk), .rst(selector_dark_gauss_blur_2_rd3_select_rst), .d0(selector_dark_gauss_blur_2_rd3_select_d0), .d1(selector_dark_gauss_blur_2_rd3_select_d1), .out(selector_dark_gauss_blur_2_rd3_select_out));
  assign selector_dark_gauss_blur_2_rd3_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd3_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd3_select

  // Bindings to dark_laplace_us_0_update_0_read_rdata
    // wr_7
  assign dark_laplace_us_0_update_0_read_rdata = rd_6;

  // Bindings to dark_laplace_us_0_update_0_read_dummy
    // rd_6
  assign rd_6 = dark_laplace_us_0_update_0_read_dummy;

  // Bindings to dark_laplace_diff_1_update_0_read_rdata
    // wr_5
  assign dark_laplace_diff_1_update_0_read_rdata = rd_4;

  // Bindings to dark_laplace_diff_1_update_0_read_dummy
    // rd_4
  assign rd_4 = dark_laplace_diff_1_update_0_read_dummy;

  // selector_dark_laplace_us_0_rd0_select
  logic [0:0] selector_dark_laplace_us_0_rd0_select_clk;
  logic [0:0] selector_dark_laplace_us_0_rd0_select_rst;
  logic [31:0] selector_dark_laplace_us_0_rd0_select_d0;
  logic [31:0] selector_dark_laplace_us_0_rd0_select_d1;
  logic [31:0] selector_dark_laplace_us_0_rd0_select_out;
  dark_laplace_us_0_rd0_select selector_dark_laplace_us_0_rd0_select(.clk(selector_dark_laplace_us_0_rd0_select_clk), .rst(selector_dark_laplace_us_0_rd0_select_rst), .d0(selector_dark_laplace_us_0_rd0_select_d0), .d1(selector_dark_laplace_us_0_rd0_select_d1), .out(selector_dark_laplace_us_0_rd0_select_out));
  assign selector_dark_laplace_us_0_rd0_select_clk = clk;
  assign selector_dark_laplace_us_0_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_us_0_rd0_select

  // selector_dark_laplace_diff_1_rd0_select
  logic [0:0] selector_dark_laplace_diff_1_rd0_select_clk;
  logic [0:0] selector_dark_laplace_diff_1_rd0_select_rst;
  logic [31:0] selector_dark_laplace_diff_1_rd0_select_d0;
  logic [31:0] selector_dark_laplace_diff_1_rd0_select_d1;
  logic [31:0] selector_dark_laplace_diff_1_rd0_select_out;
  dark_laplace_diff_1_rd0_select selector_dark_laplace_diff_1_rd0_select(.clk(selector_dark_laplace_diff_1_rd0_select_clk), .rst(selector_dark_laplace_diff_1_rd0_select_rst), .d0(selector_dark_laplace_diff_1_rd0_select_d0), .d1(selector_dark_laplace_diff_1_rd0_select_d1), .out(selector_dark_laplace_diff_1_rd0_select_out));
  assign selector_dark_laplace_diff_1_rd0_select_clk = clk;
  assign selector_dark_laplace_diff_1_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_diff_1_rd0_select

  // selector_dark_gauss_blur_2_rd8_select
  logic [0:0] selector_dark_gauss_blur_2_rd8_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd8_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd8_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd8_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd8_select_out;
  dark_gauss_blur_2_rd8_select selector_dark_gauss_blur_2_rd8_select(.clk(selector_dark_gauss_blur_2_rd8_select_clk), .rst(selector_dark_gauss_blur_2_rd8_select_rst), .d0(selector_dark_gauss_blur_2_rd8_select_d0), .d1(selector_dark_gauss_blur_2_rd8_select_d1), .out(selector_dark_gauss_blur_2_rd8_select_out));
  assign selector_dark_gauss_blur_2_rd8_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd8_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd8_select

  // selector_dark_gauss_blur_2_rd7_select
  logic [0:0] selector_dark_gauss_blur_2_rd7_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd7_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd7_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd7_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd7_select_out;
  dark_gauss_blur_2_rd7_select selector_dark_gauss_blur_2_rd7_select(.clk(selector_dark_gauss_blur_2_rd7_select_clk), .rst(selector_dark_gauss_blur_2_rd7_select_rst), .d0(selector_dark_gauss_blur_2_rd7_select_d0), .d1(selector_dark_gauss_blur_2_rd7_select_d1), .out(selector_dark_gauss_blur_2_rd7_select_out));
  assign selector_dark_gauss_blur_2_rd7_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd7_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd7_select

  // selector_dark_gauss_blur_2_rd4_select
  logic [0:0] selector_dark_gauss_blur_2_rd4_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd4_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd4_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd4_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd4_select_out;
  dark_gauss_blur_2_rd4_select selector_dark_gauss_blur_2_rd4_select(.clk(selector_dark_gauss_blur_2_rd4_select_clk), .rst(selector_dark_gauss_blur_2_rd4_select_rst), .d0(selector_dark_gauss_blur_2_rd4_select_d0), .d1(selector_dark_gauss_blur_2_rd4_select_d1), .out(selector_dark_gauss_blur_2_rd4_select_out));
  assign selector_dark_gauss_blur_2_rd4_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd4_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd4_select

  // selector_dark_gauss_blur_2_rd6_select
  logic [0:0] selector_dark_gauss_blur_2_rd6_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd6_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd6_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd6_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd6_select_out;
  dark_gauss_blur_2_rd6_select selector_dark_gauss_blur_2_rd6_select(.clk(selector_dark_gauss_blur_2_rd6_select_clk), .rst(selector_dark_gauss_blur_2_rd6_select_rst), .d0(selector_dark_gauss_blur_2_rd6_select_d0), .d1(selector_dark_gauss_blur_2_rd6_select_d1), .out(selector_dark_gauss_blur_2_rd6_select_out));
  assign selector_dark_gauss_blur_2_rd6_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd6_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd6_select

  // selector_dark_gauss_blur_2_rd5_select
  logic [0:0] selector_dark_gauss_blur_2_rd5_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd5_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd5_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd5_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd5_select_out;
  dark_gauss_blur_2_rd5_select selector_dark_gauss_blur_2_rd5_select(.clk(selector_dark_gauss_blur_2_rd5_select_clk), .rst(selector_dark_gauss_blur_2_rd5_select_rst), .d0(selector_dark_gauss_blur_2_rd5_select_d0), .d1(selector_dark_gauss_blur_2_rd5_select_d1), .out(selector_dark_gauss_blur_2_rd5_select_out));
  assign selector_dark_gauss_blur_2_rd5_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd5_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd5_select

  // selector_dark_gauss_blur_2_rd2_select
  logic [0:0] selector_dark_gauss_blur_2_rd2_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd2_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd2_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd2_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd2_select_out;
  dark_gauss_blur_2_rd2_select selector_dark_gauss_blur_2_rd2_select(.clk(selector_dark_gauss_blur_2_rd2_select_clk), .rst(selector_dark_gauss_blur_2_rd2_select_rst), .d0(selector_dark_gauss_blur_2_rd2_select_d0), .d1(selector_dark_gauss_blur_2_rd2_select_d1), .out(selector_dark_gauss_blur_2_rd2_select_out));
  assign selector_dark_gauss_blur_2_rd2_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd2_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd2_select

  // Bindings to dark_gauss_blur_2_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_gauss_blur_2_update_0_read_dummy;

  // selector_dark_gauss_blur_2_rd0_select
  logic [0:0] selector_dark_gauss_blur_2_rd0_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd0_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd0_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd0_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd0_select_out;
  dark_gauss_blur_2_rd0_select selector_dark_gauss_blur_2_rd0_select(.clk(selector_dark_gauss_blur_2_rd0_select_clk), .rst(selector_dark_gauss_blur_2_rd0_select_rst), .d0(selector_dark_gauss_blur_2_rd0_select_d0), .d1(selector_dark_gauss_blur_2_rd0_select_d1), .out(selector_dark_gauss_blur_2_rd0_select_out));
  assign selector_dark_gauss_blur_2_rd0_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd0_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd0_select

  // dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_clk;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_rst;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_start;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_done;
  dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0 dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0(.clk(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_clk), .rst(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_rst), .start(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_start), .done(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_done));
  assign dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_clk = clk;
  assign dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_rst = rst;
  // Bindings to dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0

  // Bindings to dark_gauss_ds_1_update_0_write_wen
    // rd_0
  assign rd_0 = dark_gauss_ds_1_update_0_write_wen;

  // selector_dark_gauss_blur_2_rd1_select
  logic [0:0] selector_dark_gauss_blur_2_rd1_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd1_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd1_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd1_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd1_select_out;
  dark_gauss_blur_2_rd1_select selector_dark_gauss_blur_2_rd1_select(.clk(selector_dark_gauss_blur_2_rd1_select_clk), .rst(selector_dark_gauss_blur_2_rd1_select_rst), .d0(selector_dark_gauss_blur_2_rd1_select_d0), .d1(selector_dark_gauss_blur_2_rd1_select_d1), .out(selector_dark_gauss_blur_2_rd1_select_out));
  assign selector_dark_gauss_blur_2_rd1_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd1_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd1_select

  // Bindings to dark_gauss_ds_1_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_gauss_ds_1_update_0_write_wdata;

  // dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9_clk;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9_rst;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9_start;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9_done;
  dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9 dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9(.clk(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9_clk), .rst(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9_rst), .start(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9_start), .done(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9_done));
  assign dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9_clk = clk;
  assign dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9_rst = rst;
  // Bindings to dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_9

  // dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0_clk;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0_rst;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0_start;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0_done;
  dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0 dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0(.clk(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0_clk), .rst(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0_rst), .start(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0_start), .done(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0_done));
  assign dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0_clk = clk;
  assign dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0_rst = rst;
  // Bindings to dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0



endmodule


module dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_diff_1_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_279 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114



endmodule


module in_wire_dark_gauss_ds_3_update_0_write_wen(output [0:0] dark_gauss_ds_3_update_0_write_wen);

endmodule


module in_wire_dark_gauss_ds_3_update_0_write_wdata(output [31:0] dark_gauss_ds_3_update_0_write_wdata);

endmodule


module dark_laplace_us_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = ((-1 - d1) % 2 == 0 && 23 - d0 >= 0) ? ((12 - floord(2*d0, 4))) : 0;
    end
  end

endmodule


module in_wire_dark_laplace_us_2_update_0_read_dummy(output [31:0] dark_laplace_us_2_update_0_read_dummy);

endmodule


module out_wire_dark_laplace_us_2_update_0_read_rdata(input [31:0] dark_laplace_us_2_update_0_read_rdata);

endmodule


module dark_gauss_ds_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_gauss_ds_3_update_0_write_wen, input [31:0] dark_gauss_ds_3_update_0_write_wdata, input [31:0] dark_laplace_us_2_update_0_read_dummy, output [31:0] dark_laplace_us_2_update_0_read_rdata, input [31:0] fused_level_3_update_0_read_dummy, output [31:0] fused_level_3_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_clk;
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_rst;
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_start;
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_done;
  dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0 dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0(.clk(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_clk), .rst(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_rst), .start(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_start), .done(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_done));
  assign dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_clk = clk;
  assign dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_rst = rst;
  // Bindings to dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0

  // dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_done;
  dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1 dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1(.clk(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_clk), .rst(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_rst), .start(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_start), .done(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_done));
  assign dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_clk = clk;
  assign dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1

  // Bindings to dark_gauss_ds_3_update_0_write_wen
    // rd_0
  assign rd_0 = dark_gauss_ds_3_update_0_write_wen;

  // Bindings to dark_gauss_ds_3_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_gauss_ds_3_update_0_write_wdata;

  // selector_dark_laplace_us_2_rd0_select
  logic [0:0] selector_dark_laplace_us_2_rd0_select_clk;
  logic [0:0] selector_dark_laplace_us_2_rd0_select_rst;
  logic [31:0] selector_dark_laplace_us_2_rd0_select_d0;
  logic [31:0] selector_dark_laplace_us_2_rd0_select_d1;
  logic [31:0] selector_dark_laplace_us_2_rd0_select_out;
  dark_laplace_us_2_rd0_select selector_dark_laplace_us_2_rd0_select(.clk(selector_dark_laplace_us_2_rd0_select_clk), .rst(selector_dark_laplace_us_2_rd0_select_rst), .d0(selector_dark_laplace_us_2_rd0_select_d0), .d1(selector_dark_laplace_us_2_rd0_select_d1), .out(selector_dark_laplace_us_2_rd0_select_out));
  assign selector_dark_laplace_us_2_rd0_select_clk = clk;
  assign selector_dark_laplace_us_2_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_us_2_rd0_select

  // selector_fused_level_3_rd0_select
  logic [0:0] selector_fused_level_3_rd0_select_clk;
  logic [0:0] selector_fused_level_3_rd0_select_rst;
  logic [31:0] selector_fused_level_3_rd0_select_d0;
  logic [31:0] selector_fused_level_3_rd0_select_d1;
  logic [31:0] selector_fused_level_3_rd0_select_out;
  fused_level_3_rd0_select selector_fused_level_3_rd0_select(.clk(selector_fused_level_3_rd0_select_clk), .rst(selector_fused_level_3_rd0_select_rst), .d0(selector_fused_level_3_rd0_select_d0), .d1(selector_fused_level_3_rd0_select_d1), .out(selector_fused_level_3_rd0_select_out));
  assign selector_fused_level_3_rd0_select_clk = clk;
  assign selector_fused_level_3_rd0_select_rst = rst;
  // Bindings to selector_fused_level_3_rd0_select

  // Bindings to dark_laplace_us_2_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_laplace_us_2_update_0_read_dummy;

  // Bindings to dark_laplace_us_2_update_0_read_rdata
    // wr_3
  assign dark_laplace_us_2_update_0_read_rdata = rd_2;

  // Bindings to fused_level_3_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_3_update_0_read_dummy;

  // Bindings to fused_level_3_update_0_read_rdata
    // wr_5
  assign fused_level_3_update_0_read_rdata = rd_4;



endmodule


module dark_weights_normed(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] fused_level_0_update_0_read_dummy, input [0:0] dark_weights_normed_update_0_write_wen, input [31:0] dark_weights_normed_update_0_write_wdata, input [287:0] dark_weights_normed_gauss_blur_1_update_0_read_dummy, output [287:0] dark_weights_normed_gauss_blur_1_update_0_read_rdata, output [31:0] fused_level_0_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_clk;
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_rst;
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_start;
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_done;
  dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0 dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0(.clk(dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_clk), .rst(dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_rst), .start(dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_start), .done(dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_done));
  assign dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_clk = clk;
  assign dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_rst = rst;
  // Bindings to dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0

  // Bindings to fused_level_0_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_0_update_0_read_dummy;

  // selector_dark_weights_normed_gauss_blur_1_rd1_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd1_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd1_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd1_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd1_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd1_select_out;
  dark_weights_normed_gauss_blur_1_rd1_select selector_dark_weights_normed_gauss_blur_1_rd1_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd1_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd1_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd1_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd1_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd1_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd1_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd1_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd1_select

  // selector_dark_weights_normed_gauss_blur_1_rd0_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd0_select_out;
  dark_weights_normed_gauss_blur_1_rd0_select selector_dark_weights_normed_gauss_blur_1_rd0_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd0_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd0_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd0_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd0_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd0_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd0_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd0_select

  // selector_fused_level_0_rd0_select
  logic [0:0] selector_fused_level_0_rd0_select_clk;
  logic [0:0] selector_fused_level_0_rd0_select_rst;
  logic [31:0] selector_fused_level_0_rd0_select_d0;
  logic [31:0] selector_fused_level_0_rd0_select_d1;
  logic [31:0] selector_fused_level_0_rd0_select_out;
  fused_level_0_rd0_select selector_fused_level_0_rd0_select(.clk(selector_fused_level_0_rd0_select_clk), .rst(selector_fused_level_0_rd0_select_rst), .d0(selector_fused_level_0_rd0_select_d0), .d1(selector_fused_level_0_rd0_select_d1), .out(selector_fused_level_0_rd0_select_out));
  assign selector_fused_level_0_rd0_select_clk = clk;
  assign selector_fused_level_0_rd0_select_rst = rst;
  // Bindings to selector_fused_level_0_rd0_select

  // selector_dark_weights_normed_gauss_blur_1_rd2_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd2_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd2_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd2_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd2_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd2_select_out;
  dark_weights_normed_gauss_blur_1_rd2_select selector_dark_weights_normed_gauss_blur_1_rd2_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd2_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd2_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd2_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd2_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd2_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd2_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd2_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd2_select

  // selector_dark_weights_normed_gauss_blur_1_rd3_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd3_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd3_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd3_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd3_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd3_select_out;
  dark_weights_normed_gauss_blur_1_rd3_select selector_dark_weights_normed_gauss_blur_1_rd3_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd3_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd3_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd3_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd3_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd3_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd3_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd3_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd3_select

  // selector_dark_weights_normed_gauss_blur_1_rd4_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd4_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd4_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd4_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd4_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd4_select_out;
  dark_weights_normed_gauss_blur_1_rd4_select selector_dark_weights_normed_gauss_blur_1_rd4_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd4_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd4_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd4_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd4_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd4_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd4_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd4_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd4_select

  // selector_dark_weights_normed_gauss_blur_1_rd6_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd6_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd6_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd6_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd6_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd6_select_out;
  dark_weights_normed_gauss_blur_1_rd6_select selector_dark_weights_normed_gauss_blur_1_rd6_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd6_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd6_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd6_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd6_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd6_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd6_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd6_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd6_select

  // selector_dark_weights_normed_gauss_blur_1_rd5_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd5_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd5_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd5_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd5_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd5_select_out;
  dark_weights_normed_gauss_blur_1_rd5_select selector_dark_weights_normed_gauss_blur_1_rd5_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd5_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd5_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd5_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd5_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd5_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd5_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd5_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd5_select

  // Bindings to dark_weights_normed_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_normed_update_0_write_wen;

  // selector_dark_weights_normed_gauss_blur_1_rd7_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd7_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd7_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd7_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd7_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd7_select_out;
  dark_weights_normed_gauss_blur_1_rd7_select selector_dark_weights_normed_gauss_blur_1_rd7_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd7_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd7_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd7_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd7_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd7_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd7_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd7_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd7_select

  // selector_dark_weights_normed_gauss_blur_1_rd8_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd8_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd8_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd8_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd8_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd8_select_out;
  dark_weights_normed_gauss_blur_1_rd8_select selector_dark_weights_normed_gauss_blur_1_rd8_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd8_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd8_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd8_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd8_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd8_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd8_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd8_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd8_select

  // Bindings to dark_weights_normed_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_normed_update_0_write_wdata;

  // Bindings to dark_weights_normed_gauss_blur_1_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_weights_normed_gauss_blur_1_update_0_read_dummy;

  // Bindings to dark_weights_normed_gauss_blur_1_update_0_read_rdata
    // wr_3
  assign dark_weights_normed_gauss_blur_1_update_0_read_rdata = rd_2;

  // Bindings to fused_level_0_update_0_read_rdata
    // wr_5
  assign fused_level_0_update_0_read_rdata = rd_4;

  // dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_clk;
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_rst;
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_start;
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_done;
  dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9 dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9(.clk(dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_clk), .rst(dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_rst), .start(dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_start), .done(dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_done));
  assign dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_clk = clk;
  assign dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_rst = rst;
  // Bindings to dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9



endmodule


module in_wire_dark_laplace_diff_1_update_0_write_wen(output [0:0] dark_laplace_diff_1_update_0_write_wen);

endmodule


module in_wire_dark_laplace_diff_1_update_0_write_wdata(output [31:0] dark_laplace_diff_1_update_0_write_wdata);

endmodule


module dark_weights_normed_gauss_blur_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] dark_weights_normed_gauss_blur_1_update_0_write_wdata, input [31:0] dark_weights_normed_gauss_ds_1_update_0_read_dummy, input [0:0] dark_weights_normed_gauss_blur_1_update_0_write_wen, output [31:0] dark_weights_normed_gauss_ds_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_weights_normed_gauss_blur_1_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_normed_gauss_blur_1_update_0_write_wdata;

  // Bindings to dark_weights_normed_gauss_ds_1_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_weights_normed_gauss_ds_1_update_0_read_dummy;

  // selector_dark_weights_normed_gauss_ds_1_rd0_select
  logic [0:0] selector_dark_weights_normed_gauss_ds_1_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_ds_1_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_ds_1_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_ds_1_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_ds_1_rd0_select_out;
  dark_weights_normed_gauss_ds_1_rd0_select selector_dark_weights_normed_gauss_ds_1_rd0_select(.clk(selector_dark_weights_normed_gauss_ds_1_rd0_select_clk), .rst(selector_dark_weights_normed_gauss_ds_1_rd0_select_rst), .d0(selector_dark_weights_normed_gauss_ds_1_rd0_select_d0), .d1(selector_dark_weights_normed_gauss_ds_1_rd0_select_d1), .out(selector_dark_weights_normed_gauss_ds_1_rd0_select_out));
  assign selector_dark_weights_normed_gauss_ds_1_rd0_select_clk = clk;
  assign selector_dark_weights_normed_gauss_ds_1_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_ds_1_rd0_select

  // dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1
  logic [0:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_done;
  dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1 dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1(.clk(dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_clk), .rst(dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_rst), .start(dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_start), .done(dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_done));
  assign dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_clk = clk;
  assign dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1

  // Bindings to dark_weights_normed_gauss_blur_1_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_normed_gauss_blur_1_update_0_write_wen;

  // Bindings to dark_weights_normed_gauss_ds_1_update_0_read_rdata
    // wr_3
  assign dark_weights_normed_gauss_ds_1_update_0_read_rdata = rd_2;



endmodule


module in_wire_dark_weights_normed_gauss_blur_3_update_0_write_wen(output [0:0] dark_weights_normed_gauss_blur_3_update_0_write_wen);

endmodule


module dark_weights_normed_gauss_ds_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_gauss_blur_3_update_0_write_wdata(output [31:0] dark_weights_normed_gauss_blur_3_update_0_write_wdata);

endmodule


module dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_weights_normed_gauss_ds_3_update_0_read_dummy(output [31:0] dark_weights_normed_gauss_ds_3_update_0_read_dummy);

endmodule


module out_wire_dark_weights_normed_gauss_ds_3_update_0_read_rdata(input [31:0] dark_weights_normed_gauss_ds_3_update_0_read_rdata);

endmodule


module in_wire_dark_weights_normed_gauss_ds_3_update_0_write_wen(output [0:0] dark_weights_normed_gauss_ds_3_update_0_write_wen);

endmodule


module fused_level_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_gauss_ds_3_update_0_write_wdata(output [31:0] dark_weights_normed_gauss_ds_3_update_0_write_wdata);

endmodule


module dark_weights_normed_gauss_ds_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] fused_level_3_update_0_read_dummy, input [0:0] dark_weights_normed_gauss_ds_3_update_0_write_wen, input [31:0] dark_weights_normed_gauss_ds_3_update_0_write_wdata, output [31:0] fused_level_3_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1
  logic [0:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_done;
  dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1 dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1(.clk(dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_clk), .rst(dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_rst), .start(dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_start), .done(dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_done));
  assign dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_clk = clk;
  assign dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1

  // Bindings to fused_level_3_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_3_update_0_read_dummy;

  // Bindings to dark_weights_normed_gauss_ds_3_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_normed_gauss_ds_3_update_0_write_wen;

  // selector_fused_level_3_rd0_select
  logic [0:0] selector_fused_level_3_rd0_select_clk;
  logic [0:0] selector_fused_level_3_rd0_select_rst;
  logic [31:0] selector_fused_level_3_rd0_select_d0;
  logic [31:0] selector_fused_level_3_rd0_select_d1;
  logic [31:0] selector_fused_level_3_rd0_select_out;
  fused_level_3_rd0_select selector_fused_level_3_rd0_select(.clk(selector_fused_level_3_rd0_select_clk), .rst(selector_fused_level_3_rd0_select_rst), .d0(selector_fused_level_3_rd0_select_d0), .d1(selector_fused_level_3_rd0_select_d1), .out(selector_fused_level_3_rd0_select_out));
  assign selector_fused_level_3_rd0_select_clk = clk;
  assign selector_fused_level_3_rd0_select_rst = rst;
  // Bindings to selector_fused_level_3_rd0_select

  // Bindings to dark_weights_normed_gauss_ds_3_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_normed_gauss_ds_3_update_0_write_wdata;

  // Bindings to fused_level_3_update_0_read_rdata
    // wr_3
  assign fused_level_3_update_0_read_rdata = rd_2;



endmodule


module final_merged_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] final_merged_0_update_0_write_wen, input [31:0] final_merged_0_update_0_write_wdata, input [31:0] pyramid_synthetic_exposure_fusion_update_0_read_dummy, output [31:0] pyramid_synthetic_exposure_fusion_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // final_merged_0_final_merged_0_update_0_write0_merged_banks_1
  logic [0:0] final_merged_0_final_merged_0_update_0_write0_merged_banks_1_clk;
  logic [0:0] final_merged_0_final_merged_0_update_0_write0_merged_banks_1_rst;
  logic [0:0] final_merged_0_final_merged_0_update_0_write0_merged_banks_1_start;
  logic [0:0] final_merged_0_final_merged_0_update_0_write0_merged_banks_1_done;
  final_merged_0_final_merged_0_update_0_write0_merged_banks_1 final_merged_0_final_merged_0_update_0_write0_merged_banks_1(.clk(final_merged_0_final_merged_0_update_0_write0_merged_banks_1_clk), .rst(final_merged_0_final_merged_0_update_0_write0_merged_banks_1_rst), .start(final_merged_0_final_merged_0_update_0_write0_merged_banks_1_start), .done(final_merged_0_final_merged_0_update_0_write0_merged_banks_1_done));
  assign final_merged_0_final_merged_0_update_0_write0_merged_banks_1_clk = clk;
  assign final_merged_0_final_merged_0_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to final_merged_0_final_merged_0_update_0_write0_merged_banks_1

  // Bindings to final_merged_0_update_0_write_wen
    // rd_0
  assign rd_0 = final_merged_0_update_0_write_wen;

  // selector_pyramid_synthetic_exposure_fusion_rd0_select
  logic [0:0] selector_pyramid_synthetic_exposure_fusion_rd0_select_clk;
  logic [0:0] selector_pyramid_synthetic_exposure_fusion_rd0_select_rst;
  logic [31:0] selector_pyramid_synthetic_exposure_fusion_rd0_select_d0;
  logic [31:0] selector_pyramid_synthetic_exposure_fusion_rd0_select_d1;
  logic [31:0] selector_pyramid_synthetic_exposure_fusion_rd0_select_out;
  pyramid_synthetic_exposure_fusion_rd0_select selector_pyramid_synthetic_exposure_fusion_rd0_select(.clk(selector_pyramid_synthetic_exposure_fusion_rd0_select_clk), .rst(selector_pyramid_synthetic_exposure_fusion_rd0_select_rst), .d0(selector_pyramid_synthetic_exposure_fusion_rd0_select_d0), .d1(selector_pyramid_synthetic_exposure_fusion_rd0_select_d1), .out(selector_pyramid_synthetic_exposure_fusion_rd0_select_out));
  assign selector_pyramid_synthetic_exposure_fusion_rd0_select_clk = clk;
  assign selector_pyramid_synthetic_exposure_fusion_rd0_select_rst = rst;
  // Bindings to selector_pyramid_synthetic_exposure_fusion_rd0_select

  // Bindings to final_merged_0_update_0_write_wdata
    // rd_1
  assign rd_1 = final_merged_0_update_0_write_wdata;

  // Bindings to pyramid_synthetic_exposure_fusion_update_0_read_dummy
    // rd_2
  assign rd_2 = pyramid_synthetic_exposure_fusion_update_0_read_dummy;

  // Bindings to pyramid_synthetic_exposure_fusion_update_0_read_rdata
    // wr_3
  assign pyramid_synthetic_exposure_fusion_update_0_read_rdata = rd_2;



endmodule


module fused_level_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] fused_level_0_update_0_write_wen, input [31:0] fused_level_0_update_0_write_wdata, input [31:0] final_merged_0_update_0_read_dummy, output [31:0] final_merged_0_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to fused_level_0_update_0_write_wen
    // rd_0
  assign rd_0 = fused_level_0_update_0_write_wen;

  // fused_level_0_fused_level_0_update_0_write0_merged_banks_1
  logic [0:0] fused_level_0_fused_level_0_update_0_write0_merged_banks_1_clk;
  logic [0:0] fused_level_0_fused_level_0_update_0_write0_merged_banks_1_rst;
  logic [0:0] fused_level_0_fused_level_0_update_0_write0_merged_banks_1_start;
  logic [0:0] fused_level_0_fused_level_0_update_0_write0_merged_banks_1_done;
  fused_level_0_fused_level_0_update_0_write0_merged_banks_1 fused_level_0_fused_level_0_update_0_write0_merged_banks_1(.clk(fused_level_0_fused_level_0_update_0_write0_merged_banks_1_clk), .rst(fused_level_0_fused_level_0_update_0_write0_merged_banks_1_rst), .start(fused_level_0_fused_level_0_update_0_write0_merged_banks_1_start), .done(fused_level_0_fused_level_0_update_0_write0_merged_banks_1_done));
  assign fused_level_0_fused_level_0_update_0_write0_merged_banks_1_clk = clk;
  assign fused_level_0_fused_level_0_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to fused_level_0_fused_level_0_update_0_write0_merged_banks_1

  // selector_final_merged_0_rd0_select
  logic [0:0] selector_final_merged_0_rd0_select_clk;
  logic [0:0] selector_final_merged_0_rd0_select_rst;
  logic [31:0] selector_final_merged_0_rd0_select_d0;
  logic [31:0] selector_final_merged_0_rd0_select_d1;
  logic [31:0] selector_final_merged_0_rd0_select_out;
  final_merged_0_rd0_select selector_final_merged_0_rd0_select(.clk(selector_final_merged_0_rd0_select_clk), .rst(selector_final_merged_0_rd0_select_rst), .d0(selector_final_merged_0_rd0_select_d0), .d1(selector_final_merged_0_rd0_select_d1), .out(selector_final_merged_0_rd0_select_out));
  assign selector_final_merged_0_rd0_select_clk = clk;
  assign selector_final_merged_0_rd0_select_rst = rst;
  // Bindings to selector_final_merged_0_rd0_select

  // Bindings to fused_level_0_update_0_write_wdata
    // rd_1
  assign rd_1 = fused_level_0_update_0_write_wdata;

  // Bindings to final_merged_0_update_0_read_dummy
    // rd_2
  assign rd_2 = final_merged_0_update_0_read_dummy;

  // Bindings to final_merged_0_update_0_read_rdata
    // wr_3
  assign final_merged_0_update_0_read_rdata = rd_2;



endmodule


module fused_level_1_fused_level_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module fused_level_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] fused_level_1_update_0_write_wen, input [31:0] fused_level_1_update_0_write_wdata, input [31:0] final_merged_1_update_0_read_dummy, output [31:0] final_merged_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to fused_level_1_update_0_write_wen
    // rd_0
  assign rd_0 = fused_level_1_update_0_write_wen;

  // fused_level_1_fused_level_1_update_0_write0_merged_banks_1
  logic [0:0] fused_level_1_fused_level_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] fused_level_1_fused_level_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] fused_level_1_fused_level_1_update_0_write0_merged_banks_1_start;
  logic [0:0] fused_level_1_fused_level_1_update_0_write0_merged_banks_1_done;
  fused_level_1_fused_level_1_update_0_write0_merged_banks_1 fused_level_1_fused_level_1_update_0_write0_merged_banks_1(.clk(fused_level_1_fused_level_1_update_0_write0_merged_banks_1_clk), .rst(fused_level_1_fused_level_1_update_0_write0_merged_banks_1_rst), .start(fused_level_1_fused_level_1_update_0_write0_merged_banks_1_start), .done(fused_level_1_fused_level_1_update_0_write0_merged_banks_1_done));
  assign fused_level_1_fused_level_1_update_0_write0_merged_banks_1_clk = clk;
  assign fused_level_1_fused_level_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to fused_level_1_fused_level_1_update_0_write0_merged_banks_1

  // selector_final_merged_1_rd0_select
  logic [0:0] selector_final_merged_1_rd0_select_clk;
  logic [0:0] selector_final_merged_1_rd0_select_rst;
  logic [31:0] selector_final_merged_1_rd0_select_d0;
  logic [31:0] selector_final_merged_1_rd0_select_d1;
  logic [31:0] selector_final_merged_1_rd0_select_out;
  final_merged_1_rd0_select selector_final_merged_1_rd0_select(.clk(selector_final_merged_1_rd0_select_clk), .rst(selector_final_merged_1_rd0_select_rst), .d0(selector_final_merged_1_rd0_select_d0), .d1(selector_final_merged_1_rd0_select_d1), .out(selector_final_merged_1_rd0_select_out));
  assign selector_final_merged_1_rd0_select_clk = clk;
  assign selector_final_merged_1_rd0_select_rst = rst;
  // Bindings to selector_final_merged_1_rd0_select

  // Bindings to fused_level_1_update_0_write_wdata
    // rd_1
  assign rd_1 = fused_level_1_update_0_write_wdata;

  // Bindings to final_merged_1_update_0_read_dummy
    // rd_2
  assign rd_2 = final_merged_1_update_0_read_dummy;

  // Bindings to final_merged_1_update_0_read_rdata
    // wr_3
  assign final_merged_1_update_0_read_rdata = rd_2;



endmodule


module fused_level_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] fused_level_2_update_0_write_wen, input [31:0] fused_level_2_update_0_write_wdata, input [31:0] final_merged_2_update_0_read_dummy, output [31:0] final_merged_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // selector_final_merged_2_rd0_select
  logic [0:0] selector_final_merged_2_rd0_select_clk;
  logic [0:0] selector_final_merged_2_rd0_select_rst;
  logic [31:0] selector_final_merged_2_rd0_select_d0;
  logic [31:0] selector_final_merged_2_rd0_select_d1;
  logic [31:0] selector_final_merged_2_rd0_select_out;
  final_merged_2_rd0_select selector_final_merged_2_rd0_select(.clk(selector_final_merged_2_rd0_select_clk), .rst(selector_final_merged_2_rd0_select_rst), .d0(selector_final_merged_2_rd0_select_d0), .d1(selector_final_merged_2_rd0_select_d1), .out(selector_final_merged_2_rd0_select_out));
  assign selector_final_merged_2_rd0_select_clk = clk;
  assign selector_final_merged_2_rd0_select_rst = rst;
  // Bindings to selector_final_merged_2_rd0_select

  // fused_level_2_fused_level_2_update_0_write0_merged_banks_1
  logic [0:0] fused_level_2_fused_level_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] fused_level_2_fused_level_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] fused_level_2_fused_level_2_update_0_write0_merged_banks_1_start;
  logic [0:0] fused_level_2_fused_level_2_update_0_write0_merged_banks_1_done;
  fused_level_2_fused_level_2_update_0_write0_merged_banks_1 fused_level_2_fused_level_2_update_0_write0_merged_banks_1(.clk(fused_level_2_fused_level_2_update_0_write0_merged_banks_1_clk), .rst(fused_level_2_fused_level_2_update_0_write0_merged_banks_1_rst), .start(fused_level_2_fused_level_2_update_0_write0_merged_banks_1_start), .done(fused_level_2_fused_level_2_update_0_write0_merged_banks_1_done));
  assign fused_level_2_fused_level_2_update_0_write0_merged_banks_1_clk = clk;
  assign fused_level_2_fused_level_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to fused_level_2_fused_level_2_update_0_write0_merged_banks_1

  // Bindings to fused_level_2_update_0_write_wen
    // rd_0
  assign rd_0 = fused_level_2_update_0_write_wen;

  // Bindings to fused_level_2_update_0_write_wdata
    // rd_1
  assign rd_1 = fused_level_2_update_0_write_wdata;

  // Bindings to final_merged_2_update_0_read_dummy
    // rd_2
  assign rd_2 = final_merged_2_update_0_read_dummy;

  // Bindings to final_merged_2_update_0_read_rdata
    // wr_3
  assign final_merged_2_update_0_read_rdata = rd_2;



endmodule


module in_wire_in_update_0_write_wen(output [0:0] in_update_0_write_wen);

endmodule


module bright_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_in_update_0_write_wdata(output [31:0] in_update_0_write_wdata);

endmodule


module in_wire_bright_update_0_read_dummy(output [31:0] bright_update_0_read_dummy);

endmodule


module out_wire_bright_update_0_read_rdata(input [31:0] bright_update_0_read_rdata);

endmodule


module in_wire_dark_update_0_read_dummy(output [31:0] dark_update_0_read_dummy);

endmodule


module out_wire_dark_update_0_read_rdata(input [31:0] dark_update_0_read_rdata);

endmodule


module in(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] in_update_0_write_wen, input [31:0] in_update_0_write_wdata, input [31:0] bright_update_0_read_dummy, output [31:0] bright_update_0_read_rdata, input [31:0] dark_update_0_read_dummy, output [31:0] dark_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // selector_bright_rd0_select
  logic [0:0] selector_bright_rd0_select_clk;
  logic [0:0] selector_bright_rd0_select_rst;
  logic [31:0] selector_bright_rd0_select_d0;
  logic [31:0] selector_bright_rd0_select_d1;
  logic [31:0] selector_bright_rd0_select_out;
  bright_rd0_select selector_bright_rd0_select(.clk(selector_bright_rd0_select_clk), .rst(selector_bright_rd0_select_rst), .d0(selector_bright_rd0_select_d0), .d1(selector_bright_rd0_select_d1), .out(selector_bright_rd0_select_out));
  assign selector_bright_rd0_select_clk = clk;
  assign selector_bright_rd0_select_rst = rst;
  // Bindings to selector_bright_rd0_select

  // selector_dark_rd0_select
  logic [0:0] selector_dark_rd0_select_clk;
  logic [0:0] selector_dark_rd0_select_rst;
  logic [31:0] selector_dark_rd0_select_d0;
  logic [31:0] selector_dark_rd0_select_d1;
  logic [31:0] selector_dark_rd0_select_out;
  dark_rd0_select selector_dark_rd0_select(.clk(selector_dark_rd0_select_clk), .rst(selector_dark_rd0_select_rst), .d0(selector_dark_rd0_select_d0), .d1(selector_dark_rd0_select_d1), .out(selector_dark_rd0_select_out));
  assign selector_dark_rd0_select_clk = clk;
  assign selector_dark_rd0_select_rst = rst;
  // Bindings to selector_dark_rd0_select

  // Bindings to in_update_0_write_wen
    // rd_0
  assign rd_0 = in_update_0_write_wen;

  // Bindings to in_update_0_write_wdata
    // rd_1
  assign rd_1 = in_update_0_write_wdata;

  // Bindings to bright_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_update_0_read_dummy;

  // Bindings to bright_update_0_read_rdata
    // wr_3
  assign bright_update_0_read_rdata = rd_2;

  // Bindings to dark_update_0_read_dummy
    // rd_4
  assign rd_4 = dark_update_0_read_dummy;

  // Bindings to dark_update_0_read_rdata
    // wr_5
  assign dark_update_0_read_rdata = rd_4;

  // in_in_update_0_write0_merged_banks_2
  logic [0:0] in_in_update_0_write0_merged_banks_2_clk;
  logic [0:0] in_in_update_0_write0_merged_banks_2_rst;
  logic [0:0] in_in_update_0_write0_merged_banks_2_start;
  logic [0:0] in_in_update_0_write0_merged_banks_2_done;
  in_in_update_0_write0_merged_banks_2 in_in_update_0_write0_merged_banks_2(.clk(in_in_update_0_write0_merged_banks_2_clk), .rst(in_in_update_0_write0_merged_banks_2_rst), .start(in_in_update_0_write0_merged_banks_2_start), .done(in_in_update_0_write0_merged_banks_2_done));
  assign in_in_update_0_write0_merged_banks_2_clk = clk;
  assign in_in_update_0_write0_merged_banks_2_rst = rst;
  // Bindings to in_in_update_0_write0_merged_banks_2



endmodule


module in_wire_in_off_chip_update_0_write_wen(output [0:0] in_off_chip_update_0_write_wen);

endmodule


module in_wire_in_off_chip_update_0_write_wdata(output [31:0] in_off_chip_update_0_write_wdata);

endmodule


module in_wire_in_update_0_read_dummy(output [31:0] in_update_0_read_dummy);

endmodule


module out_wire_in_update_0_read_rdata(input [31:0] in_update_0_read_rdata);

endmodule


module in_wire_pyramid_synthetic_exposure_fusion_update_0_write_wen(output [0:0] pyramid_synthetic_exposure_fusion_update_0_write_wen);

endmodule


module in_wire_pyramid_synthetic_exposure_fusion_update_0_write_wdata(output [31:0] pyramid_synthetic_exposure_fusion_update_0_write_wdata);

endmodule


module pyramid_synthetic_exposure_fusion(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] pyramid_synthetic_exposure_fusion_update_0_write_wen, input [31:0] pyramid_synthetic_exposure_fusion_update_0_write_wdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;


    end

  end


  // Data processing units...
  // Bindings to pyramid_synthetic_exposure_fusion_update_0_write_wen
    // rd_0
  assign rd_0 = pyramid_synthetic_exposure_fusion_update_0_write_wen;

  // Bindings to pyramid_synthetic_exposure_fusion_update_0_write_wdata
    // rd_1
  assign rd_1 = pyramid_synthetic_exposure_fusion_update_0_write_wdata;



endmodule


module weight_sums_weight_sums_update_0_write0_merged_banks_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_weight_sums_update_0_write_wen(output [0:0] weight_sums_update_0_write_wen);

endmodule


module bright_weights_normed_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_weights_normed_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_weight_sums_update_0_write_wdata(output [31:0] weight_sums_update_0_write_wdata);

endmodule


module weight_sums(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] weight_sums_update_0_write_wen, input [31:0] weight_sums_update_0_write_wdata, input [31:0] bright_weights_normed_update_0_read_dummy, output [31:0] bright_weights_normed_update_0_read_rdata, input [31:0] dark_weights_normed_update_0_read_dummy, output [31:0] dark_weights_normed_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // weight_sums_weight_sums_update_0_write0_merged_banks_2
  logic [0:0] weight_sums_weight_sums_update_0_write0_merged_banks_2_clk;
  logic [0:0] weight_sums_weight_sums_update_0_write0_merged_banks_2_rst;
  logic [0:0] weight_sums_weight_sums_update_0_write0_merged_banks_2_start;
  logic [0:0] weight_sums_weight_sums_update_0_write0_merged_banks_2_done;
  weight_sums_weight_sums_update_0_write0_merged_banks_2 weight_sums_weight_sums_update_0_write0_merged_banks_2(.clk(weight_sums_weight_sums_update_0_write0_merged_banks_2_clk), .rst(weight_sums_weight_sums_update_0_write0_merged_banks_2_rst), .start(weight_sums_weight_sums_update_0_write0_merged_banks_2_start), .done(weight_sums_weight_sums_update_0_write0_merged_banks_2_done));
  assign weight_sums_weight_sums_update_0_write0_merged_banks_2_clk = clk;
  assign weight_sums_weight_sums_update_0_write0_merged_banks_2_rst = rst;
  // Bindings to weight_sums_weight_sums_update_0_write0_merged_banks_2

  // Bindings to weight_sums_update_0_write_wen
    // rd_0
  assign rd_0 = weight_sums_update_0_write_wen;

  // selector_bright_weights_normed_rd0_select
  logic [0:0] selector_bright_weights_normed_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_rd0_select_out;
  bright_weights_normed_rd0_select selector_bright_weights_normed_rd0_select(.clk(selector_bright_weights_normed_rd0_select_clk), .rst(selector_bright_weights_normed_rd0_select_rst), .d0(selector_bright_weights_normed_rd0_select_d0), .d1(selector_bright_weights_normed_rd0_select_d1), .out(selector_bright_weights_normed_rd0_select_out));
  assign selector_bright_weights_normed_rd0_select_clk = clk;
  assign selector_bright_weights_normed_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_rd0_select

  // selector_dark_weights_normed_rd0_select
  logic [0:0] selector_dark_weights_normed_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_rd0_select_out;
  dark_weights_normed_rd0_select selector_dark_weights_normed_rd0_select(.clk(selector_dark_weights_normed_rd0_select_clk), .rst(selector_dark_weights_normed_rd0_select_rst), .d0(selector_dark_weights_normed_rd0_select_d0), .d1(selector_dark_weights_normed_rd0_select_d1), .out(selector_dark_weights_normed_rd0_select_out));
  assign selector_dark_weights_normed_rd0_select_clk = clk;
  assign selector_dark_weights_normed_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_rd0_select

  // Bindings to weight_sums_update_0_write_wdata
    // rd_1
  assign rd_1 = weight_sums_update_0_write_wdata;

  // Bindings to bright_weights_normed_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_update_0_read_dummy;

  // Bindings to bright_weights_normed_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_update_0_read_rdata = rd_2;

  // Bindings to dark_weights_normed_update_0_read_dummy
    // rd_4
  assign rd_4 = dark_weights_normed_update_0_read_dummy;

  // Bindings to dark_weights_normed_update_0_read_rdata
    // wr_5
  assign dark_weights_normed_update_0_read_rdata = rd_4;



endmodule


module wire_32(input [31:0] in, output [31:0] out);
  assign out = in;
endmodule


module out_wire_out(input [31:0] out);

endmodule


module bright_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_weights_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module fused_level_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] fused_level_3_update_0_write_wen, input [31:0] fused_level_3_update_0_write_wdata, input [31:0] final_merged_2_update_0_read_dummy, output [31:0] final_merged_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0
  logic [0:0] fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_clk;
  logic [0:0] fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_rst;
  logic [0:0] fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_start;
  logic [0:0] fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_done;
  fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0 fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0(.clk(fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_clk), .rst(fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_rst), .start(fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_start), .done(fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_done));
  assign fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_clk = clk;
  assign fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_rst = rst;
  // Bindings to fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0

  // Bindings to fused_level_3_update_0_write_wen
    // rd_0
  assign rd_0 = fused_level_3_update_0_write_wen;

  // selector_final_merged_2_rd0_select
  logic [0:0] selector_final_merged_2_rd0_select_clk;
  logic [0:0] selector_final_merged_2_rd0_select_rst;
  logic [31:0] selector_final_merged_2_rd0_select_d0;
  logic [31:0] selector_final_merged_2_rd0_select_d1;
  logic [31:0] selector_final_merged_2_rd0_select_out;
  final_merged_2_rd0_select selector_final_merged_2_rd0_select(.clk(selector_final_merged_2_rd0_select_clk), .rst(selector_final_merged_2_rd0_select_rst), .d0(selector_final_merged_2_rd0_select_d0), .d1(selector_final_merged_2_rd0_select_d1), .out(selector_final_merged_2_rd0_select_out));
  assign selector_final_merged_2_rd0_select_clk = clk;
  assign selector_final_merged_2_rd0_select_rst = rst;
  // Bindings to selector_final_merged_2_rd0_select

  // Bindings to fused_level_3_update_0_write_wdata
    // rd_1
  assign rd_1 = fused_level_3_update_0_write_wdata;

  // Bindings to final_merged_2_update_0_read_dummy
    // rd_2
  assign rd_2 = final_merged_2_update_0_read_dummy;

  // Bindings to final_merged_2_update_0_read_rdata
    // wr_3
  assign final_merged_2_update_0_read_rdata = rd_2;



endmodule


module in_off_chip(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] in_update_0_read_dummy, input [0:0] in_off_chip_update_0_write_wen, input [31:0] in_off_chip_update_0_write_wdata, output [31:0] in_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to in_update_0_read_dummy
    // rd_2
  assign rd_2 = in_update_0_read_dummy;

  // Bindings to in_off_chip_update_0_write_wen
    // rd_0
  assign rd_0 = in_off_chip_update_0_write_wen;

  // Bindings to in_off_chip_update_0_write_wdata
    // rd_1
  assign rd_1 = in_off_chip_update_0_write_wdata;

  // Bindings to in_update_0_read_rdata
    // wr_3
  assign in_update_0_read_rdata = rd_2;



endmodule


module in_in_update_0_write0_merged_banks_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_weights_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_gauss_blur_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_gauss_blur_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_laplace_us_0_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_gauss_ds_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_gauss_blur_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_gauss_ds_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module weight_sums_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_gauss_blur_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_laplace_diff_0_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_laplace_us_0_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_gauss_ds_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_gauss_ds_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_gauss_blur_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module bright_gauss_ds_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_laplace_us_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_laplace_diff_0_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_weights_normed_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module bright_weights_normed_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_weights_normed_gauss_blur_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_weights_normed_gauss_ds_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_weights_normed_gauss_blur_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_weights_normed_gauss_blur_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_laplace_us_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_laplace_us_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_weights_normed_gauss_ds_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_gauss_blur_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_laplace_diff_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_weights_normed_gauss_ds_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_weights_normed_gauss_blur_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_laplace_diff_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module fused_level_0_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_laplace_diff_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule



