// Module `hw_kernel_global_wrapper_stencil_ub` defined externally
// Module `hw_input_global_wrapper_stencil_ub` defined externally
// Module `conv_stencil_ub` defined externally
module op_hcompute_hw_output_stencil_write_start_pt__U1941 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_write_start_control_vars_pt__U1944 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_read_start_pt__U1925 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_read_start_control_vars_pt__U1926 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_exe_start_pt__U1927 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U1930 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_7_write_start_pt__U2270 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_7_write_start_control_vars_pt__U2273 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_7_read_start_pt__U2254 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_7_read_start_control_vars_pt__U2255 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_7_exe_start_pt__U2256 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_7_exe_start_control_vars_pt__U2259 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_6_write_start_pt__U2223 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_6_write_start_control_vars_pt__U2226 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_6_read_start_pt__U2207 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_6_read_start_control_vars_pt__U2208 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_6_exe_start_pt__U2209 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_6_exe_start_control_vars_pt__U2212 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_5_write_start_pt__U2176 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_5_write_start_control_vars_pt__U2179 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_5_read_start_pt__U2160 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_5_read_start_control_vars_pt__U2161 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_5_exe_start_pt__U2162 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_5_exe_start_control_vars_pt__U2165 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_4_write_start_pt__U2129 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_4_write_start_control_vars_pt__U2132 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_4_read_start_pt__U2113 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_4_read_start_control_vars_pt__U2114 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_4_exe_start_pt__U2115 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_4_exe_start_control_vars_pt__U2118 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_3_write_start_pt__U2082 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_3_write_start_control_vars_pt__U2085 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_3_read_start_pt__U2066 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_3_read_start_control_vars_pt__U2067 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_3_exe_start_pt__U2068 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_3_exe_start_control_vars_pt__U2071 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_2_write_start_pt__U2035 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_2_write_start_control_vars_pt__U2038 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_2_read_start_pt__U2019 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_2_read_start_control_vars_pt__U2020 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_2_exe_start_pt__U2021 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_2_exe_start_control_vars_pt__U2024 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_1_write_start_pt__U1988 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_1_write_start_control_vars_pt__U1991 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_1_read_start_pt__U1972 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_1_read_start_control_vars_pt__U1973 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_1_exe_start_pt__U1974 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_1_exe_start_control_vars_pt__U1977 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U218 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U219 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U214 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U215 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U216 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U217 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U21 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U22 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U17 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U18 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U19 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U20 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_7_write_start_pt__U182 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_pt__U183 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_7_read_start_pt__U178 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_pt__U179 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_pt__U180 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_pt__U181 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_6_write_start_pt__U159 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_pt__U160 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_6_read_start_pt__U155 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_pt__U156 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_pt__U157 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_pt__U158 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_5_write_start_pt__U136 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_pt__U137 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_5_read_start_pt__U132 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_pt__U133 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_pt__U134 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_pt__U135 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_4_write_start_pt__U113 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_pt__U114 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_4_read_start_pt__U109 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_pt__U110 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_pt__U111 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_pt__U112 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_3_write_start_pt__U90 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_pt__U91 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_3_read_start_pt__U86 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_pt__U87 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_pt__U88 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_pt__U89 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_2_write_start_pt__U67 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_pt__U68 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_2_read_start_pt__U63 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_pt__U64 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_pt__U65 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_pt__U66 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_1_write_start_pt__U44 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_pt__U45 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_1_read_start_pt__U40 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_pt__U41 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_pt__U42 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_pt__U43 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_write_start_pt__U241 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_write_start_control_vars_pt__U242 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_read_start_pt__U237 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_read_start_control_vars_pt__U238 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_exe_start_pt__U239 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_exe_start_control_vars_pt__U240 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_9_write_start_pt__U642 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_9_write_start_control_vars_pt__U660 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_9_read_start_pt__U622 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_9_read_start_control_vars_pt__U623 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_9_exe_start_pt__U624 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_9_exe_start_control_vars_pt__U627 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_8_write_start_pt__U454 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_8_write_start_control_vars_pt__U472 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_8_read_start_pt__U434 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_8_read_start_control_vars_pt__U435 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_8_exe_start_pt__U436 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_8_exe_start_control_vars_pt__U439 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_7_write_start_pt__U402 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_7_write_start_control_vars_pt__U403 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_7_read_start_pt__U398 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_7_read_start_control_vars_pt__U399 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_7_exe_start_pt__U400 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_7_exe_start_control_vars_pt__U401 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_6_write_start_pt__U379 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_6_write_start_control_vars_pt__U380 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_6_read_start_pt__U375 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_6_read_start_control_vars_pt__U376 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_6_exe_start_pt__U377 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_6_exe_start_control_vars_pt__U378 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_write_start_pt__U356 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_write_start_control_vars_pt__U357 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_read_start_pt__U352 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_read_start_control_vars_pt__U353 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_exe_start_pt__U354 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U355 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_write_start_pt__U333 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_write_start_control_vars_pt__U334 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_read_start_pt__U329 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_read_start_control_vars_pt__U330 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_exe_start_pt__U331 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U332 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_write_start_pt__U310 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_write_start_control_vars_pt__U311 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_read_start_pt__U306 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_read_start_control_vars_pt__U307 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_exe_start_pt__U308 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U309 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_write_start_pt__U287 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_write_start_control_vars_pt__U288 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_read_start_pt__U283 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_read_start_control_vars_pt__U284 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_exe_start_pt__U285 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U286 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_write_start_pt__U264 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_write_start_control_vars_pt__U265 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_read_start_pt__U260 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_read_start_control_vars_pt__U261 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_exe_start_pt__U262 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U263 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_15_write_start_pt__U1770 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_15_write_start_control_vars_pt__U1788 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_15_read_start_pt__U1750 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_15_read_start_control_vars_pt__U1751 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_15_exe_start_pt__U1752 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_15_exe_start_control_vars_pt__U1755 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_14_write_start_pt__U1582 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_14_write_start_control_vars_pt__U1600 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_14_read_start_pt__U1562 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_14_read_start_control_vars_pt__U1563 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_14_exe_start_pt__U1564 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_14_exe_start_control_vars_pt__U1567 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_13_write_start_pt__U1394 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_13_write_start_control_vars_pt__U1412 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_13_read_start_pt__U1374 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_13_read_start_control_vars_pt__U1375 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_13_exe_start_pt__U1376 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_13_exe_start_control_vars_pt__U1379 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_12_write_start_pt__U1206 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_12_write_start_control_vars_pt__U1224 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_12_read_start_pt__U1186 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_12_read_start_control_vars_pt__U1187 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_12_exe_start_pt__U1188 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_12_exe_start_control_vars_pt__U1191 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_11_write_start_pt__U1018 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_11_write_start_control_vars_pt__U1036 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_11_read_start_pt__U998 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_11_read_start_control_vars_pt__U999 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_11_exe_start_pt__U1000 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_11_exe_start_control_vars_pt__U1003 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_10_write_start_pt__U830 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_10_write_start_control_vars_pt__U848 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_10_read_start_pt__U810 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_10_read_start_control_vars_pt__U811 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_10_exe_start_pt__U812 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_10_exe_start_control_vars_pt__U815 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module coreir_reg #(
    parameter width = 1,
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input [width-1:0] in,
    output [width-1:0] out
);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out
);
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(clk),
    .in(in),
    .out(out)
);
endmodule

module mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out,
    input en
);
wire [15:0] enMux_out;
assign enMux_out = en ? in : out;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(clk),
    .in(enMux_out),
    .out(out)
);
endmodule

module corebit_reg #(
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input in,
    output out
);
reg outReg = init;
always @(posedge clk) begin
  outReg <= in;
end
assign out = outReg;
endmodule

module array_delay_U962 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U963_out;
wire [15:0] _U964_out;
wire [15:0] _U965_out;
wire [15:0] _U966_out;
wire [15:0] _U967_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U963 (
    .in(in[0]),
    .clk(clk),
    .out(_U963_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U964 (
    .in(in[1]),
    .clk(clk),
    .out(_U964_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U965 (
    .in(in[2]),
    .clk(clk),
    .out(_U965_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U966 (
    .in(in[3]),
    .clk(clk),
    .out(_U966_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U967 (
    .in(in[4]),
    .clk(clk),
    .out(_U967_out)
);
assign out[4] = _U967_out;
assign out[3] = _U966_out;
assign out[2] = _U965_out;
assign out[1] = _U964_out;
assign out[0] = _U963_out;
endmodule

module array_delay_U955 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U956_out;
wire [15:0] _U957_out;
wire [15:0] _U958_out;
wire [15:0] _U959_out;
wire [15:0] _U960_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U956 (
    .in(in[0]),
    .clk(clk),
    .out(_U956_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U957 (
    .in(in[1]),
    .clk(clk),
    .out(_U957_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U958 (
    .in(in[2]),
    .clk(clk),
    .out(_U958_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U959 (
    .in(in[3]),
    .clk(clk),
    .out(_U959_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U960 (
    .in(in[4]),
    .clk(clk),
    .out(_U960_out)
);
assign out[4] = _U960_out;
assign out[3] = _U959_out;
assign out[2] = _U958_out;
assign out[1] = _U957_out;
assign out[0] = _U956_out;
endmodule

module array_delay_U948 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U949_out;
wire [15:0] _U950_out;
wire [15:0] _U951_out;
wire [15:0] _U952_out;
wire [15:0] _U953_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U949 (
    .in(in[0]),
    .clk(clk),
    .out(_U949_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U950 (
    .in(in[1]),
    .clk(clk),
    .out(_U950_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U951 (
    .in(in[2]),
    .clk(clk),
    .out(_U951_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U952 (
    .in(in[3]),
    .clk(clk),
    .out(_U952_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U953 (
    .in(in[4]),
    .clk(clk),
    .out(_U953_out)
);
assign out[4] = _U953_out;
assign out[3] = _U952_out;
assign out[2] = _U951_out;
assign out[1] = _U950_out;
assign out[0] = _U949_out;
endmodule

module array_delay_U941 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U942_out;
wire [15:0] _U943_out;
wire [15:0] _U944_out;
wire [15:0] _U945_out;
wire [15:0] _U946_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U942 (
    .in(in[0]),
    .clk(clk),
    .out(_U942_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U943 (
    .in(in[1]),
    .clk(clk),
    .out(_U943_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U944 (
    .in(in[2]),
    .clk(clk),
    .out(_U944_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U945 (
    .in(in[3]),
    .clk(clk),
    .out(_U945_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U946 (
    .in(in[4]),
    .clk(clk),
    .out(_U946_out)
);
assign out[4] = _U946_out;
assign out[3] = _U945_out;
assign out[2] = _U944_out;
assign out[1] = _U943_out;
assign out[0] = _U942_out;
endmodule

module array_delay_U934 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U935_out;
wire [15:0] _U936_out;
wire [15:0] _U937_out;
wire [15:0] _U938_out;
wire [15:0] _U939_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U935 (
    .in(in[0]),
    .clk(clk),
    .out(_U935_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U936 (
    .in(in[1]),
    .clk(clk),
    .out(_U936_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U937 (
    .in(in[2]),
    .clk(clk),
    .out(_U937_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U938 (
    .in(in[3]),
    .clk(clk),
    .out(_U938_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U939 (
    .in(in[4]),
    .clk(clk),
    .out(_U939_out)
);
assign out[4] = _U939_out;
assign out[3] = _U938_out;
assign out[2] = _U937_out;
assign out[1] = _U936_out;
assign out[0] = _U935_out;
endmodule

module array_delay_U927 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U928_out;
wire [15:0] _U929_out;
wire [15:0] _U930_out;
wire [15:0] _U931_out;
wire [15:0] _U932_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U928 (
    .in(in[0]),
    .clk(clk),
    .out(_U928_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U929 (
    .in(in[1]),
    .clk(clk),
    .out(_U929_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U930 (
    .in(in[2]),
    .clk(clk),
    .out(_U930_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U931 (
    .in(in[3]),
    .clk(clk),
    .out(_U931_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U932 (
    .in(in[4]),
    .clk(clk),
    .out(_U932_out)
);
assign out[4] = _U932_out;
assign out[3] = _U931_out;
assign out[2] = _U930_out;
assign out[1] = _U929_out;
assign out[0] = _U928_out;
endmodule

module array_delay_U920 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U921_out;
wire [15:0] _U922_out;
wire [15:0] _U923_out;
wire [15:0] _U924_out;
wire [15:0] _U925_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U921 (
    .in(in[0]),
    .clk(clk),
    .out(_U921_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U922 (
    .in(in[1]),
    .clk(clk),
    .out(_U922_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U923 (
    .in(in[2]),
    .clk(clk),
    .out(_U923_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U924 (
    .in(in[3]),
    .clk(clk),
    .out(_U924_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U925 (
    .in(in[4]),
    .clk(clk),
    .out(_U925_out)
);
assign out[4] = _U925_out;
assign out[3] = _U924_out;
assign out[2] = _U923_out;
assign out[1] = _U922_out;
assign out[0] = _U921_out;
endmodule

module array_delay_U913 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U914_out;
wire [15:0] _U915_out;
wire [15:0] _U916_out;
wire [15:0] _U917_out;
wire [15:0] _U918_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U914 (
    .in(in[0]),
    .clk(clk),
    .out(_U914_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U915 (
    .in(in[1]),
    .clk(clk),
    .out(_U915_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U916 (
    .in(in[2]),
    .clk(clk),
    .out(_U916_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U917 (
    .in(in[3]),
    .clk(clk),
    .out(_U917_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U918 (
    .in(in[4]),
    .clk(clk),
    .out(_U918_out)
);
assign out[4] = _U918_out;
assign out[3] = _U917_out;
assign out[2] = _U916_out;
assign out[1] = _U915_out;
assign out[0] = _U914_out;
endmodule

module array_delay_U906 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U907_out;
wire [15:0] _U908_out;
wire [15:0] _U909_out;
wire [15:0] _U910_out;
wire [15:0] _U911_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U907 (
    .in(in[0]),
    .clk(clk),
    .out(_U907_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U908 (
    .in(in[1]),
    .clk(clk),
    .out(_U908_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U909 (
    .in(in[2]),
    .clk(clk),
    .out(_U909_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U910 (
    .in(in[3]),
    .clk(clk),
    .out(_U910_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U911 (
    .in(in[4]),
    .clk(clk),
    .out(_U911_out)
);
assign out[4] = _U911_out;
assign out[3] = _U910_out;
assign out[2] = _U909_out;
assign out[1] = _U908_out;
assign out[0] = _U907_out;
endmodule

module array_delay_U899 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U900_out;
wire [15:0] _U901_out;
wire [15:0] _U902_out;
wire [15:0] _U903_out;
wire [15:0] _U904_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U900 (
    .in(in[0]),
    .clk(clk),
    .out(_U900_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U901 (
    .in(in[1]),
    .clk(clk),
    .out(_U901_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U902 (
    .in(in[2]),
    .clk(clk),
    .out(_U902_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U903 (
    .in(in[3]),
    .clk(clk),
    .out(_U903_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U904 (
    .in(in[4]),
    .clk(clk),
    .out(_U904_out)
);
assign out[4] = _U904_out;
assign out[3] = _U903_out;
assign out[2] = _U902_out;
assign out[1] = _U901_out;
assign out[0] = _U900_out;
endmodule

module array_delay_U892 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U893_out;
wire [15:0] _U894_out;
wire [15:0] _U895_out;
wire [15:0] _U896_out;
wire [15:0] _U897_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U893 (
    .in(in[0]),
    .clk(clk),
    .out(_U893_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U894 (
    .in(in[1]),
    .clk(clk),
    .out(_U894_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U895 (
    .in(in[2]),
    .clk(clk),
    .out(_U895_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U896 (
    .in(in[3]),
    .clk(clk),
    .out(_U896_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U897 (
    .in(in[4]),
    .clk(clk),
    .out(_U897_out)
);
assign out[4] = _U897_out;
assign out[3] = _U896_out;
assign out[2] = _U895_out;
assign out[1] = _U894_out;
assign out[0] = _U893_out;
endmodule

module array_delay_U885 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U886_out;
wire [15:0] _U887_out;
wire [15:0] _U888_out;
wire [15:0] _U889_out;
wire [15:0] _U890_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U886 (
    .in(in[0]),
    .clk(clk),
    .out(_U886_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U887 (
    .in(in[1]),
    .clk(clk),
    .out(_U887_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U888 (
    .in(in[2]),
    .clk(clk),
    .out(_U888_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U889 (
    .in(in[3]),
    .clk(clk),
    .out(_U889_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U890 (
    .in(in[4]),
    .clk(clk),
    .out(_U890_out)
);
assign out[4] = _U890_out;
assign out[3] = _U889_out;
assign out[2] = _U888_out;
assign out[1] = _U887_out;
assign out[0] = _U886_out;
endmodule

module array_delay_U878 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U879_out;
wire [15:0] _U880_out;
wire [15:0] _U881_out;
wire [15:0] _U882_out;
wire [15:0] _U883_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U879 (
    .in(in[0]),
    .clk(clk),
    .out(_U879_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U880 (
    .in(in[1]),
    .clk(clk),
    .out(_U880_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U881 (
    .in(in[2]),
    .clk(clk),
    .out(_U881_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U882 (
    .in(in[3]),
    .clk(clk),
    .out(_U882_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U883 (
    .in(in[4]),
    .clk(clk),
    .out(_U883_out)
);
assign out[4] = _U883_out;
assign out[3] = _U882_out;
assign out[2] = _U881_out;
assign out[1] = _U880_out;
assign out[0] = _U879_out;
endmodule

module array_delay_U871 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U872_out;
wire [15:0] _U873_out;
wire [15:0] _U874_out;
wire [15:0] _U875_out;
wire [15:0] _U876_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U872 (
    .in(in[0]),
    .clk(clk),
    .out(_U872_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U873 (
    .in(in[1]),
    .clk(clk),
    .out(_U873_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U874 (
    .in(in[2]),
    .clk(clk),
    .out(_U874_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U875 (
    .in(in[3]),
    .clk(clk),
    .out(_U875_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U876 (
    .in(in[4]),
    .clk(clk),
    .out(_U876_out)
);
assign out[4] = _U876_out;
assign out[3] = _U875_out;
assign out[2] = _U874_out;
assign out[1] = _U873_out;
assign out[0] = _U872_out;
endmodule

module array_delay_U864 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U865_out;
wire [15:0] _U866_out;
wire [15:0] _U867_out;
wire [15:0] _U868_out;
wire [15:0] _U869_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U865 (
    .in(in[0]),
    .clk(clk),
    .out(_U865_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U866 (
    .in(in[1]),
    .clk(clk),
    .out(_U866_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U867 (
    .in(in[2]),
    .clk(clk),
    .out(_U867_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U868 (
    .in(in[3]),
    .clk(clk),
    .out(_U868_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U869 (
    .in(in[4]),
    .clk(clk),
    .out(_U869_out)
);
assign out[4] = _U869_out;
assign out[3] = _U868_out;
assign out[2] = _U867_out;
assign out[1] = _U866_out;
assign out[0] = _U865_out;
endmodule

module array_delay_U857 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U858_out;
wire [15:0] _U859_out;
wire [15:0] _U860_out;
wire [15:0] _U861_out;
wire [15:0] _U862_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U858 (
    .in(in[0]),
    .clk(clk),
    .out(_U858_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U859 (
    .in(in[1]),
    .clk(clk),
    .out(_U859_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U860 (
    .in(in[2]),
    .clk(clk),
    .out(_U860_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U861 (
    .in(in[3]),
    .clk(clk),
    .out(_U861_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U862 (
    .in(in[4]),
    .clk(clk),
    .out(_U862_out)
);
assign out[4] = _U862_out;
assign out[3] = _U861_out;
assign out[2] = _U860_out;
assign out[1] = _U859_out;
assign out[0] = _U858_out;
endmodule

module array_delay_U850 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U851_out;
wire [15:0] _U852_out;
wire [15:0] _U853_out;
wire [15:0] _U854_out;
wire [15:0] _U855_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U851 (
    .in(in[0]),
    .clk(clk),
    .out(_U851_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U852 (
    .in(in[1]),
    .clk(clk),
    .out(_U852_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U853 (
    .in(in[2]),
    .clk(clk),
    .out(_U853_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U854 (
    .in(in[3]),
    .clk(clk),
    .out(_U854_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U855 (
    .in(in[4]),
    .clk(clk),
    .out(_U855_out)
);
assign out[4] = _U855_out;
assign out[3] = _U854_out;
assign out[2] = _U853_out;
assign out[1] = _U852_out;
assign out[0] = _U851_out;
endmodule

module array_delay_U824 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U825_out;
wire [15:0] _U826_out;
wire [15:0] _U827_out;
wire [15:0] _U828_out;
wire [15:0] _U829_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U825 (
    .in(in[0]),
    .clk(clk),
    .out(_U825_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U826 (
    .in(in[1]),
    .clk(clk),
    .out(_U826_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U827 (
    .in(in[2]),
    .clk(clk),
    .out(_U827_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U828 (
    .in(in[3]),
    .clk(clk),
    .out(_U828_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U829 (
    .in(in[4]),
    .clk(clk),
    .out(_U829_out)
);
assign out[4] = _U829_out;
assign out[3] = _U828_out;
assign out[2] = _U827_out;
assign out[1] = _U826_out;
assign out[0] = _U825_out;
endmodule

module array_delay_U817 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U818_out;
wire [15:0] _U819_out;
wire [15:0] _U820_out;
wire [15:0] _U821_out;
wire [15:0] _U822_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U818 (
    .in(in[0]),
    .clk(clk),
    .out(_U818_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U819 (
    .in(in[1]),
    .clk(clk),
    .out(_U819_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U820 (
    .in(in[2]),
    .clk(clk),
    .out(_U820_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U821 (
    .in(in[3]),
    .clk(clk),
    .out(_U821_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U822 (
    .in(in[4]),
    .clk(clk),
    .out(_U822_out)
);
assign out[4] = _U822_out;
assign out[3] = _U821_out;
assign out[2] = _U820_out;
assign out[1] = _U819_out;
assign out[0] = _U818_out;
endmodule

module array_delay_U774 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U775_out;
wire [15:0] _U776_out;
wire [15:0] _U777_out;
wire [15:0] _U778_out;
wire [15:0] _U779_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U775 (
    .in(in[0]),
    .clk(clk),
    .out(_U775_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U776 (
    .in(in[1]),
    .clk(clk),
    .out(_U776_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U777 (
    .in(in[2]),
    .clk(clk),
    .out(_U777_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U778 (
    .in(in[3]),
    .clk(clk),
    .out(_U778_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U779 (
    .in(in[4]),
    .clk(clk),
    .out(_U779_out)
);
assign out[4] = _U779_out;
assign out[3] = _U778_out;
assign out[2] = _U777_out;
assign out[1] = _U776_out;
assign out[0] = _U775_out;
endmodule

module array_delay_U767 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U768_out;
wire [15:0] _U769_out;
wire [15:0] _U770_out;
wire [15:0] _U771_out;
wire [15:0] _U772_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U768 (
    .in(in[0]),
    .clk(clk),
    .out(_U768_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U769 (
    .in(in[1]),
    .clk(clk),
    .out(_U769_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U770 (
    .in(in[2]),
    .clk(clk),
    .out(_U770_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U771 (
    .in(in[3]),
    .clk(clk),
    .out(_U771_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U772 (
    .in(in[4]),
    .clk(clk),
    .out(_U772_out)
);
assign out[4] = _U772_out;
assign out[3] = _U771_out;
assign out[2] = _U770_out;
assign out[1] = _U769_out;
assign out[0] = _U768_out;
endmodule

module array_delay_U760 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U761_out;
wire [15:0] _U762_out;
wire [15:0] _U763_out;
wire [15:0] _U764_out;
wire [15:0] _U765_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U761 (
    .in(in[0]),
    .clk(clk),
    .out(_U761_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U762 (
    .in(in[1]),
    .clk(clk),
    .out(_U762_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U763 (
    .in(in[2]),
    .clk(clk),
    .out(_U763_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U764 (
    .in(in[3]),
    .clk(clk),
    .out(_U764_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U765 (
    .in(in[4]),
    .clk(clk),
    .out(_U765_out)
);
assign out[4] = _U765_out;
assign out[3] = _U764_out;
assign out[2] = _U763_out;
assign out[1] = _U762_out;
assign out[0] = _U761_out;
endmodule

module array_delay_U753 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U754_out;
wire [15:0] _U755_out;
wire [15:0] _U756_out;
wire [15:0] _U757_out;
wire [15:0] _U758_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U754 (
    .in(in[0]),
    .clk(clk),
    .out(_U754_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U755 (
    .in(in[1]),
    .clk(clk),
    .out(_U755_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U756 (
    .in(in[2]),
    .clk(clk),
    .out(_U756_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U757 (
    .in(in[3]),
    .clk(clk),
    .out(_U757_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U758 (
    .in(in[4]),
    .clk(clk),
    .out(_U758_out)
);
assign out[4] = _U758_out;
assign out[3] = _U757_out;
assign out[2] = _U756_out;
assign out[1] = _U755_out;
assign out[0] = _U754_out;
endmodule

module array_delay_U746 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U747_out;
wire [15:0] _U748_out;
wire [15:0] _U749_out;
wire [15:0] _U750_out;
wire [15:0] _U751_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U747 (
    .in(in[0]),
    .clk(clk),
    .out(_U747_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U748 (
    .in(in[1]),
    .clk(clk),
    .out(_U748_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U749 (
    .in(in[2]),
    .clk(clk),
    .out(_U749_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U750 (
    .in(in[3]),
    .clk(clk),
    .out(_U750_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U751 (
    .in(in[4]),
    .clk(clk),
    .out(_U751_out)
);
assign out[4] = _U751_out;
assign out[3] = _U750_out;
assign out[2] = _U749_out;
assign out[1] = _U748_out;
assign out[0] = _U747_out;
endmodule

module array_delay_U739 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U740_out;
wire [15:0] _U741_out;
wire [15:0] _U742_out;
wire [15:0] _U743_out;
wire [15:0] _U744_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U740 (
    .in(in[0]),
    .clk(clk),
    .out(_U740_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U741 (
    .in(in[1]),
    .clk(clk),
    .out(_U741_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U742 (
    .in(in[2]),
    .clk(clk),
    .out(_U742_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U743 (
    .in(in[3]),
    .clk(clk),
    .out(_U743_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U744 (
    .in(in[4]),
    .clk(clk),
    .out(_U744_out)
);
assign out[4] = _U744_out;
assign out[3] = _U743_out;
assign out[2] = _U742_out;
assign out[1] = _U741_out;
assign out[0] = _U740_out;
endmodule

module array_delay_U732 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U733_out;
wire [15:0] _U734_out;
wire [15:0] _U735_out;
wire [15:0] _U736_out;
wire [15:0] _U737_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U733 (
    .in(in[0]),
    .clk(clk),
    .out(_U733_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U734 (
    .in(in[1]),
    .clk(clk),
    .out(_U734_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U735 (
    .in(in[2]),
    .clk(clk),
    .out(_U735_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U736 (
    .in(in[3]),
    .clk(clk),
    .out(_U736_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U737 (
    .in(in[4]),
    .clk(clk),
    .out(_U737_out)
);
assign out[4] = _U737_out;
assign out[3] = _U736_out;
assign out[2] = _U735_out;
assign out[1] = _U734_out;
assign out[0] = _U733_out;
endmodule

module array_delay_U725 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U726_out;
wire [15:0] _U727_out;
wire [15:0] _U728_out;
wire [15:0] _U729_out;
wire [15:0] _U730_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U726 (
    .in(in[0]),
    .clk(clk),
    .out(_U726_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U727 (
    .in(in[1]),
    .clk(clk),
    .out(_U727_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U728 (
    .in(in[2]),
    .clk(clk),
    .out(_U728_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U729 (
    .in(in[3]),
    .clk(clk),
    .out(_U729_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U730 (
    .in(in[4]),
    .clk(clk),
    .out(_U730_out)
);
assign out[4] = _U730_out;
assign out[3] = _U729_out;
assign out[2] = _U728_out;
assign out[1] = _U727_out;
assign out[0] = _U726_out;
endmodule

module array_delay_U718 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U719_out;
wire [15:0] _U720_out;
wire [15:0] _U721_out;
wire [15:0] _U722_out;
wire [15:0] _U723_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U719 (
    .in(in[0]),
    .clk(clk),
    .out(_U719_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U720 (
    .in(in[1]),
    .clk(clk),
    .out(_U720_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U721 (
    .in(in[2]),
    .clk(clk),
    .out(_U721_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U722 (
    .in(in[3]),
    .clk(clk),
    .out(_U722_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U723 (
    .in(in[4]),
    .clk(clk),
    .out(_U723_out)
);
assign out[4] = _U723_out;
assign out[3] = _U722_out;
assign out[2] = _U721_out;
assign out[1] = _U720_out;
assign out[0] = _U719_out;
endmodule

module array_delay_U711 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U712_out;
wire [15:0] _U713_out;
wire [15:0] _U714_out;
wire [15:0] _U715_out;
wire [15:0] _U716_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U712 (
    .in(in[0]),
    .clk(clk),
    .out(_U712_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U713 (
    .in(in[1]),
    .clk(clk),
    .out(_U713_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U714 (
    .in(in[2]),
    .clk(clk),
    .out(_U714_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U715 (
    .in(in[3]),
    .clk(clk),
    .out(_U715_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U716 (
    .in(in[4]),
    .clk(clk),
    .out(_U716_out)
);
assign out[4] = _U716_out;
assign out[3] = _U715_out;
assign out[2] = _U714_out;
assign out[1] = _U713_out;
assign out[0] = _U712_out;
endmodule

module array_delay_U704 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U705_out;
wire [15:0] _U706_out;
wire [15:0] _U707_out;
wire [15:0] _U708_out;
wire [15:0] _U709_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U705 (
    .in(in[0]),
    .clk(clk),
    .out(_U705_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U706 (
    .in(in[1]),
    .clk(clk),
    .out(_U706_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U707 (
    .in(in[2]),
    .clk(clk),
    .out(_U707_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U708 (
    .in(in[3]),
    .clk(clk),
    .out(_U708_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U709 (
    .in(in[4]),
    .clk(clk),
    .out(_U709_out)
);
assign out[4] = _U709_out;
assign out[3] = _U708_out;
assign out[2] = _U707_out;
assign out[1] = _U706_out;
assign out[0] = _U705_out;
endmodule

module array_delay_U697 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U698_out;
wire [15:0] _U699_out;
wire [15:0] _U700_out;
wire [15:0] _U701_out;
wire [15:0] _U702_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U698 (
    .in(in[0]),
    .clk(clk),
    .out(_U698_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U699 (
    .in(in[1]),
    .clk(clk),
    .out(_U699_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U700 (
    .in(in[2]),
    .clk(clk),
    .out(_U700_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U701 (
    .in(in[3]),
    .clk(clk),
    .out(_U701_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U702 (
    .in(in[4]),
    .clk(clk),
    .out(_U702_out)
);
assign out[4] = _U702_out;
assign out[3] = _U701_out;
assign out[2] = _U700_out;
assign out[1] = _U699_out;
assign out[0] = _U698_out;
endmodule

module array_delay_U690 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U691_out;
wire [15:0] _U692_out;
wire [15:0] _U693_out;
wire [15:0] _U694_out;
wire [15:0] _U695_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U691 (
    .in(in[0]),
    .clk(clk),
    .out(_U691_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U692 (
    .in(in[1]),
    .clk(clk),
    .out(_U692_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U693 (
    .in(in[2]),
    .clk(clk),
    .out(_U693_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U694 (
    .in(in[3]),
    .clk(clk),
    .out(_U694_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U695 (
    .in(in[4]),
    .clk(clk),
    .out(_U695_out)
);
assign out[4] = _U695_out;
assign out[3] = _U694_out;
assign out[2] = _U693_out;
assign out[1] = _U692_out;
assign out[0] = _U691_out;
endmodule

module array_delay_U683 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U684_out;
wire [15:0] _U685_out;
wire [15:0] _U686_out;
wire [15:0] _U687_out;
wire [15:0] _U688_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U684 (
    .in(in[0]),
    .clk(clk),
    .out(_U684_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U685 (
    .in(in[1]),
    .clk(clk),
    .out(_U685_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U686 (
    .in(in[2]),
    .clk(clk),
    .out(_U686_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U687 (
    .in(in[3]),
    .clk(clk),
    .out(_U687_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U688 (
    .in(in[4]),
    .clk(clk),
    .out(_U688_out)
);
assign out[4] = _U688_out;
assign out[3] = _U687_out;
assign out[2] = _U686_out;
assign out[1] = _U685_out;
assign out[0] = _U684_out;
endmodule

module array_delay_U676 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U677_out;
wire [15:0] _U678_out;
wire [15:0] _U679_out;
wire [15:0] _U680_out;
wire [15:0] _U681_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U677 (
    .in(in[0]),
    .clk(clk),
    .out(_U677_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U678 (
    .in(in[1]),
    .clk(clk),
    .out(_U678_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U679 (
    .in(in[2]),
    .clk(clk),
    .out(_U679_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U680 (
    .in(in[3]),
    .clk(clk),
    .out(_U680_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U681 (
    .in(in[4]),
    .clk(clk),
    .out(_U681_out)
);
assign out[4] = _U681_out;
assign out[3] = _U680_out;
assign out[2] = _U679_out;
assign out[1] = _U678_out;
assign out[0] = _U677_out;
endmodule

module array_delay_U669 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U670_out;
wire [15:0] _U671_out;
wire [15:0] _U672_out;
wire [15:0] _U673_out;
wire [15:0] _U674_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U670 (
    .in(in[0]),
    .clk(clk),
    .out(_U670_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U671 (
    .in(in[1]),
    .clk(clk),
    .out(_U671_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U672 (
    .in(in[2]),
    .clk(clk),
    .out(_U672_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U673 (
    .in(in[3]),
    .clk(clk),
    .out(_U673_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U674 (
    .in(in[4]),
    .clk(clk),
    .out(_U674_out)
);
assign out[4] = _U674_out;
assign out[3] = _U673_out;
assign out[2] = _U672_out;
assign out[1] = _U671_out;
assign out[0] = _U670_out;
endmodule

module array_delay_U662 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U663_out;
wire [15:0] _U664_out;
wire [15:0] _U665_out;
wire [15:0] _U666_out;
wire [15:0] _U667_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U663 (
    .in(in[0]),
    .clk(clk),
    .out(_U663_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U664 (
    .in(in[1]),
    .clk(clk),
    .out(_U664_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U665 (
    .in(in[2]),
    .clk(clk),
    .out(_U665_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U666 (
    .in(in[3]),
    .clk(clk),
    .out(_U666_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U667 (
    .in(in[4]),
    .clk(clk),
    .out(_U667_out)
);
assign out[4] = _U667_out;
assign out[3] = _U666_out;
assign out[2] = _U665_out;
assign out[1] = _U664_out;
assign out[0] = _U663_out;
endmodule

module array_delay_U636 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U637_out;
wire [15:0] _U638_out;
wire [15:0] _U639_out;
wire [15:0] _U640_out;
wire [15:0] _U641_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U637 (
    .in(in[0]),
    .clk(clk),
    .out(_U637_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U638 (
    .in(in[1]),
    .clk(clk),
    .out(_U638_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U639 (
    .in(in[2]),
    .clk(clk),
    .out(_U639_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U640 (
    .in(in[3]),
    .clk(clk),
    .out(_U640_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U641 (
    .in(in[4]),
    .clk(clk),
    .out(_U641_out)
);
assign out[4] = _U641_out;
assign out[3] = _U640_out;
assign out[2] = _U639_out;
assign out[1] = _U638_out;
assign out[0] = _U637_out;
endmodule

module array_delay_U629 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U630_out;
wire [15:0] _U631_out;
wire [15:0] _U632_out;
wire [15:0] _U633_out;
wire [15:0] _U634_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U630 (
    .in(in[0]),
    .clk(clk),
    .out(_U630_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U631 (
    .in(in[1]),
    .clk(clk),
    .out(_U631_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U632 (
    .in(in[2]),
    .clk(clk),
    .out(_U632_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U633 (
    .in(in[3]),
    .clk(clk),
    .out(_U633_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U634 (
    .in(in[4]),
    .clk(clk),
    .out(_U634_out)
);
assign out[4] = _U634_out;
assign out[3] = _U633_out;
assign out[2] = _U632_out;
assign out[1] = _U631_out;
assign out[0] = _U630_out;
endmodule

module array_delay_U586 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U587_out;
wire [15:0] _U588_out;
wire [15:0] _U589_out;
wire [15:0] _U590_out;
wire [15:0] _U591_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U587 (
    .in(in[0]),
    .clk(clk),
    .out(_U587_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U588 (
    .in(in[1]),
    .clk(clk),
    .out(_U588_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U589 (
    .in(in[2]),
    .clk(clk),
    .out(_U589_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U590 (
    .in(in[3]),
    .clk(clk),
    .out(_U590_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U591 (
    .in(in[4]),
    .clk(clk),
    .out(_U591_out)
);
assign out[4] = _U591_out;
assign out[3] = _U590_out;
assign out[2] = _U589_out;
assign out[1] = _U588_out;
assign out[0] = _U587_out;
endmodule

module array_delay_U579 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U580_out;
wire [15:0] _U581_out;
wire [15:0] _U582_out;
wire [15:0] _U583_out;
wire [15:0] _U584_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U580 (
    .in(in[0]),
    .clk(clk),
    .out(_U580_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U581 (
    .in(in[1]),
    .clk(clk),
    .out(_U581_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U582 (
    .in(in[2]),
    .clk(clk),
    .out(_U582_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U583 (
    .in(in[3]),
    .clk(clk),
    .out(_U583_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U584 (
    .in(in[4]),
    .clk(clk),
    .out(_U584_out)
);
assign out[4] = _U584_out;
assign out[3] = _U583_out;
assign out[2] = _U582_out;
assign out[1] = _U581_out;
assign out[0] = _U580_out;
endmodule

module array_delay_U572 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U573_out;
wire [15:0] _U574_out;
wire [15:0] _U575_out;
wire [15:0] _U576_out;
wire [15:0] _U577_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U573 (
    .in(in[0]),
    .clk(clk),
    .out(_U573_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U574 (
    .in(in[1]),
    .clk(clk),
    .out(_U574_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U575 (
    .in(in[2]),
    .clk(clk),
    .out(_U575_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U576 (
    .in(in[3]),
    .clk(clk),
    .out(_U576_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U577 (
    .in(in[4]),
    .clk(clk),
    .out(_U577_out)
);
assign out[4] = _U577_out;
assign out[3] = _U576_out;
assign out[2] = _U575_out;
assign out[1] = _U574_out;
assign out[0] = _U573_out;
endmodule

module array_delay_U565 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U566_out;
wire [15:0] _U567_out;
wire [15:0] _U568_out;
wire [15:0] _U569_out;
wire [15:0] _U570_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U566 (
    .in(in[0]),
    .clk(clk),
    .out(_U566_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U567 (
    .in(in[1]),
    .clk(clk),
    .out(_U567_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U568 (
    .in(in[2]),
    .clk(clk),
    .out(_U568_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U569 (
    .in(in[3]),
    .clk(clk),
    .out(_U569_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U570 (
    .in(in[4]),
    .clk(clk),
    .out(_U570_out)
);
assign out[4] = _U570_out;
assign out[3] = _U569_out;
assign out[2] = _U568_out;
assign out[1] = _U567_out;
assign out[0] = _U566_out;
endmodule

module array_delay_U558 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U559_out;
wire [15:0] _U560_out;
wire [15:0] _U561_out;
wire [15:0] _U562_out;
wire [15:0] _U563_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U559 (
    .in(in[0]),
    .clk(clk),
    .out(_U559_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U560 (
    .in(in[1]),
    .clk(clk),
    .out(_U560_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U561 (
    .in(in[2]),
    .clk(clk),
    .out(_U561_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U562 (
    .in(in[3]),
    .clk(clk),
    .out(_U562_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U563 (
    .in(in[4]),
    .clk(clk),
    .out(_U563_out)
);
assign out[4] = _U563_out;
assign out[3] = _U562_out;
assign out[2] = _U561_out;
assign out[1] = _U560_out;
assign out[0] = _U559_out;
endmodule

module array_delay_U551 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U552_out;
wire [15:0] _U553_out;
wire [15:0] _U554_out;
wire [15:0] _U555_out;
wire [15:0] _U556_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U552 (
    .in(in[0]),
    .clk(clk),
    .out(_U552_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U553 (
    .in(in[1]),
    .clk(clk),
    .out(_U553_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U554 (
    .in(in[2]),
    .clk(clk),
    .out(_U554_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U555 (
    .in(in[3]),
    .clk(clk),
    .out(_U555_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U556 (
    .in(in[4]),
    .clk(clk),
    .out(_U556_out)
);
assign out[4] = _U556_out;
assign out[3] = _U555_out;
assign out[2] = _U554_out;
assign out[1] = _U553_out;
assign out[0] = _U552_out;
endmodule

module array_delay_U544 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U545_out;
wire [15:0] _U546_out;
wire [15:0] _U547_out;
wire [15:0] _U548_out;
wire [15:0] _U549_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U545 (
    .in(in[0]),
    .clk(clk),
    .out(_U545_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U546 (
    .in(in[1]),
    .clk(clk),
    .out(_U546_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U547 (
    .in(in[2]),
    .clk(clk),
    .out(_U547_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U548 (
    .in(in[3]),
    .clk(clk),
    .out(_U548_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U549 (
    .in(in[4]),
    .clk(clk),
    .out(_U549_out)
);
assign out[4] = _U549_out;
assign out[3] = _U548_out;
assign out[2] = _U547_out;
assign out[1] = _U546_out;
assign out[0] = _U545_out;
endmodule

module array_delay_U537 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U538_out;
wire [15:0] _U539_out;
wire [15:0] _U540_out;
wire [15:0] _U541_out;
wire [15:0] _U542_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U538 (
    .in(in[0]),
    .clk(clk),
    .out(_U538_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U539 (
    .in(in[1]),
    .clk(clk),
    .out(_U539_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U540 (
    .in(in[2]),
    .clk(clk),
    .out(_U540_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U541 (
    .in(in[3]),
    .clk(clk),
    .out(_U541_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U542 (
    .in(in[4]),
    .clk(clk),
    .out(_U542_out)
);
assign out[4] = _U542_out;
assign out[3] = _U541_out;
assign out[2] = _U540_out;
assign out[1] = _U539_out;
assign out[0] = _U538_out;
endmodule

module array_delay_U530 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U531_out;
wire [15:0] _U532_out;
wire [15:0] _U533_out;
wire [15:0] _U534_out;
wire [15:0] _U535_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U531 (
    .in(in[0]),
    .clk(clk),
    .out(_U531_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U532 (
    .in(in[1]),
    .clk(clk),
    .out(_U532_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U533 (
    .in(in[2]),
    .clk(clk),
    .out(_U533_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U534 (
    .in(in[3]),
    .clk(clk),
    .out(_U534_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U535 (
    .in(in[4]),
    .clk(clk),
    .out(_U535_out)
);
assign out[4] = _U535_out;
assign out[3] = _U534_out;
assign out[2] = _U533_out;
assign out[1] = _U532_out;
assign out[0] = _U531_out;
endmodule

module array_delay_U523 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U524_out;
wire [15:0] _U525_out;
wire [15:0] _U526_out;
wire [15:0] _U527_out;
wire [15:0] _U528_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U524 (
    .in(in[0]),
    .clk(clk),
    .out(_U524_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U525 (
    .in(in[1]),
    .clk(clk),
    .out(_U525_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U526 (
    .in(in[2]),
    .clk(clk),
    .out(_U526_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U527 (
    .in(in[3]),
    .clk(clk),
    .out(_U527_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U528 (
    .in(in[4]),
    .clk(clk),
    .out(_U528_out)
);
assign out[4] = _U528_out;
assign out[3] = _U527_out;
assign out[2] = _U526_out;
assign out[1] = _U525_out;
assign out[0] = _U524_out;
endmodule

module array_delay_U516 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U517_out;
wire [15:0] _U518_out;
wire [15:0] _U519_out;
wire [15:0] _U520_out;
wire [15:0] _U521_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U517 (
    .in(in[0]),
    .clk(clk),
    .out(_U517_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U518 (
    .in(in[1]),
    .clk(clk),
    .out(_U518_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U519 (
    .in(in[2]),
    .clk(clk),
    .out(_U519_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U520 (
    .in(in[3]),
    .clk(clk),
    .out(_U520_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U521 (
    .in(in[4]),
    .clk(clk),
    .out(_U521_out)
);
assign out[4] = _U521_out;
assign out[3] = _U520_out;
assign out[2] = _U519_out;
assign out[1] = _U518_out;
assign out[0] = _U517_out;
endmodule

module array_delay_U509 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U510_out;
wire [15:0] _U511_out;
wire [15:0] _U512_out;
wire [15:0] _U513_out;
wire [15:0] _U514_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U510 (
    .in(in[0]),
    .clk(clk),
    .out(_U510_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U511 (
    .in(in[1]),
    .clk(clk),
    .out(_U511_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U512 (
    .in(in[2]),
    .clk(clk),
    .out(_U512_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U513 (
    .in(in[3]),
    .clk(clk),
    .out(_U513_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U514 (
    .in(in[4]),
    .clk(clk),
    .out(_U514_out)
);
assign out[4] = _U514_out;
assign out[3] = _U513_out;
assign out[2] = _U512_out;
assign out[1] = _U511_out;
assign out[0] = _U510_out;
endmodule

module array_delay_U502 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U503_out;
wire [15:0] _U504_out;
wire [15:0] _U505_out;
wire [15:0] _U506_out;
wire [15:0] _U507_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U503 (
    .in(in[0]),
    .clk(clk),
    .out(_U503_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U504 (
    .in(in[1]),
    .clk(clk),
    .out(_U504_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U505 (
    .in(in[2]),
    .clk(clk),
    .out(_U505_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U506 (
    .in(in[3]),
    .clk(clk),
    .out(_U506_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U507 (
    .in(in[4]),
    .clk(clk),
    .out(_U507_out)
);
assign out[4] = _U507_out;
assign out[3] = _U506_out;
assign out[2] = _U505_out;
assign out[1] = _U504_out;
assign out[0] = _U503_out;
endmodule

module array_delay_U495 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U496_out;
wire [15:0] _U497_out;
wire [15:0] _U498_out;
wire [15:0] _U499_out;
wire [15:0] _U500_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U496 (
    .in(in[0]),
    .clk(clk),
    .out(_U496_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U497 (
    .in(in[1]),
    .clk(clk),
    .out(_U497_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U498 (
    .in(in[2]),
    .clk(clk),
    .out(_U498_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U499 (
    .in(in[3]),
    .clk(clk),
    .out(_U499_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U500 (
    .in(in[4]),
    .clk(clk),
    .out(_U500_out)
);
assign out[4] = _U500_out;
assign out[3] = _U499_out;
assign out[2] = _U498_out;
assign out[1] = _U497_out;
assign out[0] = _U496_out;
endmodule

module array_delay_U488 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U489_out;
wire [15:0] _U490_out;
wire [15:0] _U491_out;
wire [15:0] _U492_out;
wire [15:0] _U493_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U489 (
    .in(in[0]),
    .clk(clk),
    .out(_U489_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U490 (
    .in(in[1]),
    .clk(clk),
    .out(_U490_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U491 (
    .in(in[2]),
    .clk(clk),
    .out(_U491_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U492 (
    .in(in[3]),
    .clk(clk),
    .out(_U492_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U493 (
    .in(in[4]),
    .clk(clk),
    .out(_U493_out)
);
assign out[4] = _U493_out;
assign out[3] = _U492_out;
assign out[2] = _U491_out;
assign out[1] = _U490_out;
assign out[0] = _U489_out;
endmodule

module array_delay_U481 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U482_out;
wire [15:0] _U483_out;
wire [15:0] _U484_out;
wire [15:0] _U485_out;
wire [15:0] _U486_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U482 (
    .in(in[0]),
    .clk(clk),
    .out(_U482_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U483 (
    .in(in[1]),
    .clk(clk),
    .out(_U483_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U484 (
    .in(in[2]),
    .clk(clk),
    .out(_U484_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U485 (
    .in(in[3]),
    .clk(clk),
    .out(_U485_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U486 (
    .in(in[4]),
    .clk(clk),
    .out(_U486_out)
);
assign out[4] = _U486_out;
assign out[3] = _U485_out;
assign out[2] = _U484_out;
assign out[1] = _U483_out;
assign out[0] = _U482_out;
endmodule

module array_delay_U474 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U475_out;
wire [15:0] _U476_out;
wire [15:0] _U477_out;
wire [15:0] _U478_out;
wire [15:0] _U479_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U475 (
    .in(in[0]),
    .clk(clk),
    .out(_U475_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U476 (
    .in(in[1]),
    .clk(clk),
    .out(_U476_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U477 (
    .in(in[2]),
    .clk(clk),
    .out(_U477_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U478 (
    .in(in[3]),
    .clk(clk),
    .out(_U478_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U479 (
    .in(in[4]),
    .clk(clk),
    .out(_U479_out)
);
assign out[4] = _U479_out;
assign out[3] = _U478_out;
assign out[2] = _U477_out;
assign out[1] = _U476_out;
assign out[0] = _U475_out;
endmodule

module array_delay_U448 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U449_out;
wire [15:0] _U450_out;
wire [15:0] _U451_out;
wire [15:0] _U452_out;
wire [15:0] _U453_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U449 (
    .in(in[0]),
    .clk(clk),
    .out(_U449_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U450 (
    .in(in[1]),
    .clk(clk),
    .out(_U450_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U451 (
    .in(in[2]),
    .clk(clk),
    .out(_U451_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U452 (
    .in(in[3]),
    .clk(clk),
    .out(_U452_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U453 (
    .in(in[4]),
    .clk(clk),
    .out(_U453_out)
);
assign out[4] = _U453_out;
assign out[3] = _U452_out;
assign out[2] = _U451_out;
assign out[1] = _U450_out;
assign out[0] = _U449_out;
endmodule

module array_delay_U441 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U442_out;
wire [15:0] _U443_out;
wire [15:0] _U444_out;
wire [15:0] _U445_out;
wire [15:0] _U446_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U442 (
    .in(in[0]),
    .clk(clk),
    .out(_U442_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U443 (
    .in(in[1]),
    .clk(clk),
    .out(_U443_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U444 (
    .in(in[2]),
    .clk(clk),
    .out(_U444_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U445 (
    .in(in[3]),
    .clk(clk),
    .out(_U445_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U446 (
    .in(in[4]),
    .clk(clk),
    .out(_U446_out)
);
assign out[4] = _U446_out;
assign out[3] = _U445_out;
assign out[2] = _U444_out;
assign out[1] = _U443_out;
assign out[0] = _U442_out;
endmodule

module array_delay_U2280 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2281_out;
wire [15:0] _U2282_out;
wire [15:0] _U2283_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2281 (
    .in(in[0]),
    .clk(clk),
    .out(_U2281_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2282 (
    .in(in[1]),
    .clk(clk),
    .out(_U2282_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2283 (
    .in(in[2]),
    .clk(clk),
    .out(_U2283_out)
);
assign out[2] = _U2283_out;
assign out[1] = _U2282_out;
assign out[0] = _U2281_out;
endmodule

module array_delay_U2275 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2276_out;
wire [15:0] _U2277_out;
wire [15:0] _U2278_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2276 (
    .in(in[0]),
    .clk(clk),
    .out(_U2276_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2277 (
    .in(in[1]),
    .clk(clk),
    .out(_U2277_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2278 (
    .in(in[2]),
    .clk(clk),
    .out(_U2278_out)
);
assign out[2] = _U2278_out;
assign out[1] = _U2277_out;
assign out[0] = _U2276_out;
endmodule

module array_delay_U2266 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2267_out;
wire [15:0] _U2268_out;
wire [15:0] _U2269_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2267 (
    .in(in[0]),
    .clk(clk),
    .out(_U2267_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2268 (
    .in(in[1]),
    .clk(clk),
    .out(_U2268_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2269 (
    .in(in[2]),
    .clk(clk),
    .out(_U2269_out)
);
assign out[2] = _U2269_out;
assign out[1] = _U2268_out;
assign out[0] = _U2267_out;
endmodule

module array_delay_U2261 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2262_out;
wire [15:0] _U2263_out;
wire [15:0] _U2264_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2262 (
    .in(in[0]),
    .clk(clk),
    .out(_U2262_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2263 (
    .in(in[1]),
    .clk(clk),
    .out(_U2263_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2264 (
    .in(in[2]),
    .clk(clk),
    .out(_U2264_out)
);
assign out[2] = _U2264_out;
assign out[1] = _U2263_out;
assign out[0] = _U2262_out;
endmodule

module array_delay_U2233 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2234_out;
wire [15:0] _U2235_out;
wire [15:0] _U2236_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2234 (
    .in(in[0]),
    .clk(clk),
    .out(_U2234_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2235 (
    .in(in[1]),
    .clk(clk),
    .out(_U2235_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2236 (
    .in(in[2]),
    .clk(clk),
    .out(_U2236_out)
);
assign out[2] = _U2236_out;
assign out[1] = _U2235_out;
assign out[0] = _U2234_out;
endmodule

module array_delay_U2228 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2229_out;
wire [15:0] _U2230_out;
wire [15:0] _U2231_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2229 (
    .in(in[0]),
    .clk(clk),
    .out(_U2229_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2230 (
    .in(in[1]),
    .clk(clk),
    .out(_U2230_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2231 (
    .in(in[2]),
    .clk(clk),
    .out(_U2231_out)
);
assign out[2] = _U2231_out;
assign out[1] = _U2230_out;
assign out[0] = _U2229_out;
endmodule

module array_delay_U2219 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2220_out;
wire [15:0] _U2221_out;
wire [15:0] _U2222_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2220 (
    .in(in[0]),
    .clk(clk),
    .out(_U2220_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2221 (
    .in(in[1]),
    .clk(clk),
    .out(_U2221_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2222 (
    .in(in[2]),
    .clk(clk),
    .out(_U2222_out)
);
assign out[2] = _U2222_out;
assign out[1] = _U2221_out;
assign out[0] = _U2220_out;
endmodule

module array_delay_U2214 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2215_out;
wire [15:0] _U2216_out;
wire [15:0] _U2217_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2215 (
    .in(in[0]),
    .clk(clk),
    .out(_U2215_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2216 (
    .in(in[1]),
    .clk(clk),
    .out(_U2216_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2217 (
    .in(in[2]),
    .clk(clk),
    .out(_U2217_out)
);
assign out[2] = _U2217_out;
assign out[1] = _U2216_out;
assign out[0] = _U2215_out;
endmodule

module array_delay_U2186 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2187_out;
wire [15:0] _U2188_out;
wire [15:0] _U2189_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2187 (
    .in(in[0]),
    .clk(clk),
    .out(_U2187_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2188 (
    .in(in[1]),
    .clk(clk),
    .out(_U2188_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2189 (
    .in(in[2]),
    .clk(clk),
    .out(_U2189_out)
);
assign out[2] = _U2189_out;
assign out[1] = _U2188_out;
assign out[0] = _U2187_out;
endmodule

module array_delay_U2181 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2182_out;
wire [15:0] _U2183_out;
wire [15:0] _U2184_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2182 (
    .in(in[0]),
    .clk(clk),
    .out(_U2182_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2183 (
    .in(in[1]),
    .clk(clk),
    .out(_U2183_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2184 (
    .in(in[2]),
    .clk(clk),
    .out(_U2184_out)
);
assign out[2] = _U2184_out;
assign out[1] = _U2183_out;
assign out[0] = _U2182_out;
endmodule

module array_delay_U2172 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2173_out;
wire [15:0] _U2174_out;
wire [15:0] _U2175_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2173 (
    .in(in[0]),
    .clk(clk),
    .out(_U2173_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2174 (
    .in(in[1]),
    .clk(clk),
    .out(_U2174_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2175 (
    .in(in[2]),
    .clk(clk),
    .out(_U2175_out)
);
assign out[2] = _U2175_out;
assign out[1] = _U2174_out;
assign out[0] = _U2173_out;
endmodule

module array_delay_U2167 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2168_out;
wire [15:0] _U2169_out;
wire [15:0] _U2170_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2168 (
    .in(in[0]),
    .clk(clk),
    .out(_U2168_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2169 (
    .in(in[1]),
    .clk(clk),
    .out(_U2169_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2170 (
    .in(in[2]),
    .clk(clk),
    .out(_U2170_out)
);
assign out[2] = _U2170_out;
assign out[1] = _U2169_out;
assign out[0] = _U2168_out;
endmodule

module array_delay_U2139 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2140_out;
wire [15:0] _U2141_out;
wire [15:0] _U2142_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2140 (
    .in(in[0]),
    .clk(clk),
    .out(_U2140_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2141 (
    .in(in[1]),
    .clk(clk),
    .out(_U2141_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2142 (
    .in(in[2]),
    .clk(clk),
    .out(_U2142_out)
);
assign out[2] = _U2142_out;
assign out[1] = _U2141_out;
assign out[0] = _U2140_out;
endmodule

module array_delay_U2134 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2135_out;
wire [15:0] _U2136_out;
wire [15:0] _U2137_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2135 (
    .in(in[0]),
    .clk(clk),
    .out(_U2135_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2136 (
    .in(in[1]),
    .clk(clk),
    .out(_U2136_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2137 (
    .in(in[2]),
    .clk(clk),
    .out(_U2137_out)
);
assign out[2] = _U2137_out;
assign out[1] = _U2136_out;
assign out[0] = _U2135_out;
endmodule

module array_delay_U2125 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2126_out;
wire [15:0] _U2127_out;
wire [15:0] _U2128_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2126 (
    .in(in[0]),
    .clk(clk),
    .out(_U2126_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2127 (
    .in(in[1]),
    .clk(clk),
    .out(_U2127_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2128 (
    .in(in[2]),
    .clk(clk),
    .out(_U2128_out)
);
assign out[2] = _U2128_out;
assign out[1] = _U2127_out;
assign out[0] = _U2126_out;
endmodule

module array_delay_U2120 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2121_out;
wire [15:0] _U2122_out;
wire [15:0] _U2123_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2121 (
    .in(in[0]),
    .clk(clk),
    .out(_U2121_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2122 (
    .in(in[1]),
    .clk(clk),
    .out(_U2122_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2123 (
    .in(in[2]),
    .clk(clk),
    .out(_U2123_out)
);
assign out[2] = _U2123_out;
assign out[1] = _U2122_out;
assign out[0] = _U2121_out;
endmodule

module array_delay_U2092 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2093_out;
wire [15:0] _U2094_out;
wire [15:0] _U2095_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2093 (
    .in(in[0]),
    .clk(clk),
    .out(_U2093_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2094 (
    .in(in[1]),
    .clk(clk),
    .out(_U2094_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2095 (
    .in(in[2]),
    .clk(clk),
    .out(_U2095_out)
);
assign out[2] = _U2095_out;
assign out[1] = _U2094_out;
assign out[0] = _U2093_out;
endmodule

module array_delay_U2087 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2088_out;
wire [15:0] _U2089_out;
wire [15:0] _U2090_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2088 (
    .in(in[0]),
    .clk(clk),
    .out(_U2088_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2089 (
    .in(in[1]),
    .clk(clk),
    .out(_U2089_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2090 (
    .in(in[2]),
    .clk(clk),
    .out(_U2090_out)
);
assign out[2] = _U2090_out;
assign out[1] = _U2089_out;
assign out[0] = _U2088_out;
endmodule

module array_delay_U2078 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2079_out;
wire [15:0] _U2080_out;
wire [15:0] _U2081_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2079 (
    .in(in[0]),
    .clk(clk),
    .out(_U2079_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2080 (
    .in(in[1]),
    .clk(clk),
    .out(_U2080_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2081 (
    .in(in[2]),
    .clk(clk),
    .out(_U2081_out)
);
assign out[2] = _U2081_out;
assign out[1] = _U2080_out;
assign out[0] = _U2079_out;
endmodule

module array_delay_U2073 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2074_out;
wire [15:0] _U2075_out;
wire [15:0] _U2076_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2074 (
    .in(in[0]),
    .clk(clk),
    .out(_U2074_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2075 (
    .in(in[1]),
    .clk(clk),
    .out(_U2075_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2076 (
    .in(in[2]),
    .clk(clk),
    .out(_U2076_out)
);
assign out[2] = _U2076_out;
assign out[1] = _U2075_out;
assign out[0] = _U2074_out;
endmodule

module array_delay_U2045 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2046_out;
wire [15:0] _U2047_out;
wire [15:0] _U2048_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2046 (
    .in(in[0]),
    .clk(clk),
    .out(_U2046_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2047 (
    .in(in[1]),
    .clk(clk),
    .out(_U2047_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2048 (
    .in(in[2]),
    .clk(clk),
    .out(_U2048_out)
);
assign out[2] = _U2048_out;
assign out[1] = _U2047_out;
assign out[0] = _U2046_out;
endmodule

module array_delay_U2040 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2041_out;
wire [15:0] _U2042_out;
wire [15:0] _U2043_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2041 (
    .in(in[0]),
    .clk(clk),
    .out(_U2041_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2042 (
    .in(in[1]),
    .clk(clk),
    .out(_U2042_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2043 (
    .in(in[2]),
    .clk(clk),
    .out(_U2043_out)
);
assign out[2] = _U2043_out;
assign out[1] = _U2042_out;
assign out[0] = _U2041_out;
endmodule

module array_delay_U2031 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2032_out;
wire [15:0] _U2033_out;
wire [15:0] _U2034_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2032 (
    .in(in[0]),
    .clk(clk),
    .out(_U2032_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2033 (
    .in(in[1]),
    .clk(clk),
    .out(_U2033_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2034 (
    .in(in[2]),
    .clk(clk),
    .out(_U2034_out)
);
assign out[2] = _U2034_out;
assign out[1] = _U2033_out;
assign out[0] = _U2032_out;
endmodule

module array_delay_U2026 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2027_out;
wire [15:0] _U2028_out;
wire [15:0] _U2029_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2027 (
    .in(in[0]),
    .clk(clk),
    .out(_U2027_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2028 (
    .in(in[1]),
    .clk(clk),
    .out(_U2028_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2029 (
    .in(in[2]),
    .clk(clk),
    .out(_U2029_out)
);
assign out[2] = _U2029_out;
assign out[1] = _U2028_out;
assign out[0] = _U2027_out;
endmodule

module array_delay_U1998 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1999_out;
wire [15:0] _U2000_out;
wire [15:0] _U2001_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1999 (
    .in(in[0]),
    .clk(clk),
    .out(_U1999_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2000 (
    .in(in[1]),
    .clk(clk),
    .out(_U2000_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2001 (
    .in(in[2]),
    .clk(clk),
    .out(_U2001_out)
);
assign out[2] = _U2001_out;
assign out[1] = _U2000_out;
assign out[0] = _U1999_out;
endmodule

module array_delay_U1993 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1994_out;
wire [15:0] _U1995_out;
wire [15:0] _U1996_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1994 (
    .in(in[0]),
    .clk(clk),
    .out(_U1994_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1995 (
    .in(in[1]),
    .clk(clk),
    .out(_U1995_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1996 (
    .in(in[2]),
    .clk(clk),
    .out(_U1996_out)
);
assign out[2] = _U1996_out;
assign out[1] = _U1995_out;
assign out[0] = _U1994_out;
endmodule

module array_delay_U1984 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1985_out;
wire [15:0] _U1986_out;
wire [15:0] _U1987_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1985 (
    .in(in[0]),
    .clk(clk),
    .out(_U1985_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1986 (
    .in(in[1]),
    .clk(clk),
    .out(_U1986_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1987 (
    .in(in[2]),
    .clk(clk),
    .out(_U1987_out)
);
assign out[2] = _U1987_out;
assign out[1] = _U1986_out;
assign out[0] = _U1985_out;
endmodule

module array_delay_U1979 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1980_out;
wire [15:0] _U1981_out;
wire [15:0] _U1982_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1980 (
    .in(in[0]),
    .clk(clk),
    .out(_U1980_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1981 (
    .in(in[1]),
    .clk(clk),
    .out(_U1981_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1982 (
    .in(in[2]),
    .clk(clk),
    .out(_U1982_out)
);
assign out[2] = _U1982_out;
assign out[1] = _U1981_out;
assign out[0] = _U1980_out;
endmodule

module array_delay_U1951 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1952_out;
wire [15:0] _U1953_out;
wire [15:0] _U1954_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1952 (
    .in(in[0]),
    .clk(clk),
    .out(_U1952_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1953 (
    .in(in[1]),
    .clk(clk),
    .out(_U1953_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1954 (
    .in(in[2]),
    .clk(clk),
    .out(_U1954_out)
);
assign out[2] = _U1954_out;
assign out[1] = _U1953_out;
assign out[0] = _U1952_out;
endmodule

module array_delay_U1946 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1947_out;
wire [15:0] _U1948_out;
wire [15:0] _U1949_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1947 (
    .in(in[0]),
    .clk(clk),
    .out(_U1947_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1948 (
    .in(in[1]),
    .clk(clk),
    .out(_U1948_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1949 (
    .in(in[2]),
    .clk(clk),
    .out(_U1949_out)
);
assign out[2] = _U1949_out;
assign out[1] = _U1948_out;
assign out[0] = _U1947_out;
endmodule

module array_delay_U1937 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1938_out;
wire [15:0] _U1939_out;
wire [15:0] _U1940_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1938 (
    .in(in[0]),
    .clk(clk),
    .out(_U1938_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1939 (
    .in(in[1]),
    .clk(clk),
    .out(_U1939_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1940 (
    .in(in[2]),
    .clk(clk),
    .out(_U1940_out)
);
assign out[2] = _U1940_out;
assign out[1] = _U1939_out;
assign out[0] = _U1938_out;
endmodule

module array_delay_U1932 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1933_out;
wire [15:0] _U1934_out;
wire [15:0] _U1935_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1933 (
    .in(in[0]),
    .clk(clk),
    .out(_U1933_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1934 (
    .in(in[1]),
    .clk(clk),
    .out(_U1934_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1935 (
    .in(in[2]),
    .clk(clk),
    .out(_U1935_out)
);
assign out[2] = _U1935_out;
assign out[1] = _U1934_out;
assign out[0] = _U1933_out;
endmodule

module array_delay_U1902 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1903_out;
wire [15:0] _U1904_out;
wire [15:0] _U1905_out;
wire [15:0] _U1906_out;
wire [15:0] _U1907_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1903 (
    .in(in[0]),
    .clk(clk),
    .out(_U1903_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1904 (
    .in(in[1]),
    .clk(clk),
    .out(_U1904_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1905 (
    .in(in[2]),
    .clk(clk),
    .out(_U1905_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1906 (
    .in(in[3]),
    .clk(clk),
    .out(_U1906_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1907 (
    .in(in[4]),
    .clk(clk),
    .out(_U1907_out)
);
assign out[4] = _U1907_out;
assign out[3] = _U1906_out;
assign out[2] = _U1905_out;
assign out[1] = _U1904_out;
assign out[0] = _U1903_out;
endmodule

module array_delay_U1895 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1896_out;
wire [15:0] _U1897_out;
wire [15:0] _U1898_out;
wire [15:0] _U1899_out;
wire [15:0] _U1900_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1896 (
    .in(in[0]),
    .clk(clk),
    .out(_U1896_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1897 (
    .in(in[1]),
    .clk(clk),
    .out(_U1897_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1898 (
    .in(in[2]),
    .clk(clk),
    .out(_U1898_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1899 (
    .in(in[3]),
    .clk(clk),
    .out(_U1899_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1900 (
    .in(in[4]),
    .clk(clk),
    .out(_U1900_out)
);
assign out[4] = _U1900_out;
assign out[3] = _U1899_out;
assign out[2] = _U1898_out;
assign out[1] = _U1897_out;
assign out[0] = _U1896_out;
endmodule

module array_delay_U1888 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1889_out;
wire [15:0] _U1890_out;
wire [15:0] _U1891_out;
wire [15:0] _U1892_out;
wire [15:0] _U1893_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1889 (
    .in(in[0]),
    .clk(clk),
    .out(_U1889_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1890 (
    .in(in[1]),
    .clk(clk),
    .out(_U1890_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1891 (
    .in(in[2]),
    .clk(clk),
    .out(_U1891_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1892 (
    .in(in[3]),
    .clk(clk),
    .out(_U1892_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1893 (
    .in(in[4]),
    .clk(clk),
    .out(_U1893_out)
);
assign out[4] = _U1893_out;
assign out[3] = _U1892_out;
assign out[2] = _U1891_out;
assign out[1] = _U1890_out;
assign out[0] = _U1889_out;
endmodule

module array_delay_U1881 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1882_out;
wire [15:0] _U1883_out;
wire [15:0] _U1884_out;
wire [15:0] _U1885_out;
wire [15:0] _U1886_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1882 (
    .in(in[0]),
    .clk(clk),
    .out(_U1882_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1883 (
    .in(in[1]),
    .clk(clk),
    .out(_U1883_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1884 (
    .in(in[2]),
    .clk(clk),
    .out(_U1884_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1885 (
    .in(in[3]),
    .clk(clk),
    .out(_U1885_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1886 (
    .in(in[4]),
    .clk(clk),
    .out(_U1886_out)
);
assign out[4] = _U1886_out;
assign out[3] = _U1885_out;
assign out[2] = _U1884_out;
assign out[1] = _U1883_out;
assign out[0] = _U1882_out;
endmodule

module array_delay_U1874 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1875_out;
wire [15:0] _U1876_out;
wire [15:0] _U1877_out;
wire [15:0] _U1878_out;
wire [15:0] _U1879_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1875 (
    .in(in[0]),
    .clk(clk),
    .out(_U1875_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1876 (
    .in(in[1]),
    .clk(clk),
    .out(_U1876_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1877 (
    .in(in[2]),
    .clk(clk),
    .out(_U1877_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1878 (
    .in(in[3]),
    .clk(clk),
    .out(_U1878_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1879 (
    .in(in[4]),
    .clk(clk),
    .out(_U1879_out)
);
assign out[4] = _U1879_out;
assign out[3] = _U1878_out;
assign out[2] = _U1877_out;
assign out[1] = _U1876_out;
assign out[0] = _U1875_out;
endmodule

module array_delay_U1867 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1868_out;
wire [15:0] _U1869_out;
wire [15:0] _U1870_out;
wire [15:0] _U1871_out;
wire [15:0] _U1872_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1868 (
    .in(in[0]),
    .clk(clk),
    .out(_U1868_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1869 (
    .in(in[1]),
    .clk(clk),
    .out(_U1869_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1870 (
    .in(in[2]),
    .clk(clk),
    .out(_U1870_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1871 (
    .in(in[3]),
    .clk(clk),
    .out(_U1871_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1872 (
    .in(in[4]),
    .clk(clk),
    .out(_U1872_out)
);
assign out[4] = _U1872_out;
assign out[3] = _U1871_out;
assign out[2] = _U1870_out;
assign out[1] = _U1869_out;
assign out[0] = _U1868_out;
endmodule

module array_delay_U1860 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1861_out;
wire [15:0] _U1862_out;
wire [15:0] _U1863_out;
wire [15:0] _U1864_out;
wire [15:0] _U1865_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1861 (
    .in(in[0]),
    .clk(clk),
    .out(_U1861_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1862 (
    .in(in[1]),
    .clk(clk),
    .out(_U1862_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1863 (
    .in(in[2]),
    .clk(clk),
    .out(_U1863_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1864 (
    .in(in[3]),
    .clk(clk),
    .out(_U1864_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1865 (
    .in(in[4]),
    .clk(clk),
    .out(_U1865_out)
);
assign out[4] = _U1865_out;
assign out[3] = _U1864_out;
assign out[2] = _U1863_out;
assign out[1] = _U1862_out;
assign out[0] = _U1861_out;
endmodule

module array_delay_U1853 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1854_out;
wire [15:0] _U1855_out;
wire [15:0] _U1856_out;
wire [15:0] _U1857_out;
wire [15:0] _U1858_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1854 (
    .in(in[0]),
    .clk(clk),
    .out(_U1854_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1855 (
    .in(in[1]),
    .clk(clk),
    .out(_U1855_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1856 (
    .in(in[2]),
    .clk(clk),
    .out(_U1856_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1857 (
    .in(in[3]),
    .clk(clk),
    .out(_U1857_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1858 (
    .in(in[4]),
    .clk(clk),
    .out(_U1858_out)
);
assign out[4] = _U1858_out;
assign out[3] = _U1857_out;
assign out[2] = _U1856_out;
assign out[1] = _U1855_out;
assign out[0] = _U1854_out;
endmodule

module array_delay_U1846 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1847_out;
wire [15:0] _U1848_out;
wire [15:0] _U1849_out;
wire [15:0] _U1850_out;
wire [15:0] _U1851_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1847 (
    .in(in[0]),
    .clk(clk),
    .out(_U1847_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1848 (
    .in(in[1]),
    .clk(clk),
    .out(_U1848_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1849 (
    .in(in[2]),
    .clk(clk),
    .out(_U1849_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1850 (
    .in(in[3]),
    .clk(clk),
    .out(_U1850_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1851 (
    .in(in[4]),
    .clk(clk),
    .out(_U1851_out)
);
assign out[4] = _U1851_out;
assign out[3] = _U1850_out;
assign out[2] = _U1849_out;
assign out[1] = _U1848_out;
assign out[0] = _U1847_out;
endmodule

module array_delay_U1839 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1840_out;
wire [15:0] _U1841_out;
wire [15:0] _U1842_out;
wire [15:0] _U1843_out;
wire [15:0] _U1844_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1840 (
    .in(in[0]),
    .clk(clk),
    .out(_U1840_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1841 (
    .in(in[1]),
    .clk(clk),
    .out(_U1841_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1842 (
    .in(in[2]),
    .clk(clk),
    .out(_U1842_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1843 (
    .in(in[3]),
    .clk(clk),
    .out(_U1843_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1844 (
    .in(in[4]),
    .clk(clk),
    .out(_U1844_out)
);
assign out[4] = _U1844_out;
assign out[3] = _U1843_out;
assign out[2] = _U1842_out;
assign out[1] = _U1841_out;
assign out[0] = _U1840_out;
endmodule

module array_delay_U1832 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1833_out;
wire [15:0] _U1834_out;
wire [15:0] _U1835_out;
wire [15:0] _U1836_out;
wire [15:0] _U1837_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1833 (
    .in(in[0]),
    .clk(clk),
    .out(_U1833_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1834 (
    .in(in[1]),
    .clk(clk),
    .out(_U1834_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1835 (
    .in(in[2]),
    .clk(clk),
    .out(_U1835_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1836 (
    .in(in[3]),
    .clk(clk),
    .out(_U1836_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1837 (
    .in(in[4]),
    .clk(clk),
    .out(_U1837_out)
);
assign out[4] = _U1837_out;
assign out[3] = _U1836_out;
assign out[2] = _U1835_out;
assign out[1] = _U1834_out;
assign out[0] = _U1833_out;
endmodule

module array_delay_U1825 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1826_out;
wire [15:0] _U1827_out;
wire [15:0] _U1828_out;
wire [15:0] _U1829_out;
wire [15:0] _U1830_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1826 (
    .in(in[0]),
    .clk(clk),
    .out(_U1826_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1827 (
    .in(in[1]),
    .clk(clk),
    .out(_U1827_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1828 (
    .in(in[2]),
    .clk(clk),
    .out(_U1828_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1829 (
    .in(in[3]),
    .clk(clk),
    .out(_U1829_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1830 (
    .in(in[4]),
    .clk(clk),
    .out(_U1830_out)
);
assign out[4] = _U1830_out;
assign out[3] = _U1829_out;
assign out[2] = _U1828_out;
assign out[1] = _U1827_out;
assign out[0] = _U1826_out;
endmodule

module array_delay_U1818 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1819_out;
wire [15:0] _U1820_out;
wire [15:0] _U1821_out;
wire [15:0] _U1822_out;
wire [15:0] _U1823_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1819 (
    .in(in[0]),
    .clk(clk),
    .out(_U1819_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1820 (
    .in(in[1]),
    .clk(clk),
    .out(_U1820_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1821 (
    .in(in[2]),
    .clk(clk),
    .out(_U1821_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1822 (
    .in(in[3]),
    .clk(clk),
    .out(_U1822_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1823 (
    .in(in[4]),
    .clk(clk),
    .out(_U1823_out)
);
assign out[4] = _U1823_out;
assign out[3] = _U1822_out;
assign out[2] = _U1821_out;
assign out[1] = _U1820_out;
assign out[0] = _U1819_out;
endmodule

module array_delay_U1811 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1812_out;
wire [15:0] _U1813_out;
wire [15:0] _U1814_out;
wire [15:0] _U1815_out;
wire [15:0] _U1816_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1812 (
    .in(in[0]),
    .clk(clk),
    .out(_U1812_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1813 (
    .in(in[1]),
    .clk(clk),
    .out(_U1813_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1814 (
    .in(in[2]),
    .clk(clk),
    .out(_U1814_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1815 (
    .in(in[3]),
    .clk(clk),
    .out(_U1815_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1816 (
    .in(in[4]),
    .clk(clk),
    .out(_U1816_out)
);
assign out[4] = _U1816_out;
assign out[3] = _U1815_out;
assign out[2] = _U1814_out;
assign out[1] = _U1813_out;
assign out[0] = _U1812_out;
endmodule

module array_delay_U1804 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1805_out;
wire [15:0] _U1806_out;
wire [15:0] _U1807_out;
wire [15:0] _U1808_out;
wire [15:0] _U1809_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1805 (
    .in(in[0]),
    .clk(clk),
    .out(_U1805_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1806 (
    .in(in[1]),
    .clk(clk),
    .out(_U1806_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1807 (
    .in(in[2]),
    .clk(clk),
    .out(_U1807_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1808 (
    .in(in[3]),
    .clk(clk),
    .out(_U1808_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1809 (
    .in(in[4]),
    .clk(clk),
    .out(_U1809_out)
);
assign out[4] = _U1809_out;
assign out[3] = _U1808_out;
assign out[2] = _U1807_out;
assign out[1] = _U1806_out;
assign out[0] = _U1805_out;
endmodule

module array_delay_U1797 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1798_out;
wire [15:0] _U1799_out;
wire [15:0] _U1800_out;
wire [15:0] _U1801_out;
wire [15:0] _U1802_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1798 (
    .in(in[0]),
    .clk(clk),
    .out(_U1798_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1799 (
    .in(in[1]),
    .clk(clk),
    .out(_U1799_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1800 (
    .in(in[2]),
    .clk(clk),
    .out(_U1800_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1801 (
    .in(in[3]),
    .clk(clk),
    .out(_U1801_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1802 (
    .in(in[4]),
    .clk(clk),
    .out(_U1802_out)
);
assign out[4] = _U1802_out;
assign out[3] = _U1801_out;
assign out[2] = _U1800_out;
assign out[1] = _U1799_out;
assign out[0] = _U1798_out;
endmodule

module array_delay_U1790 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1791_out;
wire [15:0] _U1792_out;
wire [15:0] _U1793_out;
wire [15:0] _U1794_out;
wire [15:0] _U1795_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1791 (
    .in(in[0]),
    .clk(clk),
    .out(_U1791_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1792 (
    .in(in[1]),
    .clk(clk),
    .out(_U1792_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1793 (
    .in(in[2]),
    .clk(clk),
    .out(_U1793_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1794 (
    .in(in[3]),
    .clk(clk),
    .out(_U1794_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1795 (
    .in(in[4]),
    .clk(clk),
    .out(_U1795_out)
);
assign out[4] = _U1795_out;
assign out[3] = _U1794_out;
assign out[2] = _U1793_out;
assign out[1] = _U1792_out;
assign out[0] = _U1791_out;
endmodule

module array_delay_U1764 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1765_out;
wire [15:0] _U1766_out;
wire [15:0] _U1767_out;
wire [15:0] _U1768_out;
wire [15:0] _U1769_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1765 (
    .in(in[0]),
    .clk(clk),
    .out(_U1765_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1766 (
    .in(in[1]),
    .clk(clk),
    .out(_U1766_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1767 (
    .in(in[2]),
    .clk(clk),
    .out(_U1767_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1768 (
    .in(in[3]),
    .clk(clk),
    .out(_U1768_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1769 (
    .in(in[4]),
    .clk(clk),
    .out(_U1769_out)
);
assign out[4] = _U1769_out;
assign out[3] = _U1768_out;
assign out[2] = _U1767_out;
assign out[1] = _U1766_out;
assign out[0] = _U1765_out;
endmodule

module array_delay_U1757 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1758_out;
wire [15:0] _U1759_out;
wire [15:0] _U1760_out;
wire [15:0] _U1761_out;
wire [15:0] _U1762_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1758 (
    .in(in[0]),
    .clk(clk),
    .out(_U1758_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1759 (
    .in(in[1]),
    .clk(clk),
    .out(_U1759_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1760 (
    .in(in[2]),
    .clk(clk),
    .out(_U1760_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1761 (
    .in(in[3]),
    .clk(clk),
    .out(_U1761_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1762 (
    .in(in[4]),
    .clk(clk),
    .out(_U1762_out)
);
assign out[4] = _U1762_out;
assign out[3] = _U1761_out;
assign out[2] = _U1760_out;
assign out[1] = _U1759_out;
assign out[0] = _U1758_out;
endmodule

module array_delay_U1714 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1715_out;
wire [15:0] _U1716_out;
wire [15:0] _U1717_out;
wire [15:0] _U1718_out;
wire [15:0] _U1719_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1715 (
    .in(in[0]),
    .clk(clk),
    .out(_U1715_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1716 (
    .in(in[1]),
    .clk(clk),
    .out(_U1716_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1717 (
    .in(in[2]),
    .clk(clk),
    .out(_U1717_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1718 (
    .in(in[3]),
    .clk(clk),
    .out(_U1718_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1719 (
    .in(in[4]),
    .clk(clk),
    .out(_U1719_out)
);
assign out[4] = _U1719_out;
assign out[3] = _U1718_out;
assign out[2] = _U1717_out;
assign out[1] = _U1716_out;
assign out[0] = _U1715_out;
endmodule

module array_delay_U1707 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1708_out;
wire [15:0] _U1709_out;
wire [15:0] _U1710_out;
wire [15:0] _U1711_out;
wire [15:0] _U1712_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1708 (
    .in(in[0]),
    .clk(clk),
    .out(_U1708_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1709 (
    .in(in[1]),
    .clk(clk),
    .out(_U1709_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1710 (
    .in(in[2]),
    .clk(clk),
    .out(_U1710_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1711 (
    .in(in[3]),
    .clk(clk),
    .out(_U1711_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1712 (
    .in(in[4]),
    .clk(clk),
    .out(_U1712_out)
);
assign out[4] = _U1712_out;
assign out[3] = _U1711_out;
assign out[2] = _U1710_out;
assign out[1] = _U1709_out;
assign out[0] = _U1708_out;
endmodule

module array_delay_U1700 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1701_out;
wire [15:0] _U1702_out;
wire [15:0] _U1703_out;
wire [15:0] _U1704_out;
wire [15:0] _U1705_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1701 (
    .in(in[0]),
    .clk(clk),
    .out(_U1701_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1702 (
    .in(in[1]),
    .clk(clk),
    .out(_U1702_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1703 (
    .in(in[2]),
    .clk(clk),
    .out(_U1703_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1704 (
    .in(in[3]),
    .clk(clk),
    .out(_U1704_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1705 (
    .in(in[4]),
    .clk(clk),
    .out(_U1705_out)
);
assign out[4] = _U1705_out;
assign out[3] = _U1704_out;
assign out[2] = _U1703_out;
assign out[1] = _U1702_out;
assign out[0] = _U1701_out;
endmodule

module array_delay_U1693 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1694_out;
wire [15:0] _U1695_out;
wire [15:0] _U1696_out;
wire [15:0] _U1697_out;
wire [15:0] _U1698_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1694 (
    .in(in[0]),
    .clk(clk),
    .out(_U1694_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1695 (
    .in(in[1]),
    .clk(clk),
    .out(_U1695_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1696 (
    .in(in[2]),
    .clk(clk),
    .out(_U1696_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1697 (
    .in(in[3]),
    .clk(clk),
    .out(_U1697_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1698 (
    .in(in[4]),
    .clk(clk),
    .out(_U1698_out)
);
assign out[4] = _U1698_out;
assign out[3] = _U1697_out;
assign out[2] = _U1696_out;
assign out[1] = _U1695_out;
assign out[0] = _U1694_out;
endmodule

module array_delay_U1686 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1687_out;
wire [15:0] _U1688_out;
wire [15:0] _U1689_out;
wire [15:0] _U1690_out;
wire [15:0] _U1691_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1687 (
    .in(in[0]),
    .clk(clk),
    .out(_U1687_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1688 (
    .in(in[1]),
    .clk(clk),
    .out(_U1688_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1689 (
    .in(in[2]),
    .clk(clk),
    .out(_U1689_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1690 (
    .in(in[3]),
    .clk(clk),
    .out(_U1690_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1691 (
    .in(in[4]),
    .clk(clk),
    .out(_U1691_out)
);
assign out[4] = _U1691_out;
assign out[3] = _U1690_out;
assign out[2] = _U1689_out;
assign out[1] = _U1688_out;
assign out[0] = _U1687_out;
endmodule

module array_delay_U1679 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1680_out;
wire [15:0] _U1681_out;
wire [15:0] _U1682_out;
wire [15:0] _U1683_out;
wire [15:0] _U1684_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1680 (
    .in(in[0]),
    .clk(clk),
    .out(_U1680_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1681 (
    .in(in[1]),
    .clk(clk),
    .out(_U1681_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1682 (
    .in(in[2]),
    .clk(clk),
    .out(_U1682_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1683 (
    .in(in[3]),
    .clk(clk),
    .out(_U1683_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1684 (
    .in(in[4]),
    .clk(clk),
    .out(_U1684_out)
);
assign out[4] = _U1684_out;
assign out[3] = _U1683_out;
assign out[2] = _U1682_out;
assign out[1] = _U1681_out;
assign out[0] = _U1680_out;
endmodule

module array_delay_U1672 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1673_out;
wire [15:0] _U1674_out;
wire [15:0] _U1675_out;
wire [15:0] _U1676_out;
wire [15:0] _U1677_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1673 (
    .in(in[0]),
    .clk(clk),
    .out(_U1673_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1674 (
    .in(in[1]),
    .clk(clk),
    .out(_U1674_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1675 (
    .in(in[2]),
    .clk(clk),
    .out(_U1675_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1676 (
    .in(in[3]),
    .clk(clk),
    .out(_U1676_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1677 (
    .in(in[4]),
    .clk(clk),
    .out(_U1677_out)
);
assign out[4] = _U1677_out;
assign out[3] = _U1676_out;
assign out[2] = _U1675_out;
assign out[1] = _U1674_out;
assign out[0] = _U1673_out;
endmodule

module array_delay_U1665 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1666_out;
wire [15:0] _U1667_out;
wire [15:0] _U1668_out;
wire [15:0] _U1669_out;
wire [15:0] _U1670_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1666 (
    .in(in[0]),
    .clk(clk),
    .out(_U1666_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1667 (
    .in(in[1]),
    .clk(clk),
    .out(_U1667_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1668 (
    .in(in[2]),
    .clk(clk),
    .out(_U1668_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1669 (
    .in(in[3]),
    .clk(clk),
    .out(_U1669_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1670 (
    .in(in[4]),
    .clk(clk),
    .out(_U1670_out)
);
assign out[4] = _U1670_out;
assign out[3] = _U1669_out;
assign out[2] = _U1668_out;
assign out[1] = _U1667_out;
assign out[0] = _U1666_out;
endmodule

module array_delay_U1658 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1659_out;
wire [15:0] _U1660_out;
wire [15:0] _U1661_out;
wire [15:0] _U1662_out;
wire [15:0] _U1663_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1659 (
    .in(in[0]),
    .clk(clk),
    .out(_U1659_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1660 (
    .in(in[1]),
    .clk(clk),
    .out(_U1660_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1661 (
    .in(in[2]),
    .clk(clk),
    .out(_U1661_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1662 (
    .in(in[3]),
    .clk(clk),
    .out(_U1662_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1663 (
    .in(in[4]),
    .clk(clk),
    .out(_U1663_out)
);
assign out[4] = _U1663_out;
assign out[3] = _U1662_out;
assign out[2] = _U1661_out;
assign out[1] = _U1660_out;
assign out[0] = _U1659_out;
endmodule

module array_delay_U1651 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1652_out;
wire [15:0] _U1653_out;
wire [15:0] _U1654_out;
wire [15:0] _U1655_out;
wire [15:0] _U1656_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1652 (
    .in(in[0]),
    .clk(clk),
    .out(_U1652_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1653 (
    .in(in[1]),
    .clk(clk),
    .out(_U1653_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1654 (
    .in(in[2]),
    .clk(clk),
    .out(_U1654_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1655 (
    .in(in[3]),
    .clk(clk),
    .out(_U1655_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1656 (
    .in(in[4]),
    .clk(clk),
    .out(_U1656_out)
);
assign out[4] = _U1656_out;
assign out[3] = _U1655_out;
assign out[2] = _U1654_out;
assign out[1] = _U1653_out;
assign out[0] = _U1652_out;
endmodule

module array_delay_U1644 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1645_out;
wire [15:0] _U1646_out;
wire [15:0] _U1647_out;
wire [15:0] _U1648_out;
wire [15:0] _U1649_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1645 (
    .in(in[0]),
    .clk(clk),
    .out(_U1645_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1646 (
    .in(in[1]),
    .clk(clk),
    .out(_U1646_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1647 (
    .in(in[2]),
    .clk(clk),
    .out(_U1647_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1648 (
    .in(in[3]),
    .clk(clk),
    .out(_U1648_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1649 (
    .in(in[4]),
    .clk(clk),
    .out(_U1649_out)
);
assign out[4] = _U1649_out;
assign out[3] = _U1648_out;
assign out[2] = _U1647_out;
assign out[1] = _U1646_out;
assign out[0] = _U1645_out;
endmodule

module array_delay_U1637 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1638_out;
wire [15:0] _U1639_out;
wire [15:0] _U1640_out;
wire [15:0] _U1641_out;
wire [15:0] _U1642_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1638 (
    .in(in[0]),
    .clk(clk),
    .out(_U1638_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1639 (
    .in(in[1]),
    .clk(clk),
    .out(_U1639_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1640 (
    .in(in[2]),
    .clk(clk),
    .out(_U1640_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1641 (
    .in(in[3]),
    .clk(clk),
    .out(_U1641_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1642 (
    .in(in[4]),
    .clk(clk),
    .out(_U1642_out)
);
assign out[4] = _U1642_out;
assign out[3] = _U1641_out;
assign out[2] = _U1640_out;
assign out[1] = _U1639_out;
assign out[0] = _U1638_out;
endmodule

module array_delay_U1630 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1631_out;
wire [15:0] _U1632_out;
wire [15:0] _U1633_out;
wire [15:0] _U1634_out;
wire [15:0] _U1635_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1631 (
    .in(in[0]),
    .clk(clk),
    .out(_U1631_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1632 (
    .in(in[1]),
    .clk(clk),
    .out(_U1632_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1633 (
    .in(in[2]),
    .clk(clk),
    .out(_U1633_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1634 (
    .in(in[3]),
    .clk(clk),
    .out(_U1634_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1635 (
    .in(in[4]),
    .clk(clk),
    .out(_U1635_out)
);
assign out[4] = _U1635_out;
assign out[3] = _U1634_out;
assign out[2] = _U1633_out;
assign out[1] = _U1632_out;
assign out[0] = _U1631_out;
endmodule

module array_delay_U1623 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1624_out;
wire [15:0] _U1625_out;
wire [15:0] _U1626_out;
wire [15:0] _U1627_out;
wire [15:0] _U1628_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1624 (
    .in(in[0]),
    .clk(clk),
    .out(_U1624_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1625 (
    .in(in[1]),
    .clk(clk),
    .out(_U1625_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1626 (
    .in(in[2]),
    .clk(clk),
    .out(_U1626_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1627 (
    .in(in[3]),
    .clk(clk),
    .out(_U1627_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1628 (
    .in(in[4]),
    .clk(clk),
    .out(_U1628_out)
);
assign out[4] = _U1628_out;
assign out[3] = _U1627_out;
assign out[2] = _U1626_out;
assign out[1] = _U1625_out;
assign out[0] = _U1624_out;
endmodule

module array_delay_U1616 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1617_out;
wire [15:0] _U1618_out;
wire [15:0] _U1619_out;
wire [15:0] _U1620_out;
wire [15:0] _U1621_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1617 (
    .in(in[0]),
    .clk(clk),
    .out(_U1617_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1618 (
    .in(in[1]),
    .clk(clk),
    .out(_U1618_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1619 (
    .in(in[2]),
    .clk(clk),
    .out(_U1619_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1620 (
    .in(in[3]),
    .clk(clk),
    .out(_U1620_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1621 (
    .in(in[4]),
    .clk(clk),
    .out(_U1621_out)
);
assign out[4] = _U1621_out;
assign out[3] = _U1620_out;
assign out[2] = _U1619_out;
assign out[1] = _U1618_out;
assign out[0] = _U1617_out;
endmodule

module array_delay_U1609 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1610_out;
wire [15:0] _U1611_out;
wire [15:0] _U1612_out;
wire [15:0] _U1613_out;
wire [15:0] _U1614_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1610 (
    .in(in[0]),
    .clk(clk),
    .out(_U1610_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1611 (
    .in(in[1]),
    .clk(clk),
    .out(_U1611_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1612 (
    .in(in[2]),
    .clk(clk),
    .out(_U1612_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1613 (
    .in(in[3]),
    .clk(clk),
    .out(_U1613_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1614 (
    .in(in[4]),
    .clk(clk),
    .out(_U1614_out)
);
assign out[4] = _U1614_out;
assign out[3] = _U1613_out;
assign out[2] = _U1612_out;
assign out[1] = _U1611_out;
assign out[0] = _U1610_out;
endmodule

module array_delay_U1602 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1603_out;
wire [15:0] _U1604_out;
wire [15:0] _U1605_out;
wire [15:0] _U1606_out;
wire [15:0] _U1607_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1603 (
    .in(in[0]),
    .clk(clk),
    .out(_U1603_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1604 (
    .in(in[1]),
    .clk(clk),
    .out(_U1604_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1605 (
    .in(in[2]),
    .clk(clk),
    .out(_U1605_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1606 (
    .in(in[3]),
    .clk(clk),
    .out(_U1606_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1607 (
    .in(in[4]),
    .clk(clk),
    .out(_U1607_out)
);
assign out[4] = _U1607_out;
assign out[3] = _U1606_out;
assign out[2] = _U1605_out;
assign out[1] = _U1604_out;
assign out[0] = _U1603_out;
endmodule

module array_delay_U1576 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1577_out;
wire [15:0] _U1578_out;
wire [15:0] _U1579_out;
wire [15:0] _U1580_out;
wire [15:0] _U1581_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1577 (
    .in(in[0]),
    .clk(clk),
    .out(_U1577_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1578 (
    .in(in[1]),
    .clk(clk),
    .out(_U1578_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1579 (
    .in(in[2]),
    .clk(clk),
    .out(_U1579_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1580 (
    .in(in[3]),
    .clk(clk),
    .out(_U1580_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1581 (
    .in(in[4]),
    .clk(clk),
    .out(_U1581_out)
);
assign out[4] = _U1581_out;
assign out[3] = _U1580_out;
assign out[2] = _U1579_out;
assign out[1] = _U1578_out;
assign out[0] = _U1577_out;
endmodule

module array_delay_U1569 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1570_out;
wire [15:0] _U1571_out;
wire [15:0] _U1572_out;
wire [15:0] _U1573_out;
wire [15:0] _U1574_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1570 (
    .in(in[0]),
    .clk(clk),
    .out(_U1570_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1571 (
    .in(in[1]),
    .clk(clk),
    .out(_U1571_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1572 (
    .in(in[2]),
    .clk(clk),
    .out(_U1572_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1573 (
    .in(in[3]),
    .clk(clk),
    .out(_U1573_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1574 (
    .in(in[4]),
    .clk(clk),
    .out(_U1574_out)
);
assign out[4] = _U1574_out;
assign out[3] = _U1573_out;
assign out[2] = _U1572_out;
assign out[1] = _U1571_out;
assign out[0] = _U1570_out;
endmodule

module array_delay_U1526 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1527_out;
wire [15:0] _U1528_out;
wire [15:0] _U1529_out;
wire [15:0] _U1530_out;
wire [15:0] _U1531_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1527 (
    .in(in[0]),
    .clk(clk),
    .out(_U1527_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1528 (
    .in(in[1]),
    .clk(clk),
    .out(_U1528_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1529 (
    .in(in[2]),
    .clk(clk),
    .out(_U1529_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1530 (
    .in(in[3]),
    .clk(clk),
    .out(_U1530_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1531 (
    .in(in[4]),
    .clk(clk),
    .out(_U1531_out)
);
assign out[4] = _U1531_out;
assign out[3] = _U1530_out;
assign out[2] = _U1529_out;
assign out[1] = _U1528_out;
assign out[0] = _U1527_out;
endmodule

module array_delay_U1519 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1520_out;
wire [15:0] _U1521_out;
wire [15:0] _U1522_out;
wire [15:0] _U1523_out;
wire [15:0] _U1524_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1520 (
    .in(in[0]),
    .clk(clk),
    .out(_U1520_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1521 (
    .in(in[1]),
    .clk(clk),
    .out(_U1521_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1522 (
    .in(in[2]),
    .clk(clk),
    .out(_U1522_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1523 (
    .in(in[3]),
    .clk(clk),
    .out(_U1523_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1524 (
    .in(in[4]),
    .clk(clk),
    .out(_U1524_out)
);
assign out[4] = _U1524_out;
assign out[3] = _U1523_out;
assign out[2] = _U1522_out;
assign out[1] = _U1521_out;
assign out[0] = _U1520_out;
endmodule

module array_delay_U1512 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1513_out;
wire [15:0] _U1514_out;
wire [15:0] _U1515_out;
wire [15:0] _U1516_out;
wire [15:0] _U1517_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1513 (
    .in(in[0]),
    .clk(clk),
    .out(_U1513_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1514 (
    .in(in[1]),
    .clk(clk),
    .out(_U1514_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1515 (
    .in(in[2]),
    .clk(clk),
    .out(_U1515_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1516 (
    .in(in[3]),
    .clk(clk),
    .out(_U1516_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1517 (
    .in(in[4]),
    .clk(clk),
    .out(_U1517_out)
);
assign out[4] = _U1517_out;
assign out[3] = _U1516_out;
assign out[2] = _U1515_out;
assign out[1] = _U1514_out;
assign out[0] = _U1513_out;
endmodule

module array_delay_U1505 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1506_out;
wire [15:0] _U1507_out;
wire [15:0] _U1508_out;
wire [15:0] _U1509_out;
wire [15:0] _U1510_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1506 (
    .in(in[0]),
    .clk(clk),
    .out(_U1506_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1507 (
    .in(in[1]),
    .clk(clk),
    .out(_U1507_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1508 (
    .in(in[2]),
    .clk(clk),
    .out(_U1508_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1509 (
    .in(in[3]),
    .clk(clk),
    .out(_U1509_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1510 (
    .in(in[4]),
    .clk(clk),
    .out(_U1510_out)
);
assign out[4] = _U1510_out;
assign out[3] = _U1509_out;
assign out[2] = _U1508_out;
assign out[1] = _U1507_out;
assign out[0] = _U1506_out;
endmodule

module array_delay_U1498 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1499_out;
wire [15:0] _U1500_out;
wire [15:0] _U1501_out;
wire [15:0] _U1502_out;
wire [15:0] _U1503_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1499 (
    .in(in[0]),
    .clk(clk),
    .out(_U1499_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1500 (
    .in(in[1]),
    .clk(clk),
    .out(_U1500_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1501 (
    .in(in[2]),
    .clk(clk),
    .out(_U1501_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1502 (
    .in(in[3]),
    .clk(clk),
    .out(_U1502_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1503 (
    .in(in[4]),
    .clk(clk),
    .out(_U1503_out)
);
assign out[4] = _U1503_out;
assign out[3] = _U1502_out;
assign out[2] = _U1501_out;
assign out[1] = _U1500_out;
assign out[0] = _U1499_out;
endmodule

module array_delay_U1491 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1492_out;
wire [15:0] _U1493_out;
wire [15:0] _U1494_out;
wire [15:0] _U1495_out;
wire [15:0] _U1496_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1492 (
    .in(in[0]),
    .clk(clk),
    .out(_U1492_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1493 (
    .in(in[1]),
    .clk(clk),
    .out(_U1493_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1494 (
    .in(in[2]),
    .clk(clk),
    .out(_U1494_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1495 (
    .in(in[3]),
    .clk(clk),
    .out(_U1495_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1496 (
    .in(in[4]),
    .clk(clk),
    .out(_U1496_out)
);
assign out[4] = _U1496_out;
assign out[3] = _U1495_out;
assign out[2] = _U1494_out;
assign out[1] = _U1493_out;
assign out[0] = _U1492_out;
endmodule

module array_delay_U1484 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1485_out;
wire [15:0] _U1486_out;
wire [15:0] _U1487_out;
wire [15:0] _U1488_out;
wire [15:0] _U1489_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1485 (
    .in(in[0]),
    .clk(clk),
    .out(_U1485_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1486 (
    .in(in[1]),
    .clk(clk),
    .out(_U1486_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1487 (
    .in(in[2]),
    .clk(clk),
    .out(_U1487_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1488 (
    .in(in[3]),
    .clk(clk),
    .out(_U1488_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1489 (
    .in(in[4]),
    .clk(clk),
    .out(_U1489_out)
);
assign out[4] = _U1489_out;
assign out[3] = _U1488_out;
assign out[2] = _U1487_out;
assign out[1] = _U1486_out;
assign out[0] = _U1485_out;
endmodule

module array_delay_U1477 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1478_out;
wire [15:0] _U1479_out;
wire [15:0] _U1480_out;
wire [15:0] _U1481_out;
wire [15:0] _U1482_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1478 (
    .in(in[0]),
    .clk(clk),
    .out(_U1478_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1479 (
    .in(in[1]),
    .clk(clk),
    .out(_U1479_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1480 (
    .in(in[2]),
    .clk(clk),
    .out(_U1480_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1481 (
    .in(in[3]),
    .clk(clk),
    .out(_U1481_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1482 (
    .in(in[4]),
    .clk(clk),
    .out(_U1482_out)
);
assign out[4] = _U1482_out;
assign out[3] = _U1481_out;
assign out[2] = _U1480_out;
assign out[1] = _U1479_out;
assign out[0] = _U1478_out;
endmodule

module array_delay_U1470 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1471_out;
wire [15:0] _U1472_out;
wire [15:0] _U1473_out;
wire [15:0] _U1474_out;
wire [15:0] _U1475_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1471 (
    .in(in[0]),
    .clk(clk),
    .out(_U1471_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1472 (
    .in(in[1]),
    .clk(clk),
    .out(_U1472_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1473 (
    .in(in[2]),
    .clk(clk),
    .out(_U1473_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1474 (
    .in(in[3]),
    .clk(clk),
    .out(_U1474_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1475 (
    .in(in[4]),
    .clk(clk),
    .out(_U1475_out)
);
assign out[4] = _U1475_out;
assign out[3] = _U1474_out;
assign out[2] = _U1473_out;
assign out[1] = _U1472_out;
assign out[0] = _U1471_out;
endmodule

module array_delay_U1463 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1464_out;
wire [15:0] _U1465_out;
wire [15:0] _U1466_out;
wire [15:0] _U1467_out;
wire [15:0] _U1468_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1464 (
    .in(in[0]),
    .clk(clk),
    .out(_U1464_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1465 (
    .in(in[1]),
    .clk(clk),
    .out(_U1465_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1466 (
    .in(in[2]),
    .clk(clk),
    .out(_U1466_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1467 (
    .in(in[3]),
    .clk(clk),
    .out(_U1467_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1468 (
    .in(in[4]),
    .clk(clk),
    .out(_U1468_out)
);
assign out[4] = _U1468_out;
assign out[3] = _U1467_out;
assign out[2] = _U1466_out;
assign out[1] = _U1465_out;
assign out[0] = _U1464_out;
endmodule

module array_delay_U1456 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1457_out;
wire [15:0] _U1458_out;
wire [15:0] _U1459_out;
wire [15:0] _U1460_out;
wire [15:0] _U1461_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1457 (
    .in(in[0]),
    .clk(clk),
    .out(_U1457_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1458 (
    .in(in[1]),
    .clk(clk),
    .out(_U1458_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1459 (
    .in(in[2]),
    .clk(clk),
    .out(_U1459_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1460 (
    .in(in[3]),
    .clk(clk),
    .out(_U1460_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1461 (
    .in(in[4]),
    .clk(clk),
    .out(_U1461_out)
);
assign out[4] = _U1461_out;
assign out[3] = _U1460_out;
assign out[2] = _U1459_out;
assign out[1] = _U1458_out;
assign out[0] = _U1457_out;
endmodule

module array_delay_U1449 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1450_out;
wire [15:0] _U1451_out;
wire [15:0] _U1452_out;
wire [15:0] _U1453_out;
wire [15:0] _U1454_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1450 (
    .in(in[0]),
    .clk(clk),
    .out(_U1450_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1451 (
    .in(in[1]),
    .clk(clk),
    .out(_U1451_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1452 (
    .in(in[2]),
    .clk(clk),
    .out(_U1452_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1453 (
    .in(in[3]),
    .clk(clk),
    .out(_U1453_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1454 (
    .in(in[4]),
    .clk(clk),
    .out(_U1454_out)
);
assign out[4] = _U1454_out;
assign out[3] = _U1453_out;
assign out[2] = _U1452_out;
assign out[1] = _U1451_out;
assign out[0] = _U1450_out;
endmodule

module array_delay_U1442 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1443_out;
wire [15:0] _U1444_out;
wire [15:0] _U1445_out;
wire [15:0] _U1446_out;
wire [15:0] _U1447_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1443 (
    .in(in[0]),
    .clk(clk),
    .out(_U1443_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1444 (
    .in(in[1]),
    .clk(clk),
    .out(_U1444_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1445 (
    .in(in[2]),
    .clk(clk),
    .out(_U1445_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1446 (
    .in(in[3]),
    .clk(clk),
    .out(_U1446_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1447 (
    .in(in[4]),
    .clk(clk),
    .out(_U1447_out)
);
assign out[4] = _U1447_out;
assign out[3] = _U1446_out;
assign out[2] = _U1445_out;
assign out[1] = _U1444_out;
assign out[0] = _U1443_out;
endmodule

module array_delay_U1435 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1436_out;
wire [15:0] _U1437_out;
wire [15:0] _U1438_out;
wire [15:0] _U1439_out;
wire [15:0] _U1440_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1436 (
    .in(in[0]),
    .clk(clk),
    .out(_U1436_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1437 (
    .in(in[1]),
    .clk(clk),
    .out(_U1437_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1438 (
    .in(in[2]),
    .clk(clk),
    .out(_U1438_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1439 (
    .in(in[3]),
    .clk(clk),
    .out(_U1439_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1440 (
    .in(in[4]),
    .clk(clk),
    .out(_U1440_out)
);
assign out[4] = _U1440_out;
assign out[3] = _U1439_out;
assign out[2] = _U1438_out;
assign out[1] = _U1437_out;
assign out[0] = _U1436_out;
endmodule

module array_delay_U1428 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1429_out;
wire [15:0] _U1430_out;
wire [15:0] _U1431_out;
wire [15:0] _U1432_out;
wire [15:0] _U1433_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1429 (
    .in(in[0]),
    .clk(clk),
    .out(_U1429_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1430 (
    .in(in[1]),
    .clk(clk),
    .out(_U1430_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1431 (
    .in(in[2]),
    .clk(clk),
    .out(_U1431_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1432 (
    .in(in[3]),
    .clk(clk),
    .out(_U1432_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1433 (
    .in(in[4]),
    .clk(clk),
    .out(_U1433_out)
);
assign out[4] = _U1433_out;
assign out[3] = _U1432_out;
assign out[2] = _U1431_out;
assign out[1] = _U1430_out;
assign out[0] = _U1429_out;
endmodule

module array_delay_U1421 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1422_out;
wire [15:0] _U1423_out;
wire [15:0] _U1424_out;
wire [15:0] _U1425_out;
wire [15:0] _U1426_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1422 (
    .in(in[0]),
    .clk(clk),
    .out(_U1422_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1423 (
    .in(in[1]),
    .clk(clk),
    .out(_U1423_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1424 (
    .in(in[2]),
    .clk(clk),
    .out(_U1424_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1425 (
    .in(in[3]),
    .clk(clk),
    .out(_U1425_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1426 (
    .in(in[4]),
    .clk(clk),
    .out(_U1426_out)
);
assign out[4] = _U1426_out;
assign out[3] = _U1425_out;
assign out[2] = _U1424_out;
assign out[1] = _U1423_out;
assign out[0] = _U1422_out;
endmodule

module array_delay_U1414 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1415_out;
wire [15:0] _U1416_out;
wire [15:0] _U1417_out;
wire [15:0] _U1418_out;
wire [15:0] _U1419_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1415 (
    .in(in[0]),
    .clk(clk),
    .out(_U1415_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1416 (
    .in(in[1]),
    .clk(clk),
    .out(_U1416_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1417 (
    .in(in[2]),
    .clk(clk),
    .out(_U1417_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1418 (
    .in(in[3]),
    .clk(clk),
    .out(_U1418_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1419 (
    .in(in[4]),
    .clk(clk),
    .out(_U1419_out)
);
assign out[4] = _U1419_out;
assign out[3] = _U1418_out;
assign out[2] = _U1417_out;
assign out[1] = _U1416_out;
assign out[0] = _U1415_out;
endmodule

module array_delay_U1388 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1389_out;
wire [15:0] _U1390_out;
wire [15:0] _U1391_out;
wire [15:0] _U1392_out;
wire [15:0] _U1393_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1389 (
    .in(in[0]),
    .clk(clk),
    .out(_U1389_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1390 (
    .in(in[1]),
    .clk(clk),
    .out(_U1390_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1391 (
    .in(in[2]),
    .clk(clk),
    .out(_U1391_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1392 (
    .in(in[3]),
    .clk(clk),
    .out(_U1392_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1393 (
    .in(in[4]),
    .clk(clk),
    .out(_U1393_out)
);
assign out[4] = _U1393_out;
assign out[3] = _U1392_out;
assign out[2] = _U1391_out;
assign out[1] = _U1390_out;
assign out[0] = _U1389_out;
endmodule

module array_delay_U1381 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1382_out;
wire [15:0] _U1383_out;
wire [15:0] _U1384_out;
wire [15:0] _U1385_out;
wire [15:0] _U1386_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1382 (
    .in(in[0]),
    .clk(clk),
    .out(_U1382_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1383 (
    .in(in[1]),
    .clk(clk),
    .out(_U1383_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1384 (
    .in(in[2]),
    .clk(clk),
    .out(_U1384_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1385 (
    .in(in[3]),
    .clk(clk),
    .out(_U1385_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1386 (
    .in(in[4]),
    .clk(clk),
    .out(_U1386_out)
);
assign out[4] = _U1386_out;
assign out[3] = _U1385_out;
assign out[2] = _U1384_out;
assign out[1] = _U1383_out;
assign out[0] = _U1382_out;
endmodule

module array_delay_U1338 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1339_out;
wire [15:0] _U1340_out;
wire [15:0] _U1341_out;
wire [15:0] _U1342_out;
wire [15:0] _U1343_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1339 (
    .in(in[0]),
    .clk(clk),
    .out(_U1339_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1340 (
    .in(in[1]),
    .clk(clk),
    .out(_U1340_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1341 (
    .in(in[2]),
    .clk(clk),
    .out(_U1341_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1342 (
    .in(in[3]),
    .clk(clk),
    .out(_U1342_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1343 (
    .in(in[4]),
    .clk(clk),
    .out(_U1343_out)
);
assign out[4] = _U1343_out;
assign out[3] = _U1342_out;
assign out[2] = _U1341_out;
assign out[1] = _U1340_out;
assign out[0] = _U1339_out;
endmodule

module array_delay_U1331 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1332_out;
wire [15:0] _U1333_out;
wire [15:0] _U1334_out;
wire [15:0] _U1335_out;
wire [15:0] _U1336_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1332 (
    .in(in[0]),
    .clk(clk),
    .out(_U1332_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1333 (
    .in(in[1]),
    .clk(clk),
    .out(_U1333_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1334 (
    .in(in[2]),
    .clk(clk),
    .out(_U1334_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1335 (
    .in(in[3]),
    .clk(clk),
    .out(_U1335_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1336 (
    .in(in[4]),
    .clk(clk),
    .out(_U1336_out)
);
assign out[4] = _U1336_out;
assign out[3] = _U1335_out;
assign out[2] = _U1334_out;
assign out[1] = _U1333_out;
assign out[0] = _U1332_out;
endmodule

module array_delay_U1324 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1325_out;
wire [15:0] _U1326_out;
wire [15:0] _U1327_out;
wire [15:0] _U1328_out;
wire [15:0] _U1329_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1325 (
    .in(in[0]),
    .clk(clk),
    .out(_U1325_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1326 (
    .in(in[1]),
    .clk(clk),
    .out(_U1326_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1327 (
    .in(in[2]),
    .clk(clk),
    .out(_U1327_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1328 (
    .in(in[3]),
    .clk(clk),
    .out(_U1328_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1329 (
    .in(in[4]),
    .clk(clk),
    .out(_U1329_out)
);
assign out[4] = _U1329_out;
assign out[3] = _U1328_out;
assign out[2] = _U1327_out;
assign out[1] = _U1326_out;
assign out[0] = _U1325_out;
endmodule

module array_delay_U1317 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1318_out;
wire [15:0] _U1319_out;
wire [15:0] _U1320_out;
wire [15:0] _U1321_out;
wire [15:0] _U1322_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1318 (
    .in(in[0]),
    .clk(clk),
    .out(_U1318_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1319 (
    .in(in[1]),
    .clk(clk),
    .out(_U1319_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1320 (
    .in(in[2]),
    .clk(clk),
    .out(_U1320_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1321 (
    .in(in[3]),
    .clk(clk),
    .out(_U1321_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1322 (
    .in(in[4]),
    .clk(clk),
    .out(_U1322_out)
);
assign out[4] = _U1322_out;
assign out[3] = _U1321_out;
assign out[2] = _U1320_out;
assign out[1] = _U1319_out;
assign out[0] = _U1318_out;
endmodule

module array_delay_U1310 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1311_out;
wire [15:0] _U1312_out;
wire [15:0] _U1313_out;
wire [15:0] _U1314_out;
wire [15:0] _U1315_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1311 (
    .in(in[0]),
    .clk(clk),
    .out(_U1311_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1312 (
    .in(in[1]),
    .clk(clk),
    .out(_U1312_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1313 (
    .in(in[2]),
    .clk(clk),
    .out(_U1313_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1314 (
    .in(in[3]),
    .clk(clk),
    .out(_U1314_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1315 (
    .in(in[4]),
    .clk(clk),
    .out(_U1315_out)
);
assign out[4] = _U1315_out;
assign out[3] = _U1314_out;
assign out[2] = _U1313_out;
assign out[1] = _U1312_out;
assign out[0] = _U1311_out;
endmodule

module array_delay_U1303 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1304_out;
wire [15:0] _U1305_out;
wire [15:0] _U1306_out;
wire [15:0] _U1307_out;
wire [15:0] _U1308_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1304 (
    .in(in[0]),
    .clk(clk),
    .out(_U1304_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1305 (
    .in(in[1]),
    .clk(clk),
    .out(_U1305_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1306 (
    .in(in[2]),
    .clk(clk),
    .out(_U1306_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1307 (
    .in(in[3]),
    .clk(clk),
    .out(_U1307_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1308 (
    .in(in[4]),
    .clk(clk),
    .out(_U1308_out)
);
assign out[4] = _U1308_out;
assign out[3] = _U1307_out;
assign out[2] = _U1306_out;
assign out[1] = _U1305_out;
assign out[0] = _U1304_out;
endmodule

module array_delay_U1296 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1297_out;
wire [15:0] _U1298_out;
wire [15:0] _U1299_out;
wire [15:0] _U1300_out;
wire [15:0] _U1301_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1297 (
    .in(in[0]),
    .clk(clk),
    .out(_U1297_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1298 (
    .in(in[1]),
    .clk(clk),
    .out(_U1298_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1299 (
    .in(in[2]),
    .clk(clk),
    .out(_U1299_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1300 (
    .in(in[3]),
    .clk(clk),
    .out(_U1300_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1301 (
    .in(in[4]),
    .clk(clk),
    .out(_U1301_out)
);
assign out[4] = _U1301_out;
assign out[3] = _U1300_out;
assign out[2] = _U1299_out;
assign out[1] = _U1298_out;
assign out[0] = _U1297_out;
endmodule

module array_delay_U1289 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1290_out;
wire [15:0] _U1291_out;
wire [15:0] _U1292_out;
wire [15:0] _U1293_out;
wire [15:0] _U1294_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1290 (
    .in(in[0]),
    .clk(clk),
    .out(_U1290_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1291 (
    .in(in[1]),
    .clk(clk),
    .out(_U1291_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1292 (
    .in(in[2]),
    .clk(clk),
    .out(_U1292_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1293 (
    .in(in[3]),
    .clk(clk),
    .out(_U1293_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1294 (
    .in(in[4]),
    .clk(clk),
    .out(_U1294_out)
);
assign out[4] = _U1294_out;
assign out[3] = _U1293_out;
assign out[2] = _U1292_out;
assign out[1] = _U1291_out;
assign out[0] = _U1290_out;
endmodule

module array_delay_U1282 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1283_out;
wire [15:0] _U1284_out;
wire [15:0] _U1285_out;
wire [15:0] _U1286_out;
wire [15:0] _U1287_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1283 (
    .in(in[0]),
    .clk(clk),
    .out(_U1283_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1284 (
    .in(in[1]),
    .clk(clk),
    .out(_U1284_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1285 (
    .in(in[2]),
    .clk(clk),
    .out(_U1285_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1286 (
    .in(in[3]),
    .clk(clk),
    .out(_U1286_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1287 (
    .in(in[4]),
    .clk(clk),
    .out(_U1287_out)
);
assign out[4] = _U1287_out;
assign out[3] = _U1286_out;
assign out[2] = _U1285_out;
assign out[1] = _U1284_out;
assign out[0] = _U1283_out;
endmodule

module array_delay_U1275 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1276_out;
wire [15:0] _U1277_out;
wire [15:0] _U1278_out;
wire [15:0] _U1279_out;
wire [15:0] _U1280_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1276 (
    .in(in[0]),
    .clk(clk),
    .out(_U1276_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1277 (
    .in(in[1]),
    .clk(clk),
    .out(_U1277_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1278 (
    .in(in[2]),
    .clk(clk),
    .out(_U1278_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1279 (
    .in(in[3]),
    .clk(clk),
    .out(_U1279_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1280 (
    .in(in[4]),
    .clk(clk),
    .out(_U1280_out)
);
assign out[4] = _U1280_out;
assign out[3] = _U1279_out;
assign out[2] = _U1278_out;
assign out[1] = _U1277_out;
assign out[0] = _U1276_out;
endmodule

module array_delay_U1268 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1269_out;
wire [15:0] _U1270_out;
wire [15:0] _U1271_out;
wire [15:0] _U1272_out;
wire [15:0] _U1273_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1269 (
    .in(in[0]),
    .clk(clk),
    .out(_U1269_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1270 (
    .in(in[1]),
    .clk(clk),
    .out(_U1270_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1271 (
    .in(in[2]),
    .clk(clk),
    .out(_U1271_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1272 (
    .in(in[3]),
    .clk(clk),
    .out(_U1272_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1273 (
    .in(in[4]),
    .clk(clk),
    .out(_U1273_out)
);
assign out[4] = _U1273_out;
assign out[3] = _U1272_out;
assign out[2] = _U1271_out;
assign out[1] = _U1270_out;
assign out[0] = _U1269_out;
endmodule

module array_delay_U1261 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1262_out;
wire [15:0] _U1263_out;
wire [15:0] _U1264_out;
wire [15:0] _U1265_out;
wire [15:0] _U1266_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1262 (
    .in(in[0]),
    .clk(clk),
    .out(_U1262_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1263 (
    .in(in[1]),
    .clk(clk),
    .out(_U1263_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1264 (
    .in(in[2]),
    .clk(clk),
    .out(_U1264_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1265 (
    .in(in[3]),
    .clk(clk),
    .out(_U1265_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1266 (
    .in(in[4]),
    .clk(clk),
    .out(_U1266_out)
);
assign out[4] = _U1266_out;
assign out[3] = _U1265_out;
assign out[2] = _U1264_out;
assign out[1] = _U1263_out;
assign out[0] = _U1262_out;
endmodule

module array_delay_U1254 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1255_out;
wire [15:0] _U1256_out;
wire [15:0] _U1257_out;
wire [15:0] _U1258_out;
wire [15:0] _U1259_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1255 (
    .in(in[0]),
    .clk(clk),
    .out(_U1255_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1256 (
    .in(in[1]),
    .clk(clk),
    .out(_U1256_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1257 (
    .in(in[2]),
    .clk(clk),
    .out(_U1257_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1258 (
    .in(in[3]),
    .clk(clk),
    .out(_U1258_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1259 (
    .in(in[4]),
    .clk(clk),
    .out(_U1259_out)
);
assign out[4] = _U1259_out;
assign out[3] = _U1258_out;
assign out[2] = _U1257_out;
assign out[1] = _U1256_out;
assign out[0] = _U1255_out;
endmodule

module array_delay_U1247 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1248_out;
wire [15:0] _U1249_out;
wire [15:0] _U1250_out;
wire [15:0] _U1251_out;
wire [15:0] _U1252_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1248 (
    .in(in[0]),
    .clk(clk),
    .out(_U1248_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1249 (
    .in(in[1]),
    .clk(clk),
    .out(_U1249_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1250 (
    .in(in[2]),
    .clk(clk),
    .out(_U1250_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1251 (
    .in(in[3]),
    .clk(clk),
    .out(_U1251_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1252 (
    .in(in[4]),
    .clk(clk),
    .out(_U1252_out)
);
assign out[4] = _U1252_out;
assign out[3] = _U1251_out;
assign out[2] = _U1250_out;
assign out[1] = _U1249_out;
assign out[0] = _U1248_out;
endmodule

module array_delay_U1240 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1241_out;
wire [15:0] _U1242_out;
wire [15:0] _U1243_out;
wire [15:0] _U1244_out;
wire [15:0] _U1245_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1241 (
    .in(in[0]),
    .clk(clk),
    .out(_U1241_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1242 (
    .in(in[1]),
    .clk(clk),
    .out(_U1242_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1243 (
    .in(in[2]),
    .clk(clk),
    .out(_U1243_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1244 (
    .in(in[3]),
    .clk(clk),
    .out(_U1244_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1245 (
    .in(in[4]),
    .clk(clk),
    .out(_U1245_out)
);
assign out[4] = _U1245_out;
assign out[3] = _U1244_out;
assign out[2] = _U1243_out;
assign out[1] = _U1242_out;
assign out[0] = _U1241_out;
endmodule

module array_delay_U1233 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1234_out;
wire [15:0] _U1235_out;
wire [15:0] _U1236_out;
wire [15:0] _U1237_out;
wire [15:0] _U1238_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1234 (
    .in(in[0]),
    .clk(clk),
    .out(_U1234_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1235 (
    .in(in[1]),
    .clk(clk),
    .out(_U1235_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1236 (
    .in(in[2]),
    .clk(clk),
    .out(_U1236_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1237 (
    .in(in[3]),
    .clk(clk),
    .out(_U1237_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1238 (
    .in(in[4]),
    .clk(clk),
    .out(_U1238_out)
);
assign out[4] = _U1238_out;
assign out[3] = _U1237_out;
assign out[2] = _U1236_out;
assign out[1] = _U1235_out;
assign out[0] = _U1234_out;
endmodule

module array_delay_U1226 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1227_out;
wire [15:0] _U1228_out;
wire [15:0] _U1229_out;
wire [15:0] _U1230_out;
wire [15:0] _U1231_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1227 (
    .in(in[0]),
    .clk(clk),
    .out(_U1227_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1228 (
    .in(in[1]),
    .clk(clk),
    .out(_U1228_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1229 (
    .in(in[2]),
    .clk(clk),
    .out(_U1229_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1230 (
    .in(in[3]),
    .clk(clk),
    .out(_U1230_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1231 (
    .in(in[4]),
    .clk(clk),
    .out(_U1231_out)
);
assign out[4] = _U1231_out;
assign out[3] = _U1230_out;
assign out[2] = _U1229_out;
assign out[1] = _U1228_out;
assign out[0] = _U1227_out;
endmodule

module array_delay_U1200 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1201_out;
wire [15:0] _U1202_out;
wire [15:0] _U1203_out;
wire [15:0] _U1204_out;
wire [15:0] _U1205_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1201 (
    .in(in[0]),
    .clk(clk),
    .out(_U1201_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1202 (
    .in(in[1]),
    .clk(clk),
    .out(_U1202_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1203 (
    .in(in[2]),
    .clk(clk),
    .out(_U1203_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1204 (
    .in(in[3]),
    .clk(clk),
    .out(_U1204_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1205 (
    .in(in[4]),
    .clk(clk),
    .out(_U1205_out)
);
assign out[4] = _U1205_out;
assign out[3] = _U1204_out;
assign out[2] = _U1203_out;
assign out[1] = _U1202_out;
assign out[0] = _U1201_out;
endmodule

module array_delay_U1193 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1194_out;
wire [15:0] _U1195_out;
wire [15:0] _U1196_out;
wire [15:0] _U1197_out;
wire [15:0] _U1198_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1194 (
    .in(in[0]),
    .clk(clk),
    .out(_U1194_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1195 (
    .in(in[1]),
    .clk(clk),
    .out(_U1195_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1196 (
    .in(in[2]),
    .clk(clk),
    .out(_U1196_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1197 (
    .in(in[3]),
    .clk(clk),
    .out(_U1197_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1198 (
    .in(in[4]),
    .clk(clk),
    .out(_U1198_out)
);
assign out[4] = _U1198_out;
assign out[3] = _U1197_out;
assign out[2] = _U1196_out;
assign out[1] = _U1195_out;
assign out[0] = _U1194_out;
endmodule

module array_delay_U1150 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1151_out;
wire [15:0] _U1152_out;
wire [15:0] _U1153_out;
wire [15:0] _U1154_out;
wire [15:0] _U1155_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1151 (
    .in(in[0]),
    .clk(clk),
    .out(_U1151_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1152 (
    .in(in[1]),
    .clk(clk),
    .out(_U1152_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1153 (
    .in(in[2]),
    .clk(clk),
    .out(_U1153_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1154 (
    .in(in[3]),
    .clk(clk),
    .out(_U1154_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1155 (
    .in(in[4]),
    .clk(clk),
    .out(_U1155_out)
);
assign out[4] = _U1155_out;
assign out[3] = _U1154_out;
assign out[2] = _U1153_out;
assign out[1] = _U1152_out;
assign out[0] = _U1151_out;
endmodule

module array_delay_U1143 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1144_out;
wire [15:0] _U1145_out;
wire [15:0] _U1146_out;
wire [15:0] _U1147_out;
wire [15:0] _U1148_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1144 (
    .in(in[0]),
    .clk(clk),
    .out(_U1144_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1145 (
    .in(in[1]),
    .clk(clk),
    .out(_U1145_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1146 (
    .in(in[2]),
    .clk(clk),
    .out(_U1146_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1147 (
    .in(in[3]),
    .clk(clk),
    .out(_U1147_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1148 (
    .in(in[4]),
    .clk(clk),
    .out(_U1148_out)
);
assign out[4] = _U1148_out;
assign out[3] = _U1147_out;
assign out[2] = _U1146_out;
assign out[1] = _U1145_out;
assign out[0] = _U1144_out;
endmodule

module array_delay_U1136 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1137_out;
wire [15:0] _U1138_out;
wire [15:0] _U1139_out;
wire [15:0] _U1140_out;
wire [15:0] _U1141_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1137 (
    .in(in[0]),
    .clk(clk),
    .out(_U1137_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1138 (
    .in(in[1]),
    .clk(clk),
    .out(_U1138_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1139 (
    .in(in[2]),
    .clk(clk),
    .out(_U1139_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1140 (
    .in(in[3]),
    .clk(clk),
    .out(_U1140_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1141 (
    .in(in[4]),
    .clk(clk),
    .out(_U1141_out)
);
assign out[4] = _U1141_out;
assign out[3] = _U1140_out;
assign out[2] = _U1139_out;
assign out[1] = _U1138_out;
assign out[0] = _U1137_out;
endmodule

module array_delay_U1129 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1130_out;
wire [15:0] _U1131_out;
wire [15:0] _U1132_out;
wire [15:0] _U1133_out;
wire [15:0] _U1134_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1130 (
    .in(in[0]),
    .clk(clk),
    .out(_U1130_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1131 (
    .in(in[1]),
    .clk(clk),
    .out(_U1131_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1132 (
    .in(in[2]),
    .clk(clk),
    .out(_U1132_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1133 (
    .in(in[3]),
    .clk(clk),
    .out(_U1133_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1134 (
    .in(in[4]),
    .clk(clk),
    .out(_U1134_out)
);
assign out[4] = _U1134_out;
assign out[3] = _U1133_out;
assign out[2] = _U1132_out;
assign out[1] = _U1131_out;
assign out[0] = _U1130_out;
endmodule

module array_delay_U1122 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1123_out;
wire [15:0] _U1124_out;
wire [15:0] _U1125_out;
wire [15:0] _U1126_out;
wire [15:0] _U1127_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1123 (
    .in(in[0]),
    .clk(clk),
    .out(_U1123_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1124 (
    .in(in[1]),
    .clk(clk),
    .out(_U1124_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1125 (
    .in(in[2]),
    .clk(clk),
    .out(_U1125_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1126 (
    .in(in[3]),
    .clk(clk),
    .out(_U1126_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1127 (
    .in(in[4]),
    .clk(clk),
    .out(_U1127_out)
);
assign out[4] = _U1127_out;
assign out[3] = _U1126_out;
assign out[2] = _U1125_out;
assign out[1] = _U1124_out;
assign out[0] = _U1123_out;
endmodule

module array_delay_U1115 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1116_out;
wire [15:0] _U1117_out;
wire [15:0] _U1118_out;
wire [15:0] _U1119_out;
wire [15:0] _U1120_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1116 (
    .in(in[0]),
    .clk(clk),
    .out(_U1116_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1117 (
    .in(in[1]),
    .clk(clk),
    .out(_U1117_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1118 (
    .in(in[2]),
    .clk(clk),
    .out(_U1118_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1119 (
    .in(in[3]),
    .clk(clk),
    .out(_U1119_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1120 (
    .in(in[4]),
    .clk(clk),
    .out(_U1120_out)
);
assign out[4] = _U1120_out;
assign out[3] = _U1119_out;
assign out[2] = _U1118_out;
assign out[1] = _U1117_out;
assign out[0] = _U1116_out;
endmodule

module array_delay_U1108 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1109_out;
wire [15:0] _U1110_out;
wire [15:0] _U1111_out;
wire [15:0] _U1112_out;
wire [15:0] _U1113_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1109 (
    .in(in[0]),
    .clk(clk),
    .out(_U1109_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1110 (
    .in(in[1]),
    .clk(clk),
    .out(_U1110_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1111 (
    .in(in[2]),
    .clk(clk),
    .out(_U1111_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1112 (
    .in(in[3]),
    .clk(clk),
    .out(_U1112_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1113 (
    .in(in[4]),
    .clk(clk),
    .out(_U1113_out)
);
assign out[4] = _U1113_out;
assign out[3] = _U1112_out;
assign out[2] = _U1111_out;
assign out[1] = _U1110_out;
assign out[0] = _U1109_out;
endmodule

module array_delay_U1101 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1102_out;
wire [15:0] _U1103_out;
wire [15:0] _U1104_out;
wire [15:0] _U1105_out;
wire [15:0] _U1106_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1102 (
    .in(in[0]),
    .clk(clk),
    .out(_U1102_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1103 (
    .in(in[1]),
    .clk(clk),
    .out(_U1103_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1104 (
    .in(in[2]),
    .clk(clk),
    .out(_U1104_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1105 (
    .in(in[3]),
    .clk(clk),
    .out(_U1105_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1106 (
    .in(in[4]),
    .clk(clk),
    .out(_U1106_out)
);
assign out[4] = _U1106_out;
assign out[3] = _U1105_out;
assign out[2] = _U1104_out;
assign out[1] = _U1103_out;
assign out[0] = _U1102_out;
endmodule

module array_delay_U1094 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1095_out;
wire [15:0] _U1096_out;
wire [15:0] _U1097_out;
wire [15:0] _U1098_out;
wire [15:0] _U1099_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1095 (
    .in(in[0]),
    .clk(clk),
    .out(_U1095_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1096 (
    .in(in[1]),
    .clk(clk),
    .out(_U1096_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1097 (
    .in(in[2]),
    .clk(clk),
    .out(_U1097_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1098 (
    .in(in[3]),
    .clk(clk),
    .out(_U1098_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1099 (
    .in(in[4]),
    .clk(clk),
    .out(_U1099_out)
);
assign out[4] = _U1099_out;
assign out[3] = _U1098_out;
assign out[2] = _U1097_out;
assign out[1] = _U1096_out;
assign out[0] = _U1095_out;
endmodule

module array_delay_U1087 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1088_out;
wire [15:0] _U1089_out;
wire [15:0] _U1090_out;
wire [15:0] _U1091_out;
wire [15:0] _U1092_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1088 (
    .in(in[0]),
    .clk(clk),
    .out(_U1088_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1089 (
    .in(in[1]),
    .clk(clk),
    .out(_U1089_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1090 (
    .in(in[2]),
    .clk(clk),
    .out(_U1090_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1091 (
    .in(in[3]),
    .clk(clk),
    .out(_U1091_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1092 (
    .in(in[4]),
    .clk(clk),
    .out(_U1092_out)
);
assign out[4] = _U1092_out;
assign out[3] = _U1091_out;
assign out[2] = _U1090_out;
assign out[1] = _U1089_out;
assign out[0] = _U1088_out;
endmodule

module array_delay_U1080 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1081_out;
wire [15:0] _U1082_out;
wire [15:0] _U1083_out;
wire [15:0] _U1084_out;
wire [15:0] _U1085_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1081 (
    .in(in[0]),
    .clk(clk),
    .out(_U1081_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1082 (
    .in(in[1]),
    .clk(clk),
    .out(_U1082_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1083 (
    .in(in[2]),
    .clk(clk),
    .out(_U1083_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1084 (
    .in(in[3]),
    .clk(clk),
    .out(_U1084_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1085 (
    .in(in[4]),
    .clk(clk),
    .out(_U1085_out)
);
assign out[4] = _U1085_out;
assign out[3] = _U1084_out;
assign out[2] = _U1083_out;
assign out[1] = _U1082_out;
assign out[0] = _U1081_out;
endmodule

module array_delay_U1073 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1074_out;
wire [15:0] _U1075_out;
wire [15:0] _U1076_out;
wire [15:0] _U1077_out;
wire [15:0] _U1078_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1074 (
    .in(in[0]),
    .clk(clk),
    .out(_U1074_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1075 (
    .in(in[1]),
    .clk(clk),
    .out(_U1075_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1076 (
    .in(in[2]),
    .clk(clk),
    .out(_U1076_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1077 (
    .in(in[3]),
    .clk(clk),
    .out(_U1077_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1078 (
    .in(in[4]),
    .clk(clk),
    .out(_U1078_out)
);
assign out[4] = _U1078_out;
assign out[3] = _U1077_out;
assign out[2] = _U1076_out;
assign out[1] = _U1075_out;
assign out[0] = _U1074_out;
endmodule

module array_delay_U1066 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1067_out;
wire [15:0] _U1068_out;
wire [15:0] _U1069_out;
wire [15:0] _U1070_out;
wire [15:0] _U1071_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1067 (
    .in(in[0]),
    .clk(clk),
    .out(_U1067_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1068 (
    .in(in[1]),
    .clk(clk),
    .out(_U1068_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1069 (
    .in(in[2]),
    .clk(clk),
    .out(_U1069_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1070 (
    .in(in[3]),
    .clk(clk),
    .out(_U1070_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1071 (
    .in(in[4]),
    .clk(clk),
    .out(_U1071_out)
);
assign out[4] = _U1071_out;
assign out[3] = _U1070_out;
assign out[2] = _U1069_out;
assign out[1] = _U1068_out;
assign out[0] = _U1067_out;
endmodule

module array_delay_U1059 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1060_out;
wire [15:0] _U1061_out;
wire [15:0] _U1062_out;
wire [15:0] _U1063_out;
wire [15:0] _U1064_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1060 (
    .in(in[0]),
    .clk(clk),
    .out(_U1060_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1061 (
    .in(in[1]),
    .clk(clk),
    .out(_U1061_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1062 (
    .in(in[2]),
    .clk(clk),
    .out(_U1062_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1063 (
    .in(in[3]),
    .clk(clk),
    .out(_U1063_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1064 (
    .in(in[4]),
    .clk(clk),
    .out(_U1064_out)
);
assign out[4] = _U1064_out;
assign out[3] = _U1063_out;
assign out[2] = _U1062_out;
assign out[1] = _U1061_out;
assign out[0] = _U1060_out;
endmodule

module array_delay_U1052 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1053_out;
wire [15:0] _U1054_out;
wire [15:0] _U1055_out;
wire [15:0] _U1056_out;
wire [15:0] _U1057_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1053 (
    .in(in[0]),
    .clk(clk),
    .out(_U1053_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1054 (
    .in(in[1]),
    .clk(clk),
    .out(_U1054_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1055 (
    .in(in[2]),
    .clk(clk),
    .out(_U1055_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1056 (
    .in(in[3]),
    .clk(clk),
    .out(_U1056_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1057 (
    .in(in[4]),
    .clk(clk),
    .out(_U1057_out)
);
assign out[4] = _U1057_out;
assign out[3] = _U1056_out;
assign out[2] = _U1055_out;
assign out[1] = _U1054_out;
assign out[0] = _U1053_out;
endmodule

module array_delay_U1045 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1046_out;
wire [15:0] _U1047_out;
wire [15:0] _U1048_out;
wire [15:0] _U1049_out;
wire [15:0] _U1050_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1046 (
    .in(in[0]),
    .clk(clk),
    .out(_U1046_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1047 (
    .in(in[1]),
    .clk(clk),
    .out(_U1047_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1048 (
    .in(in[2]),
    .clk(clk),
    .out(_U1048_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1049 (
    .in(in[3]),
    .clk(clk),
    .out(_U1049_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1050 (
    .in(in[4]),
    .clk(clk),
    .out(_U1050_out)
);
assign out[4] = _U1050_out;
assign out[3] = _U1049_out;
assign out[2] = _U1048_out;
assign out[1] = _U1047_out;
assign out[0] = _U1046_out;
endmodule

module array_delay_U1038 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1039_out;
wire [15:0] _U1040_out;
wire [15:0] _U1041_out;
wire [15:0] _U1042_out;
wire [15:0] _U1043_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1039 (
    .in(in[0]),
    .clk(clk),
    .out(_U1039_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1040 (
    .in(in[1]),
    .clk(clk),
    .out(_U1040_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1041 (
    .in(in[2]),
    .clk(clk),
    .out(_U1041_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1042 (
    .in(in[3]),
    .clk(clk),
    .out(_U1042_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1043 (
    .in(in[4]),
    .clk(clk),
    .out(_U1043_out)
);
assign out[4] = _U1043_out;
assign out[3] = _U1042_out;
assign out[2] = _U1041_out;
assign out[1] = _U1040_out;
assign out[0] = _U1039_out;
endmodule

module array_delay_U1012 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1013_out;
wire [15:0] _U1014_out;
wire [15:0] _U1015_out;
wire [15:0] _U1016_out;
wire [15:0] _U1017_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1013 (
    .in(in[0]),
    .clk(clk),
    .out(_U1013_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1014 (
    .in(in[1]),
    .clk(clk),
    .out(_U1014_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1015 (
    .in(in[2]),
    .clk(clk),
    .out(_U1015_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1016 (
    .in(in[3]),
    .clk(clk),
    .out(_U1016_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1017 (
    .in(in[4]),
    .clk(clk),
    .out(_U1017_out)
);
assign out[4] = _U1017_out;
assign out[3] = _U1016_out;
assign out[2] = _U1015_out;
assign out[1] = _U1014_out;
assign out[0] = _U1013_out;
endmodule

module array_delay_U1005 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1006_out;
wire [15:0] _U1007_out;
wire [15:0] _U1008_out;
wire [15:0] _U1009_out;
wire [15:0] _U1010_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1006 (
    .in(in[0]),
    .clk(clk),
    .out(_U1006_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1007 (
    .in(in[1]),
    .clk(clk),
    .out(_U1007_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1008 (
    .in(in[2]),
    .clk(clk),
    .out(_U1008_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1009 (
    .in(in[3]),
    .clk(clk),
    .out(_U1009_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1010 (
    .in(in[4]),
    .clk(clk),
    .out(_U1010_out)
);
assign out[4] = _U1010_out;
assign out[3] = _U1009_out;
assign out[2] = _U1008_out;
assign out[1] = _U1007_out;
assign out[0] = _U1006_out;
endmodule

module aff__U969 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U968 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire d_4_at_max_out;
wire [15:0] d_4_next_value_out;
wire [15:0] d_4_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [4:0];
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U969 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_next_value_out = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_next_value_out = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_next_value_out = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_next_value_out = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_next_value_out),
    .clk(clk),
    .out(d_4_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U93 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U92 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U93 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U781 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U780 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire d_4_at_max_out;
wire [15:0] d_4_next_value_out;
wire [15:0] d_4_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [4:0];
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U781 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_next_value_out = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_next_value_out = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_next_value_out = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_next_value_out = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_next_value_out),
    .clk(clk),
    .out(d_4_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U70 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U69 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U70 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U593 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U592 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire d_4_at_max_out;
wire [15:0] d_4_next_value_out;
wire [15:0] d_4_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [4:0];
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U593 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_next_value_out = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_next_value_out = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_next_value_out = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_next_value_out = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_next_value_out),
    .clk(clk),
    .out(d_4_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U47 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U46 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U47 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U405 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U404 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire d_4_at_max_out;
wire [15:0] d_4_next_value_out;
wire [15:0] d_4_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [4:0];
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U405 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_next_value_out = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_next_value_out = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_next_value_out = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_next_value_out = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_next_value_out),
    .clk(clk),
    .out(d_4_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U382 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U381 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U382 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U359 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U358 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U359 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U336 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U335 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U336 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U313 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U312 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U313 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U290 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U289 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U290 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U267 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U266 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U267 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U244 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U243 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U244 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U24 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U23 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U24 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U2238 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U2237 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U2238 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U221 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U220 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U221 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U2191 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U2190 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U2191 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U2144 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U2143 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U2144 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U2097 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U2096 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U2097 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U2050 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U2049 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U2050 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U2003 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U2002 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U2003 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1956 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U1955 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1956 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1909 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U1908 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1909 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U185 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h00d8 * d[1])))) + (16'(16'h0048 * d[2])))) + (16'(16'h0009 * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h0002);
endmodule

module affine_controller__U184 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire d_4_at_max_out;
wire [15:0] d_4_next_value_out;
wire [15:0] d_4_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [4:0];
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U185 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_next_value_out = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_next_value_out = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h0007;
assign d_3_next_value_out = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign d_4_at_max_out = d_4_reg_out == 16'h0007;
assign d_4_next_value_out = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_next_value_out),
    .clk(clk),
    .out(d_4_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1721 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U1720 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire d_4_at_max_out;
wire [15:0] d_4_next_value_out;
wire [15:0] d_4_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [4:0];
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1721 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_next_value_out = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_next_value_out = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_next_value_out = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_next_value_out = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_next_value_out),
    .clk(clk),
    .out(d_4_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U162 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U161 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U162 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1533 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U1532 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire d_4_at_max_out;
wire [15:0] d_4_next_value_out;
wire [15:0] d_4_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [4:0];
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1533 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_next_value_out = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_next_value_out = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_next_value_out = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_next_value_out = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_next_value_out),
    .clk(clk),
    .out(d_4_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U139 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U138 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U139 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1345 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U1344 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire d_4_at_max_out;
wire [15:0] d_4_next_value_out;
wire [15:0] d_4_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [4:0];
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1345 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_next_value_out = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_next_value_out = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_next_value_out = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_next_value_out = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_next_value_out),
    .clk(clk),
    .out(d_4_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U116 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U115 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U116 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1157 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U1156 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire d_4_at_max_out;
wire [15:0] d_4_next_value_out;
wire [15:0] d_4_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [4:0];
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1157 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_next_value_out = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_next_value_out = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_next_value_out = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_next_value_out = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_next_value_out),
    .clk(clk),
    .out(d_4_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U0 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module _U997_pt__U998 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U990_pt__U991 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U987_pt__U988 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U973_pt__U974 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U965_pt__U966 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U961_pt__U962 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U95_pt__U96 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U957_pt__U958 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U949_pt__U950 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U946_pt__U947 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U938_pt__U939 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U932_pt__U933 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U917_pt__U918 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U914_pt__U915 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U905_pt__U906 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U902_pt__U903 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U8_pt__U9 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_4_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
_U8_pt__U9 _U8 (
    .in(in0_hw_input_stencil[0]),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil_4 (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read[0];
hcompute_hw_input_global_wrapper_stencil_4_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U899_pt__U900 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U891_pt__U892 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U888_pt__U889 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U885_pt__U886 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U882_pt__U883 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U876_pt__U877 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U86_pt__U87 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U864_pt__U865 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U859_pt__U860 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U856_pt__U857 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U840_pt__U841 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U838_pt__U839 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U831_pt__U832 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U824_pt__U825 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U818_pt__U819 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U812_pt__U813 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U807_pt__U808 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U802_pt__U803 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U798_pt__U799 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U794_pt__U795 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U791_pt__U792 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U78_pt__U79 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U788_pt__U789 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U786_pt__U787 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U784_pt__U785 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U768_pt__U769 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U765_pt__U766 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U761_pt__U762 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U758_pt__U759 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U752_pt__U753 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U749_pt__U750 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U741_pt__U742 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U738_pt__U739 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U728_pt__U729 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U725_pt__U726 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U713_pt__U714 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U710_pt__U711 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U70_pt__U71 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U707_pt__U708 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U6_pt__U7 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_3_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
_U6_pt__U7 _U6 (
    .in(in0_hw_input_stencil[0]),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil_3 (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read[0];
hcompute_hw_input_global_wrapper_stencil_3_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U693_pt__U694 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U691_pt__U692 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U688_pt__U689 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U671_pt__U672 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U663_pt__U664 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U654_pt__U655 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U646_pt__U647 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U63_pt__U64 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U637_pt__U638 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_11_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U637_out;
wire [15:0] _U639_out;
wire [15:0] _U640_out;
wire [15:0] _U641_out;
wire [15:0] _U642_out;
wire [15:0] _U643_out;
wire [15:0] _U644_out;
wire [15:0] _U645_out;
wire [15:0] _U646_out;
wire [15:0] _U648_out;
wire [15:0] _U649_out;
wire [15:0] _U650_out;
wire [15:0] _U651_out;
wire [15:0] _U652_out;
wire [15:0] _U653_out;
wire [15:0] _U654_out;
wire [15:0] _U656_out;
wire [15:0] _U657_out;
wire [15:0] _U658_out;
wire [15:0] _U659_out;
wire [15:0] _U660_out;
wire [15:0] _U661_out;
wire [15:0] _U662_out;
wire [15:0] _U663_out;
wire [15:0] _U665_out;
wire [15:0] _U666_out;
wire [15:0] _U667_out;
wire [15:0] _U668_out;
wire [15:0] _U669_out;
wire [15:0] _U670_out;
wire [15:0] _U671_out;
wire [15:0] _U673_out;
wire [15:0] _U674_out;
wire [15:0] _U675_out;
wire [15:0] _U676_out;
wire [15:0] _U677_out;
wire [15:0] _U678_out;
wire [15:0] _U679_out;
wire [15:0] _U680_out;
wire [15:0] _U681_out;
wire [15:0] _U682_out;
wire [15:0] _U683_out;
wire [15:0] _U684_out;
wire [15:0] _U685_out;
wire [15:0] _U686_out;
wire [15:0] _U687_out;
wire [15:0] _U688_out;
wire [15:0] _U690_out;
wire [15:0] _U693_out;
wire [15:0] _U695_out;
wire [15:0] _U696_out;
wire [15:0] _U697_out;
wire [15:0] _U698_out;
wire [15:0] _U699_out;
wire [15:0] _U700_out;
wire [15:0] _U701_out;
wire [15:0] _U702_out;
wire [15:0] _U703_out;
wire [15:0] _U704_out;
wire [15:0] _U705_out;
wire [15:0] _U706_out;
wire [15:0] _U707_out;
wire [15:0] _U709_out;
wire [15:0] _U710_out;
wire [15:0] _U712_out;
wire [15:0] _U713_out;
wire [15:0] _U715_out;
wire [15:0] _U716_out;
wire [15:0] _U717_out;
wire [15:0] _U718_out;
wire [15:0] _U719_out;
wire [15:0] _U720_out;
wire [15:0] _U721_out;
wire [15:0] _U722_out;
wire [15:0] _U723_out;
wire [15:0] _U724_out;
wire [15:0] _U725_out;
wire [15:0] _U727_out;
wire [15:0] _U728_out;
wire [15:0] _U730_out;
wire [15:0] _U731_out;
wire [15:0] _U732_out;
wire [15:0] _U733_out;
wire [15:0] _U734_out;
wire [15:0] _U735_out;
wire [15:0] _U736_out;
wire [15:0] _U737_out;
wire [15:0] _U738_out;
wire [15:0] _U740_out;
wire [15:0] _U741_out;
wire [15:0] _U743_out;
wire [15:0] _U744_out;
wire [15:0] _U745_out;
wire [15:0] _U746_out;
wire [15:0] _U747_out;
wire [15:0] _U748_out;
wire [15:0] _U749_out;
wire [15:0] _U751_out;
wire [15:0] _U752_out;
wire [15:0] _U754_out;
wire [15:0] _U755_out;
wire [15:0] _U756_out;
wire [15:0] _U757_out;
wire [15:0] _U758_out;
wire [15:0] _U760_out;
wire [15:0] _U761_out;
wire [15:0] _U763_out;
wire [15:0] _U764_out;
wire [15:0] _U765_out;
wire [15:0] _U767_out;
wire [15:0] _U768_out;
wire [15:0] _U770_out;
wire [15:0] _U771_out;
wire [15:0] _U772_out;
wire [15:0] _U773_out;
wire [15:0] _U774_out;
wire [15:0] _U775_out;
wire [15:0] _U776_out;
wire [15:0] _U777_out;
wire [15:0] _U778_out;
wire [15:0] _U779_out;
wire [15:0] _U780_out;
wire [15:0] _U781_out;
wire [15:0] _U782_out;
wire [15:0] _U783_out;
wire [15:0] _U784_out;
wire [15:0] _U786_out;
wire [15:0] _U788_out;
wire [15:0] _U790_out;
wire [15:0] _U791_out;
wire [15:0] _U793_out;
wire [15:0] _U794_out;
wire [15:0] _U796_out;
wire [15:0] _U797_out;
wire [15:0] _U798_out;
wire [15:0] _U800_out;
wire [15:0] _U801_out;
wire [15:0] _U802_out;
wire [15:0] _U804_out;
wire [15:0] _U805_out;
wire [15:0] _U806_out;
wire [15:0] _U807_out;
wire [15:0] _U809_out;
wire [15:0] _U810_out;
wire [15:0] _U811_out;
wire [15:0] _U812_out;
wire [15:0] _U814_out;
wire [15:0] _U815_out;
wire [15:0] _U816_out;
wire [15:0] _U817_out;
wire [15:0] _U818_out;
wire [15:0] _U820_out;
wire [15:0] _U821_out;
wire [15:0] _U822_out;
wire [15:0] _U823_out;
wire [15:0] _U824_out;
wire [15:0] _U826_out;
wire [15:0] _U827_out;
wire [15:0] _U828_out;
wire [15:0] _U829_out;
wire [15:0] _U830_out;
wire [15:0] _U831_out;
wire [15:0] _U833_out;
wire [15:0] _U834_out;
wire [15:0] _U835_out;
wire [15:0] _U836_out;
wire [15:0] _U837_out;
wire [15:0] add_919_933_934_out;
wire [15:0] add_920_931_932_out;
wire [15:0] add_921_930_931_out;
wire [15:0] add_922_929_930_out;
wire [15:0] add_923_928_929_out;
wire [15:0] add_924_927_928_out;
wire [15:0] add_925_926_927_out;
wire [15:0] add_conv_stencil_4_932_933_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_25_hw_input_global_wrapper_stencil_25_919_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_26_hw_input_global_wrapper_stencil_26_920_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_27_hw_input_global_wrapper_stencil_27_921_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_28_hw_input_global_wrapper_stencil_28_922_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_29_hw_input_global_wrapper_stencil_29_923_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_30_hw_input_global_wrapper_stencil_30_924_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_31_hw_input_global_wrapper_stencil_31_925_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_32_hw_input_global_wrapper_stencil_32_926_out;
_U637_pt__U638 _U637 (
    .in(_U645_out),
    .out(_U637_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U639 (
    .in(in2_hw_kernel_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U639_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U640 (
    .in(_U639_out),
    .clk(clk),
    .out(_U640_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U641 (
    .in(_U640_out),
    .clk(clk),
    .out(_U641_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U642 (
    .in(_U641_out),
    .clk(clk),
    .out(_U642_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U643 (
    .in(_U642_out),
    .clk(clk),
    .out(_U643_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U644 (
    .in(_U643_out),
    .clk(clk),
    .out(_U644_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U645 (
    .in(_U644_out),
    .clk(clk),
    .out(_U645_out)
);
_U646_pt__U647 _U646 (
    .in(_U653_out),
    .out(_U646_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U648 (
    .in(in2_hw_kernel_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U648_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U649 (
    .in(_U648_out),
    .clk(clk),
    .out(_U649_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U650 (
    .in(_U649_out),
    .clk(clk),
    .out(_U650_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U651 (
    .in(_U650_out),
    .clk(clk),
    .out(_U651_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U652 (
    .in(_U651_out),
    .clk(clk),
    .out(_U652_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U653 (
    .in(_U652_out),
    .clk(clk),
    .out(_U653_out)
);
_U654_pt__U655 _U654 (
    .in(_U662_out),
    .out(_U654_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U656 (
    .in(in1_hw_input_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U656_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U657 (
    .in(_U656_out),
    .clk(clk),
    .out(_U657_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U658 (
    .in(_U657_out),
    .clk(clk),
    .out(_U658_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U659 (
    .in(_U658_out),
    .clk(clk),
    .out(_U659_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U660 (
    .in(_U659_out),
    .clk(clk),
    .out(_U660_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U661 (
    .in(_U660_out),
    .clk(clk),
    .out(_U661_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U662 (
    .in(_U661_out),
    .clk(clk),
    .out(_U662_out)
);
_U663_pt__U664 _U663 (
    .in(_U670_out),
    .out(_U663_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U665 (
    .in(in1_hw_input_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U665_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U666 (
    .in(_U665_out),
    .clk(clk),
    .out(_U666_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U667 (
    .in(_U666_out),
    .clk(clk),
    .out(_U667_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U668 (
    .in(_U667_out),
    .clk(clk),
    .out(_U668_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U669 (
    .in(_U668_out),
    .clk(clk),
    .out(_U669_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U670 (
    .in(_U669_out),
    .clk(clk),
    .out(_U670_out)
);
_U671_pt__U672 _U671 (
    .in(_U687_out),
    .out(_U671_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U673 (
    .in(mul_hw_kernel_global_wrapper_stencil_25_hw_input_global_wrapper_stencil_25_919_out),
    .clk(clk),
    .out(_U673_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U674 (
    .in(_U673_out),
    .clk(clk),
    .out(_U674_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U675 (
    .in(_U674_out),
    .clk(clk),
    .out(_U675_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U676 (
    .in(_U675_out),
    .clk(clk),
    .out(_U676_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U677 (
    .in(_U676_out),
    .clk(clk),
    .out(_U677_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U678 (
    .in(_U677_out),
    .clk(clk),
    .out(_U678_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U679 (
    .in(_U678_out),
    .clk(clk),
    .out(_U679_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U680 (
    .in(_U679_out),
    .clk(clk),
    .out(_U680_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U681 (
    .in(_U680_out),
    .clk(clk),
    .out(_U681_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U682 (
    .in(_U681_out),
    .clk(clk),
    .out(_U682_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U683 (
    .in(_U682_out),
    .clk(clk),
    .out(_U683_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U684 (
    .in(_U683_out),
    .clk(clk),
    .out(_U684_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U685 (
    .in(_U684_out),
    .clk(clk),
    .out(_U685_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U686 (
    .in(_U685_out),
    .clk(clk),
    .out(_U686_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U687 (
    .in(_U686_out),
    .clk(clk),
    .out(_U687_out)
);
_U688_pt__U689 _U688 (
    .in(_U690_out),
    .out(_U688_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U690 (
    .in(add_conv_stencil_4_932_933_out),
    .clk(clk),
    .out(_U690_out)
);
_U691_pt__U692 _U691 (
    .in(add_919_933_934_out),
    .out(out_conv_stencil)
);
_U693_pt__U694 _U693 (
    .in(_U706_out),
    .out(_U693_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U695 (
    .in(mul_hw_kernel_global_wrapper_stencil_26_hw_input_global_wrapper_stencil_26_920_out),
    .clk(clk),
    .out(_U695_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U696 (
    .in(_U695_out),
    .clk(clk),
    .out(_U696_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U697 (
    .in(_U696_out),
    .clk(clk),
    .out(_U697_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U698 (
    .in(_U697_out),
    .clk(clk),
    .out(_U698_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U699 (
    .in(_U698_out),
    .clk(clk),
    .out(_U699_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U700 (
    .in(_U699_out),
    .clk(clk),
    .out(_U700_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U701 (
    .in(_U700_out),
    .clk(clk),
    .out(_U701_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U702 (
    .in(_U701_out),
    .clk(clk),
    .out(_U702_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U703 (
    .in(_U702_out),
    .clk(clk),
    .out(_U703_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U704 (
    .in(_U703_out),
    .clk(clk),
    .out(_U704_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U705 (
    .in(_U704_out),
    .clk(clk),
    .out(_U705_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U706 (
    .in(_U705_out),
    .clk(clk),
    .out(_U706_out)
);
_U707_pt__U708 _U707 (
    .in(_U709_out),
    .out(_U707_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U709 (
    .in(add_921_930_931_out),
    .clk(clk),
    .out(_U709_out)
);
_U710_pt__U711 _U710 (
    .in(_U712_out),
    .out(_U710_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U712 (
    .in(add_920_931_932_out),
    .clk(clk),
    .out(_U712_out)
);
_U713_pt__U714 _U713 (
    .in(_U724_out),
    .out(_U713_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U715 (
    .in(mul_hw_kernel_global_wrapper_stencil_27_hw_input_global_wrapper_stencil_27_921_out),
    .clk(clk),
    .out(_U715_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U716 (
    .in(_U715_out),
    .clk(clk),
    .out(_U716_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U717 (
    .in(_U716_out),
    .clk(clk),
    .out(_U717_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U718 (
    .in(_U717_out),
    .clk(clk),
    .out(_U718_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U719 (
    .in(_U718_out),
    .clk(clk),
    .out(_U719_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U720 (
    .in(_U719_out),
    .clk(clk),
    .out(_U720_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U721 (
    .in(_U720_out),
    .clk(clk),
    .out(_U721_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U722 (
    .in(_U721_out),
    .clk(clk),
    .out(_U722_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U723 (
    .in(_U722_out),
    .clk(clk),
    .out(_U723_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U724 (
    .in(_U723_out),
    .clk(clk),
    .out(_U724_out)
);
_U725_pt__U726 _U725 (
    .in(_U727_out),
    .out(_U725_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U727 (
    .in(add_922_929_930_out),
    .clk(clk),
    .out(_U727_out)
);
_U728_pt__U729 _U728 (
    .in(_U737_out),
    .out(_U728_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U730 (
    .in(mul_hw_kernel_global_wrapper_stencil_28_hw_input_global_wrapper_stencil_28_922_out),
    .clk(clk),
    .out(_U730_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U731 (
    .in(_U730_out),
    .clk(clk),
    .out(_U731_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U732 (
    .in(_U731_out),
    .clk(clk),
    .out(_U732_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U733 (
    .in(_U732_out),
    .clk(clk),
    .out(_U733_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U734 (
    .in(_U733_out),
    .clk(clk),
    .out(_U734_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U735 (
    .in(_U734_out),
    .clk(clk),
    .out(_U735_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U736 (
    .in(_U735_out),
    .clk(clk),
    .out(_U736_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U737 (
    .in(_U736_out),
    .clk(clk),
    .out(_U737_out)
);
_U738_pt__U739 _U738 (
    .in(_U740_out),
    .out(_U738_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U740 (
    .in(add_923_928_929_out),
    .clk(clk),
    .out(_U740_out)
);
_U741_pt__U742 _U741 (
    .in(_U748_out),
    .out(_U741_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U743 (
    .in(mul_hw_kernel_global_wrapper_stencil_29_hw_input_global_wrapper_stencil_29_923_out),
    .clk(clk),
    .out(_U743_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U744 (
    .in(_U743_out),
    .clk(clk),
    .out(_U744_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U745 (
    .in(_U744_out),
    .clk(clk),
    .out(_U745_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U746 (
    .in(_U745_out),
    .clk(clk),
    .out(_U746_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U747 (
    .in(_U746_out),
    .clk(clk),
    .out(_U747_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U748 (
    .in(_U747_out),
    .clk(clk),
    .out(_U748_out)
);
_U749_pt__U750 _U749 (
    .in(_U751_out),
    .out(_U749_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U751 (
    .in(add_924_927_928_out),
    .clk(clk),
    .out(_U751_out)
);
_U752_pt__U753 _U752 (
    .in(_U757_out),
    .out(_U752_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U754 (
    .in(mul_hw_kernel_global_wrapper_stencil_30_hw_input_global_wrapper_stencil_30_924_out),
    .clk(clk),
    .out(_U754_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U755 (
    .in(_U754_out),
    .clk(clk),
    .out(_U755_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U756 (
    .in(_U755_out),
    .clk(clk),
    .out(_U756_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U757 (
    .in(_U756_out),
    .clk(clk),
    .out(_U757_out)
);
_U758_pt__U759 _U758 (
    .in(_U760_out),
    .out(_U758_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U760 (
    .in(add_925_926_927_out),
    .clk(clk),
    .out(_U760_out)
);
_U761_pt__U762 _U761 (
    .in(_U764_out),
    .out(_U761_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U763 (
    .in(mul_hw_kernel_global_wrapper_stencil_31_hw_input_global_wrapper_stencil_31_925_out),
    .clk(clk),
    .out(_U763_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U764 (
    .in(_U763_out),
    .clk(clk),
    .out(_U764_out)
);
_U765_pt__U766 _U765 (
    .in(_U767_out),
    .out(_U765_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U767 (
    .in(mul_hw_kernel_global_wrapper_stencil_32_hw_input_global_wrapper_stencil_32_926_out),
    .clk(clk),
    .out(_U767_out)
);
_U768_pt__U769 _U768 (
    .in(_U783_out),
    .out(_U768_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U770 (
    .in(in0_conv_stencil[0]),
    .clk(clk),
    .out(_U770_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U771 (
    .in(_U770_out),
    .clk(clk),
    .out(_U771_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U772 (
    .in(_U771_out),
    .clk(clk),
    .out(_U772_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U773 (
    .in(_U772_out),
    .clk(clk),
    .out(_U773_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U774 (
    .in(_U773_out),
    .clk(clk),
    .out(_U774_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U775 (
    .in(_U774_out),
    .clk(clk),
    .out(_U775_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U776 (
    .in(_U775_out),
    .clk(clk),
    .out(_U776_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U777 (
    .in(_U776_out),
    .clk(clk),
    .out(_U777_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U778 (
    .in(_U777_out),
    .clk(clk),
    .out(_U778_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U779 (
    .in(_U778_out),
    .clk(clk),
    .out(_U779_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U780 (
    .in(_U779_out),
    .clk(clk),
    .out(_U780_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U781 (
    .in(_U780_out),
    .clk(clk),
    .out(_U781_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U782 (
    .in(_U781_out),
    .clk(clk),
    .out(_U782_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U783 (
    .in(_U782_out),
    .clk(clk),
    .out(_U783_out)
);
_U784_pt__U785 _U784 (
    .in(in2_hw_kernel_global_wrapper_stencil[0]),
    .out(_U784_out)
);
_U786_pt__U787 _U786 (
    .in(in1_hw_input_global_wrapper_stencil[0]),
    .out(_U786_out)
);
_U788_pt__U789 _U788 (
    .in(_U790_out),
    .out(_U788_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U790 (
    .in(in2_hw_kernel_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U790_out)
);
_U791_pt__U792 _U791 (
    .in(_U793_out),
    .out(_U791_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U793 (
    .in(in1_hw_input_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U793_out)
);
_U794_pt__U795 _U794 (
    .in(_U797_out),
    .out(_U794_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U796 (
    .in(in2_hw_kernel_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U796_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U797 (
    .in(_U796_out),
    .clk(clk),
    .out(_U797_out)
);
_U798_pt__U799 _U798 (
    .in(_U801_out),
    .out(_U798_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U800 (
    .in(in1_hw_input_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U800_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U801 (
    .in(_U800_out),
    .clk(clk),
    .out(_U801_out)
);
_U802_pt__U803 _U802 (
    .in(_U806_out),
    .out(_U802_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U804 (
    .in(in2_hw_kernel_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U804_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U805 (
    .in(_U804_out),
    .clk(clk),
    .out(_U805_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U806 (
    .in(_U805_out),
    .clk(clk),
    .out(_U806_out)
);
_U807_pt__U808 _U807 (
    .in(_U811_out),
    .out(_U807_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U809 (
    .in(in1_hw_input_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U809_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U810 (
    .in(_U809_out),
    .clk(clk),
    .out(_U810_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U811 (
    .in(_U810_out),
    .clk(clk),
    .out(_U811_out)
);
_U812_pt__U813 _U812 (
    .in(_U817_out),
    .out(_U812_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U814 (
    .in(in2_hw_kernel_global_wrapper_stencil[4]),
    .clk(clk),
    .out(_U814_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U815 (
    .in(_U814_out),
    .clk(clk),
    .out(_U815_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U816 (
    .in(_U815_out),
    .clk(clk),
    .out(_U816_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U817 (
    .in(_U816_out),
    .clk(clk),
    .out(_U817_out)
);
_U818_pt__U819 _U818 (
    .in(_U823_out),
    .out(_U818_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U820 (
    .in(in1_hw_input_global_wrapper_stencil[4]),
    .clk(clk),
    .out(_U820_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U821 (
    .in(_U820_out),
    .clk(clk),
    .out(_U821_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U822 (
    .in(_U821_out),
    .clk(clk),
    .out(_U822_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U823 (
    .in(_U822_out),
    .clk(clk),
    .out(_U823_out)
);
_U824_pt__U825 _U824 (
    .in(_U830_out),
    .out(_U824_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U826 (
    .in(in2_hw_kernel_global_wrapper_stencil[5]),
    .clk(clk),
    .out(_U826_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U827 (
    .in(_U826_out),
    .clk(clk),
    .out(_U827_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U828 (
    .in(_U827_out),
    .clk(clk),
    .out(_U828_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U829 (
    .in(_U828_out),
    .clk(clk),
    .out(_U829_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U830 (
    .in(_U829_out),
    .clk(clk),
    .out(_U830_out)
);
_U831_pt__U832 _U831 (
    .in(_U837_out),
    .out(_U831_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U833 (
    .in(in1_hw_input_global_wrapper_stencil[5]),
    .clk(clk),
    .out(_U833_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U834 (
    .in(_U833_out),
    .clk(clk),
    .out(_U834_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U835 (
    .in(_U834_out),
    .clk(clk),
    .out(_U835_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U836 (
    .in(_U835_out),
    .clk(clk),
    .out(_U836_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U837 (
    .in(_U836_out),
    .clk(clk),
    .out(_U837_out)
);
assign add_919_933_934_out = 16'(_U671_out + _U688_out);
assign add_920_931_932_out = 16'(_U693_out + _U707_out);
assign add_921_930_931_out = 16'(_U713_out + _U725_out);
assign add_922_929_930_out = 16'(_U728_out + _U738_out);
assign add_923_928_929_out = 16'(_U741_out + _U749_out);
assign add_924_927_928_out = 16'(_U752_out + _U758_out);
assign add_925_926_927_out = 16'(_U761_out + _U765_out);
assign add_conv_stencil_4_932_933_out = 16'(_U768_out + _U710_out);
assign mul_hw_kernel_global_wrapper_stencil_25_hw_input_global_wrapper_stencil_25_919_out = 16'(_U784_out * _U786_out);
assign mul_hw_kernel_global_wrapper_stencil_26_hw_input_global_wrapper_stencil_26_920_out = 16'(_U788_out * _U791_out);
assign mul_hw_kernel_global_wrapper_stencil_27_hw_input_global_wrapper_stencil_27_921_out = 16'(_U794_out * _U798_out);
assign mul_hw_kernel_global_wrapper_stencil_28_hw_input_global_wrapper_stencil_28_922_out = 16'(_U802_out * _U807_out);
assign mul_hw_kernel_global_wrapper_stencil_29_hw_input_global_wrapper_stencil_29_923_out = 16'(_U812_out * _U818_out);
assign mul_hw_kernel_global_wrapper_stencil_30_hw_input_global_wrapper_stencil_30_924_out = 16'(_U824_out * _U831_out);
assign mul_hw_kernel_global_wrapper_stencil_31_hw_input_global_wrapper_stencil_31_925_out = 16'(_U646_out * _U663_out);
assign mul_hw_kernel_global_wrapper_stencil_32_hw_input_global_wrapper_stencil_32_926_out = 16'(_U637_out * _U654_out);
endmodule

module cu_op_hcompute_conv_stencil_11 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_11_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_11_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_11_read[0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[0];
hcompute_conv_stencil_11_pipelined inner_compute (
    .clk(clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_11_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U628_pt__U629 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U619_pt__U620 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U611_pt__U612 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U603_pt__U604 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U596_pt__U597 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U589_pt__U590 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U583_pt__U584 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U577_pt__U578 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U572_pt__U573 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U56_pt__U57 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U567_pt__U568 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U563_pt__U564 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U559_pt__U560 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U556_pt__U557 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U553_pt__U554 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U551_pt__U552 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U549_pt__U550 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U533_pt__U534 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U530_pt__U531 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U526_pt__U527 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U523_pt__U524 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U517_pt__U518 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U514_pt__U515 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U50_pt__U51 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U506_pt__U507 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U503_pt__U504 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U4_pt__U5 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_2_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
_U4_pt__U5 _U4 (
    .in(in0_hw_input_stencil[0]),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil_2 (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read[0];
hcompute_hw_input_global_wrapper_stencil_2_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U493_pt__U494 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U490_pt__U491 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U478_pt__U479 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U475_pt__U476 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U472_pt__U473 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U458_pt__U459 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U456_pt__U457 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U453_pt__U454 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U44_pt__U45 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U436_pt__U437 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_10_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U436_out;
wire [15:0] _U438_out;
wire [15:0] _U439_out;
wire [15:0] _U440_out;
wire [15:0] _U441_out;
wire [15:0] _U442_out;
wire [15:0] _U443_out;
wire [15:0] _U444_out;
wire [15:0] _U445_out;
wire [15:0] _U446_out;
wire [15:0] _U447_out;
wire [15:0] _U448_out;
wire [15:0] _U449_out;
wire [15:0] _U450_out;
wire [15:0] _U451_out;
wire [15:0] _U452_out;
wire [15:0] _U453_out;
wire [15:0] _U455_out;
wire [15:0] _U458_out;
wire [15:0] _U460_out;
wire [15:0] _U461_out;
wire [15:0] _U462_out;
wire [15:0] _U463_out;
wire [15:0] _U464_out;
wire [15:0] _U465_out;
wire [15:0] _U466_out;
wire [15:0] _U467_out;
wire [15:0] _U468_out;
wire [15:0] _U469_out;
wire [15:0] _U470_out;
wire [15:0] _U471_out;
wire [15:0] _U472_out;
wire [15:0] _U474_out;
wire [15:0] _U475_out;
wire [15:0] _U477_out;
wire [15:0] _U478_out;
wire [15:0] _U480_out;
wire [15:0] _U481_out;
wire [15:0] _U482_out;
wire [15:0] _U483_out;
wire [15:0] _U484_out;
wire [15:0] _U485_out;
wire [15:0] _U486_out;
wire [15:0] _U487_out;
wire [15:0] _U488_out;
wire [15:0] _U489_out;
wire [15:0] _U490_out;
wire [15:0] _U492_out;
wire [15:0] _U493_out;
wire [15:0] _U495_out;
wire [15:0] _U496_out;
wire [15:0] _U497_out;
wire [15:0] _U498_out;
wire [15:0] _U499_out;
wire [15:0] _U500_out;
wire [15:0] _U501_out;
wire [15:0] _U502_out;
wire [15:0] _U503_out;
wire [15:0] _U505_out;
wire [15:0] _U506_out;
wire [15:0] _U508_out;
wire [15:0] _U509_out;
wire [15:0] _U510_out;
wire [15:0] _U511_out;
wire [15:0] _U512_out;
wire [15:0] _U513_out;
wire [15:0] _U514_out;
wire [15:0] _U516_out;
wire [15:0] _U517_out;
wire [15:0] _U519_out;
wire [15:0] _U520_out;
wire [15:0] _U521_out;
wire [15:0] _U522_out;
wire [15:0] _U523_out;
wire [15:0] _U525_out;
wire [15:0] _U526_out;
wire [15:0] _U528_out;
wire [15:0] _U529_out;
wire [15:0] _U530_out;
wire [15:0] _U532_out;
wire [15:0] _U533_out;
wire [15:0] _U535_out;
wire [15:0] _U536_out;
wire [15:0] _U537_out;
wire [15:0] _U538_out;
wire [15:0] _U539_out;
wire [15:0] _U540_out;
wire [15:0] _U541_out;
wire [15:0] _U542_out;
wire [15:0] _U543_out;
wire [15:0] _U544_out;
wire [15:0] _U545_out;
wire [15:0] _U546_out;
wire [15:0] _U547_out;
wire [15:0] _U548_out;
wire [15:0] _U549_out;
wire [15:0] _U551_out;
wire [15:0] _U553_out;
wire [15:0] _U555_out;
wire [15:0] _U556_out;
wire [15:0] _U558_out;
wire [15:0] _U559_out;
wire [15:0] _U561_out;
wire [15:0] _U562_out;
wire [15:0] _U563_out;
wire [15:0] _U565_out;
wire [15:0] _U566_out;
wire [15:0] _U567_out;
wire [15:0] _U569_out;
wire [15:0] _U570_out;
wire [15:0] _U571_out;
wire [15:0] _U572_out;
wire [15:0] _U574_out;
wire [15:0] _U575_out;
wire [15:0] _U576_out;
wire [15:0] _U577_out;
wire [15:0] _U579_out;
wire [15:0] _U580_out;
wire [15:0] _U581_out;
wire [15:0] _U582_out;
wire [15:0] _U583_out;
wire [15:0] _U585_out;
wire [15:0] _U586_out;
wire [15:0] _U587_out;
wire [15:0] _U588_out;
wire [15:0] _U589_out;
wire [15:0] _U591_out;
wire [15:0] _U592_out;
wire [15:0] _U593_out;
wire [15:0] _U594_out;
wire [15:0] _U595_out;
wire [15:0] _U596_out;
wire [15:0] _U598_out;
wire [15:0] _U599_out;
wire [15:0] _U600_out;
wire [15:0] _U601_out;
wire [15:0] _U602_out;
wire [15:0] _U603_out;
wire [15:0] _U605_out;
wire [15:0] _U606_out;
wire [15:0] _U607_out;
wire [15:0] _U608_out;
wire [15:0] _U609_out;
wire [15:0] _U610_out;
wire [15:0] _U611_out;
wire [15:0] _U613_out;
wire [15:0] _U614_out;
wire [15:0] _U615_out;
wire [15:0] _U616_out;
wire [15:0] _U617_out;
wire [15:0] _U618_out;
wire [15:0] _U619_out;
wire [15:0] _U621_out;
wire [15:0] _U622_out;
wire [15:0] _U623_out;
wire [15:0] _U624_out;
wire [15:0] _U625_out;
wire [15:0] _U626_out;
wire [15:0] _U627_out;
wire [15:0] _U628_out;
wire [15:0] _U630_out;
wire [15:0] _U631_out;
wire [15:0] _U632_out;
wire [15:0] _U633_out;
wire [15:0] _U634_out;
wire [15:0] _U635_out;
wire [15:0] _U636_out;
wire [15:0] add_852_866_867_out;
wire [15:0] add_853_864_865_out;
wire [15:0] add_854_863_864_out;
wire [15:0] add_855_862_863_out;
wire [15:0] add_856_861_862_out;
wire [15:0] add_857_860_861_out;
wire [15:0] add_858_859_860_out;
wire [15:0] add_conv_stencil_3_865_866_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_17_hw_input_global_wrapper_stencil_17_852_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_18_hw_input_global_wrapper_stencil_18_853_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_19_hw_input_global_wrapper_stencil_19_854_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_20_hw_input_global_wrapper_stencil_20_855_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_21_hw_input_global_wrapper_stencil_21_856_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_22_hw_input_global_wrapper_stencil_22_857_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_23_hw_input_global_wrapper_stencil_23_858_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_24_hw_input_global_wrapper_stencil_24_859_out;
_U436_pt__U437 _U436 (
    .in(_U452_out),
    .out(_U436_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U438 (
    .in(mul_hw_kernel_global_wrapper_stencil_17_hw_input_global_wrapper_stencil_17_852_out),
    .clk(clk),
    .out(_U438_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U439 (
    .in(_U438_out),
    .clk(clk),
    .out(_U439_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U440 (
    .in(_U439_out),
    .clk(clk),
    .out(_U440_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U441 (
    .in(_U440_out),
    .clk(clk),
    .out(_U441_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U442 (
    .in(_U441_out),
    .clk(clk),
    .out(_U442_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U443 (
    .in(_U442_out),
    .clk(clk),
    .out(_U443_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U444 (
    .in(_U443_out),
    .clk(clk),
    .out(_U444_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U445 (
    .in(_U444_out),
    .clk(clk),
    .out(_U445_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U446 (
    .in(_U445_out),
    .clk(clk),
    .out(_U446_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U447 (
    .in(_U446_out),
    .clk(clk),
    .out(_U447_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U448 (
    .in(_U447_out),
    .clk(clk),
    .out(_U448_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U449 (
    .in(_U448_out),
    .clk(clk),
    .out(_U449_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U450 (
    .in(_U449_out),
    .clk(clk),
    .out(_U450_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U451 (
    .in(_U450_out),
    .clk(clk),
    .out(_U451_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U452 (
    .in(_U451_out),
    .clk(clk),
    .out(_U452_out)
);
_U453_pt__U454 _U453 (
    .in(_U455_out),
    .out(_U453_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U455 (
    .in(add_conv_stencil_3_865_866_out),
    .clk(clk),
    .out(_U455_out)
);
_U456_pt__U457 _U456 (
    .in(add_852_866_867_out),
    .out(out_conv_stencil)
);
_U458_pt__U459 _U458 (
    .in(_U471_out),
    .out(_U458_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U460 (
    .in(mul_hw_kernel_global_wrapper_stencil_18_hw_input_global_wrapper_stencil_18_853_out),
    .clk(clk),
    .out(_U460_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U461 (
    .in(_U460_out),
    .clk(clk),
    .out(_U461_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U462 (
    .in(_U461_out),
    .clk(clk),
    .out(_U462_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U463 (
    .in(_U462_out),
    .clk(clk),
    .out(_U463_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U464 (
    .in(_U463_out),
    .clk(clk),
    .out(_U464_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U465 (
    .in(_U464_out),
    .clk(clk),
    .out(_U465_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U466 (
    .in(_U465_out),
    .clk(clk),
    .out(_U466_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U467 (
    .in(_U466_out),
    .clk(clk),
    .out(_U467_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U468 (
    .in(_U467_out),
    .clk(clk),
    .out(_U468_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U469 (
    .in(_U468_out),
    .clk(clk),
    .out(_U469_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U470 (
    .in(_U469_out),
    .clk(clk),
    .out(_U470_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U471 (
    .in(_U470_out),
    .clk(clk),
    .out(_U471_out)
);
_U472_pt__U473 _U472 (
    .in(_U474_out),
    .out(_U472_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U474 (
    .in(add_854_863_864_out),
    .clk(clk),
    .out(_U474_out)
);
_U475_pt__U476 _U475 (
    .in(_U477_out),
    .out(_U475_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U477 (
    .in(add_853_864_865_out),
    .clk(clk),
    .out(_U477_out)
);
_U478_pt__U479 _U478 (
    .in(_U489_out),
    .out(_U478_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U480 (
    .in(mul_hw_kernel_global_wrapper_stencil_19_hw_input_global_wrapper_stencil_19_854_out),
    .clk(clk),
    .out(_U480_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U481 (
    .in(_U480_out),
    .clk(clk),
    .out(_U481_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U482 (
    .in(_U481_out),
    .clk(clk),
    .out(_U482_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U483 (
    .in(_U482_out),
    .clk(clk),
    .out(_U483_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U484 (
    .in(_U483_out),
    .clk(clk),
    .out(_U484_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U485 (
    .in(_U484_out),
    .clk(clk),
    .out(_U485_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U486 (
    .in(_U485_out),
    .clk(clk),
    .out(_U486_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U487 (
    .in(_U486_out),
    .clk(clk),
    .out(_U487_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U488 (
    .in(_U487_out),
    .clk(clk),
    .out(_U488_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U489 (
    .in(_U488_out),
    .clk(clk),
    .out(_U489_out)
);
_U490_pt__U491 _U490 (
    .in(_U492_out),
    .out(_U490_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U492 (
    .in(add_855_862_863_out),
    .clk(clk),
    .out(_U492_out)
);
_U493_pt__U494 _U493 (
    .in(_U502_out),
    .out(_U493_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U495 (
    .in(mul_hw_kernel_global_wrapper_stencil_20_hw_input_global_wrapper_stencil_20_855_out),
    .clk(clk),
    .out(_U495_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U496 (
    .in(_U495_out),
    .clk(clk),
    .out(_U496_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U497 (
    .in(_U496_out),
    .clk(clk),
    .out(_U497_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U498 (
    .in(_U497_out),
    .clk(clk),
    .out(_U498_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U499 (
    .in(_U498_out),
    .clk(clk),
    .out(_U499_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U500 (
    .in(_U499_out),
    .clk(clk),
    .out(_U500_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U501 (
    .in(_U500_out),
    .clk(clk),
    .out(_U501_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U502 (
    .in(_U501_out),
    .clk(clk),
    .out(_U502_out)
);
_U503_pt__U504 _U503 (
    .in(_U505_out),
    .out(_U503_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U505 (
    .in(add_856_861_862_out),
    .clk(clk),
    .out(_U505_out)
);
_U506_pt__U507 _U506 (
    .in(_U513_out),
    .out(_U506_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U508 (
    .in(mul_hw_kernel_global_wrapper_stencil_21_hw_input_global_wrapper_stencil_21_856_out),
    .clk(clk),
    .out(_U508_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U509 (
    .in(_U508_out),
    .clk(clk),
    .out(_U509_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U510 (
    .in(_U509_out),
    .clk(clk),
    .out(_U510_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U511 (
    .in(_U510_out),
    .clk(clk),
    .out(_U511_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U512 (
    .in(_U511_out),
    .clk(clk),
    .out(_U512_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U513 (
    .in(_U512_out),
    .clk(clk),
    .out(_U513_out)
);
_U514_pt__U515 _U514 (
    .in(_U516_out),
    .out(_U514_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U516 (
    .in(add_857_860_861_out),
    .clk(clk),
    .out(_U516_out)
);
_U517_pt__U518 _U517 (
    .in(_U522_out),
    .out(_U517_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U519 (
    .in(mul_hw_kernel_global_wrapper_stencil_22_hw_input_global_wrapper_stencil_22_857_out),
    .clk(clk),
    .out(_U519_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U520 (
    .in(_U519_out),
    .clk(clk),
    .out(_U520_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U521 (
    .in(_U520_out),
    .clk(clk),
    .out(_U521_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U522 (
    .in(_U521_out),
    .clk(clk),
    .out(_U522_out)
);
_U523_pt__U524 _U523 (
    .in(_U525_out),
    .out(_U523_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U525 (
    .in(add_858_859_860_out),
    .clk(clk),
    .out(_U525_out)
);
_U526_pt__U527 _U526 (
    .in(_U529_out),
    .out(_U526_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U528 (
    .in(mul_hw_kernel_global_wrapper_stencil_23_hw_input_global_wrapper_stencil_23_858_out),
    .clk(clk),
    .out(_U528_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U529 (
    .in(_U528_out),
    .clk(clk),
    .out(_U529_out)
);
_U530_pt__U531 _U530 (
    .in(_U532_out),
    .out(_U530_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U532 (
    .in(mul_hw_kernel_global_wrapper_stencil_24_hw_input_global_wrapper_stencil_24_859_out),
    .clk(clk),
    .out(_U532_out)
);
_U533_pt__U534 _U533 (
    .in(_U548_out),
    .out(_U533_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U535 (
    .in(in0_conv_stencil[0]),
    .clk(clk),
    .out(_U535_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U536 (
    .in(_U535_out),
    .clk(clk),
    .out(_U536_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U537 (
    .in(_U536_out),
    .clk(clk),
    .out(_U537_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U538 (
    .in(_U537_out),
    .clk(clk),
    .out(_U538_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U539 (
    .in(_U538_out),
    .clk(clk),
    .out(_U539_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U540 (
    .in(_U539_out),
    .clk(clk),
    .out(_U540_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U541 (
    .in(_U540_out),
    .clk(clk),
    .out(_U541_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U542 (
    .in(_U541_out),
    .clk(clk),
    .out(_U542_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U543 (
    .in(_U542_out),
    .clk(clk),
    .out(_U543_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U544 (
    .in(_U543_out),
    .clk(clk),
    .out(_U544_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U545 (
    .in(_U544_out),
    .clk(clk),
    .out(_U545_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U546 (
    .in(_U545_out),
    .clk(clk),
    .out(_U546_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U547 (
    .in(_U546_out),
    .clk(clk),
    .out(_U547_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U548 (
    .in(_U547_out),
    .clk(clk),
    .out(_U548_out)
);
_U549_pt__U550 _U549 (
    .in(in2_hw_kernel_global_wrapper_stencil[0]),
    .out(_U549_out)
);
_U551_pt__U552 _U551 (
    .in(in1_hw_input_global_wrapper_stencil[0]),
    .out(_U551_out)
);
_U553_pt__U554 _U553 (
    .in(_U555_out),
    .out(_U553_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U555 (
    .in(in2_hw_kernel_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U555_out)
);
_U556_pt__U557 _U556 (
    .in(_U558_out),
    .out(_U556_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U558 (
    .in(in1_hw_input_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U558_out)
);
_U559_pt__U560 _U559 (
    .in(_U562_out),
    .out(_U559_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U561 (
    .in(in2_hw_kernel_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U561_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U562 (
    .in(_U561_out),
    .clk(clk),
    .out(_U562_out)
);
_U563_pt__U564 _U563 (
    .in(_U566_out),
    .out(_U563_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U565 (
    .in(in1_hw_input_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U565_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U566 (
    .in(_U565_out),
    .clk(clk),
    .out(_U566_out)
);
_U567_pt__U568 _U567 (
    .in(_U571_out),
    .out(_U567_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U569 (
    .in(in2_hw_kernel_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U569_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U570 (
    .in(_U569_out),
    .clk(clk),
    .out(_U570_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U571 (
    .in(_U570_out),
    .clk(clk),
    .out(_U571_out)
);
_U572_pt__U573 _U572 (
    .in(_U576_out),
    .out(_U572_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U574 (
    .in(in1_hw_input_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U574_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U575 (
    .in(_U574_out),
    .clk(clk),
    .out(_U575_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U576 (
    .in(_U575_out),
    .clk(clk),
    .out(_U576_out)
);
_U577_pt__U578 _U577 (
    .in(_U582_out),
    .out(_U577_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U579 (
    .in(in2_hw_kernel_global_wrapper_stencil[4]),
    .clk(clk),
    .out(_U579_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U580 (
    .in(_U579_out),
    .clk(clk),
    .out(_U580_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U581 (
    .in(_U580_out),
    .clk(clk),
    .out(_U581_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U582 (
    .in(_U581_out),
    .clk(clk),
    .out(_U582_out)
);
_U583_pt__U584 _U583 (
    .in(_U588_out),
    .out(_U583_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U585 (
    .in(in1_hw_input_global_wrapper_stencil[4]),
    .clk(clk),
    .out(_U585_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U586 (
    .in(_U585_out),
    .clk(clk),
    .out(_U586_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U587 (
    .in(_U586_out),
    .clk(clk),
    .out(_U587_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U588 (
    .in(_U587_out),
    .clk(clk),
    .out(_U588_out)
);
_U589_pt__U590 _U589 (
    .in(_U595_out),
    .out(_U589_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U591 (
    .in(in2_hw_kernel_global_wrapper_stencil[5]),
    .clk(clk),
    .out(_U591_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U592 (
    .in(_U591_out),
    .clk(clk),
    .out(_U592_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U593 (
    .in(_U592_out),
    .clk(clk),
    .out(_U593_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U594 (
    .in(_U593_out),
    .clk(clk),
    .out(_U594_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U595 (
    .in(_U594_out),
    .clk(clk),
    .out(_U595_out)
);
_U596_pt__U597 _U596 (
    .in(_U602_out),
    .out(_U596_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U598 (
    .in(in1_hw_input_global_wrapper_stencil[5]),
    .clk(clk),
    .out(_U598_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U599 (
    .in(_U598_out),
    .clk(clk),
    .out(_U599_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U600 (
    .in(_U599_out),
    .clk(clk),
    .out(_U600_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U601 (
    .in(_U600_out),
    .clk(clk),
    .out(_U601_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U602 (
    .in(_U601_out),
    .clk(clk),
    .out(_U602_out)
);
_U603_pt__U604 _U603 (
    .in(_U610_out),
    .out(_U603_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U605 (
    .in(in2_hw_kernel_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U605_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U606 (
    .in(_U605_out),
    .clk(clk),
    .out(_U606_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U607 (
    .in(_U606_out),
    .clk(clk),
    .out(_U607_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U608 (
    .in(_U607_out),
    .clk(clk),
    .out(_U608_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U609 (
    .in(_U608_out),
    .clk(clk),
    .out(_U609_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U610 (
    .in(_U609_out),
    .clk(clk),
    .out(_U610_out)
);
_U611_pt__U612 _U611 (
    .in(_U618_out),
    .out(_U611_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U613 (
    .in(in1_hw_input_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U613_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U614 (
    .in(_U613_out),
    .clk(clk),
    .out(_U614_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U615 (
    .in(_U614_out),
    .clk(clk),
    .out(_U615_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U616 (
    .in(_U615_out),
    .clk(clk),
    .out(_U616_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U617 (
    .in(_U616_out),
    .clk(clk),
    .out(_U617_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U618 (
    .in(_U617_out),
    .clk(clk),
    .out(_U618_out)
);
_U619_pt__U620 _U619 (
    .in(_U627_out),
    .out(_U619_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U621 (
    .in(in2_hw_kernel_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U621_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U622 (
    .in(_U621_out),
    .clk(clk),
    .out(_U622_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U623 (
    .in(_U622_out),
    .clk(clk),
    .out(_U623_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U624 (
    .in(_U623_out),
    .clk(clk),
    .out(_U624_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U625 (
    .in(_U624_out),
    .clk(clk),
    .out(_U625_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U626 (
    .in(_U625_out),
    .clk(clk),
    .out(_U626_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U627 (
    .in(_U626_out),
    .clk(clk),
    .out(_U627_out)
);
_U628_pt__U629 _U628 (
    .in(_U636_out),
    .out(_U628_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U630 (
    .in(in1_hw_input_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U630_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U631 (
    .in(_U630_out),
    .clk(clk),
    .out(_U631_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U632 (
    .in(_U631_out),
    .clk(clk),
    .out(_U632_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U633 (
    .in(_U632_out),
    .clk(clk),
    .out(_U633_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U634 (
    .in(_U633_out),
    .clk(clk),
    .out(_U634_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U635 (
    .in(_U634_out),
    .clk(clk),
    .out(_U635_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U636 (
    .in(_U635_out),
    .clk(clk),
    .out(_U636_out)
);
assign add_852_866_867_out = 16'(_U436_out + _U453_out);
assign add_853_864_865_out = 16'(_U458_out + _U472_out);
assign add_854_863_864_out = 16'(_U478_out + _U490_out);
assign add_855_862_863_out = 16'(_U493_out + _U503_out);
assign add_856_861_862_out = 16'(_U506_out + _U514_out);
assign add_857_860_861_out = 16'(_U517_out + _U523_out);
assign add_858_859_860_out = 16'(_U526_out + _U530_out);
assign add_conv_stencil_3_865_866_out = 16'(_U533_out + _U475_out);
assign mul_hw_kernel_global_wrapper_stencil_17_hw_input_global_wrapper_stencil_17_852_out = 16'(_U549_out * _U551_out);
assign mul_hw_kernel_global_wrapper_stencil_18_hw_input_global_wrapper_stencil_18_853_out = 16'(_U553_out * _U556_out);
assign mul_hw_kernel_global_wrapper_stencil_19_hw_input_global_wrapper_stencil_19_854_out = 16'(_U559_out * _U563_out);
assign mul_hw_kernel_global_wrapper_stencil_20_hw_input_global_wrapper_stencil_20_855_out = 16'(_U567_out * _U572_out);
assign mul_hw_kernel_global_wrapper_stencil_21_hw_input_global_wrapper_stencil_21_856_out = 16'(_U577_out * _U583_out);
assign mul_hw_kernel_global_wrapper_stencil_22_hw_input_global_wrapper_stencil_22_857_out = 16'(_U589_out * _U596_out);
assign mul_hw_kernel_global_wrapper_stencil_23_hw_input_global_wrapper_stencil_23_858_out = 16'(_U603_out * _U611_out);
assign mul_hw_kernel_global_wrapper_stencil_24_hw_input_global_wrapper_stencil_24_859_out = 16'(_U619_out * _U628_out);
endmodule

module cu_op_hcompute_conv_stencil_10 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_10_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_10_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_10_read[0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[0];
hcompute_conv_stencil_10_pipelined inner_compute (
    .clk(clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_10_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U425_pt__U426 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U422_pt__U423 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U409_pt__U410 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U406_pt__U407 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U403_pt__U404 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U39_pt__U40 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U388_pt__U389 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U386_pt__U387 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U383_pt__U384 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U373_pt__U374 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U369_pt__U370 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U366_pt__U367 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U363_pt__U364 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U361_pt__U362 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U359_pt__U360 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U34_pt__U35 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U343_pt__U344 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U339_pt__U340 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U334_pt__U335 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U331_pt__U332 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U32_pt__U33 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_7_pipelined (
    output [15:0] out_conv_stencil
);
_U32_pt__U33 _U32 (
    .in(16'h0000),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_7 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_7_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_7_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_7_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U324_pt__U325 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U321_pt__U322 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U312_pt__U313 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U30_pt__U31 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_6_pipelined (
    output [15:0] out_conv_stencil
);
_U30_pt__U31 _U30 (
    .in(16'h0000),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_6 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_6_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_6_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_6_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U309_pt__U310 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U300_pt__U301 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U2_pt__U3 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_1_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
_U2_pt__U3 _U2 (
    .in(in0_hw_input_stencil[0]),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil_1 (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read[0];
hcompute_hw_input_global_wrapper_stencil_1_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U291_pt__U292 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U28_pt__U29 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_5_pipelined (
    output [15:0] out_conv_stencil
);
_U28_pt__U29 _U28 (
    .in(16'h0000),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_5 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_5_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U283_pt__U284 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U275_pt__U276 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U26_pt__U27 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_4_pipelined (
    output [15:0] out_conv_stencil
);
_U26_pt__U27 _U26 (
    .in(16'h0000),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_4 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_4_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U268_pt__U269 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U261_pt__U262 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U255_pt__U256 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U24_pt__U25 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_3_pipelined (
    output [15:0] out_conv_stencil
);
_U24_pt__U25 _U24 (
    .in(16'h0000),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_3 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_3_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U249_pt__U250 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U244_pt__U245 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U239_pt__U240 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U235_pt__U236 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_9_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U235_out;
wire [15:0] _U237_out;
wire [15:0] _U238_out;
wire [15:0] _U239_out;
wire [15:0] _U241_out;
wire [15:0] _U242_out;
wire [15:0] _U243_out;
wire [15:0] _U244_out;
wire [15:0] _U246_out;
wire [15:0] _U247_out;
wire [15:0] _U248_out;
wire [15:0] _U249_out;
wire [15:0] _U251_out;
wire [15:0] _U252_out;
wire [15:0] _U253_out;
wire [15:0] _U254_out;
wire [15:0] _U255_out;
wire [15:0] _U257_out;
wire [15:0] _U258_out;
wire [15:0] _U259_out;
wire [15:0] _U260_out;
wire [15:0] _U261_out;
wire [15:0] _U263_out;
wire [15:0] _U264_out;
wire [15:0] _U265_out;
wire [15:0] _U266_out;
wire [15:0] _U267_out;
wire [15:0] _U268_out;
wire [15:0] _U270_out;
wire [15:0] _U271_out;
wire [15:0] _U272_out;
wire [15:0] _U273_out;
wire [15:0] _U274_out;
wire [15:0] _U275_out;
wire [15:0] _U277_out;
wire [15:0] _U278_out;
wire [15:0] _U279_out;
wire [15:0] _U280_out;
wire [15:0] _U281_out;
wire [15:0] _U282_out;
wire [15:0] _U283_out;
wire [15:0] _U285_out;
wire [15:0] _U286_out;
wire [15:0] _U287_out;
wire [15:0] _U288_out;
wire [15:0] _U289_out;
wire [15:0] _U290_out;
wire [15:0] _U291_out;
wire [15:0] _U293_out;
wire [15:0] _U294_out;
wire [15:0] _U295_out;
wire [15:0] _U296_out;
wire [15:0] _U297_out;
wire [15:0] _U298_out;
wire [15:0] _U299_out;
wire [15:0] _U300_out;
wire [15:0] _U302_out;
wire [15:0] _U303_out;
wire [15:0] _U304_out;
wire [15:0] _U305_out;
wire [15:0] _U306_out;
wire [15:0] _U307_out;
wire [15:0] _U308_out;
wire [15:0] _U309_out;
wire [15:0] _U311_out;
wire [15:0] _U312_out;
wire [15:0] _U314_out;
wire [15:0] _U315_out;
wire [15:0] _U316_out;
wire [15:0] _U317_out;
wire [15:0] _U318_out;
wire [15:0] _U319_out;
wire [15:0] _U320_out;
wire [15:0] _U321_out;
wire [15:0] _U323_out;
wire [15:0] _U324_out;
wire [15:0] _U326_out;
wire [15:0] _U327_out;
wire [15:0] _U328_out;
wire [15:0] _U329_out;
wire [15:0] _U330_out;
wire [15:0] _U331_out;
wire [15:0] _U333_out;
wire [15:0] _U334_out;
wire [15:0] _U336_out;
wire [15:0] _U337_out;
wire [15:0] _U338_out;
wire [15:0] _U339_out;
wire [15:0] _U341_out;
wire [15:0] _U342_out;
wire [15:0] _U343_out;
wire [15:0] _U345_out;
wire [15:0] _U346_out;
wire [15:0] _U347_out;
wire [15:0] _U348_out;
wire [15:0] _U349_out;
wire [15:0] _U350_out;
wire [15:0] _U351_out;
wire [15:0] _U352_out;
wire [15:0] _U353_out;
wire [15:0] _U354_out;
wire [15:0] _U355_out;
wire [15:0] _U356_out;
wire [15:0] _U357_out;
wire [15:0] _U358_out;
wire [15:0] _U359_out;
wire [15:0] _U361_out;
wire [15:0] _U363_out;
wire [15:0] _U365_out;
wire [15:0] _U366_out;
wire [15:0] _U368_out;
wire [15:0] _U369_out;
wire [15:0] _U371_out;
wire [15:0] _U372_out;
wire [15:0] _U373_out;
wire [15:0] _U375_out;
wire [15:0] _U376_out;
wire [15:0] _U377_out;
wire [15:0] _U378_out;
wire [15:0] _U379_out;
wire [15:0] _U380_out;
wire [15:0] _U381_out;
wire [15:0] _U382_out;
wire [15:0] _U383_out;
wire [15:0] _U385_out;
wire [15:0] _U388_out;
wire [15:0] _U390_out;
wire [15:0] _U391_out;
wire [15:0] _U392_out;
wire [15:0] _U393_out;
wire [15:0] _U394_out;
wire [15:0] _U395_out;
wire [15:0] _U396_out;
wire [15:0] _U397_out;
wire [15:0] _U398_out;
wire [15:0] _U399_out;
wire [15:0] _U400_out;
wire [15:0] _U401_out;
wire [15:0] _U402_out;
wire [15:0] _U403_out;
wire [15:0] _U405_out;
wire [15:0] _U406_out;
wire [15:0] _U408_out;
wire [15:0] _U409_out;
wire [15:0] _U411_out;
wire [15:0] _U412_out;
wire [15:0] _U413_out;
wire [15:0] _U414_out;
wire [15:0] _U415_out;
wire [15:0] _U416_out;
wire [15:0] _U417_out;
wire [15:0] _U418_out;
wire [15:0] _U419_out;
wire [15:0] _U420_out;
wire [15:0] _U421_out;
wire [15:0] _U422_out;
wire [15:0] _U424_out;
wire [15:0] _U425_out;
wire [15:0] _U427_out;
wire [15:0] _U428_out;
wire [15:0] _U429_out;
wire [15:0] _U430_out;
wire [15:0] _U431_out;
wire [15:0] _U432_out;
wire [15:0] _U433_out;
wire [15:0] _U434_out;
wire [15:0] _U435_out;
wire [15:0] add_785_799_800_out;
wire [15:0] add_786_797_798_out;
wire [15:0] add_787_796_797_out;
wire [15:0] add_788_795_796_out;
wire [15:0] add_789_794_795_out;
wire [15:0] add_790_793_794_out;
wire [15:0] add_791_792_793_out;
wire [15:0] add_conv_stencil_2_798_799_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_10_hw_input_global_wrapper_stencil_10_786_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_11_hw_input_global_wrapper_stencil_11_787_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_12_hw_input_global_wrapper_stencil_12_788_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_13_hw_input_global_wrapper_stencil_13_789_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_14_hw_input_global_wrapper_stencil_14_790_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_15_hw_input_global_wrapper_stencil_15_791_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_16_hw_input_global_wrapper_stencil_16_792_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_9_hw_input_global_wrapper_stencil_9_785_out;
_U235_pt__U236 _U235 (
    .in(_U238_out),
    .out(_U235_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U237 (
    .in(in1_hw_input_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U237_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U238 (
    .in(_U237_out),
    .clk(clk),
    .out(_U238_out)
);
_U239_pt__U240 _U239 (
    .in(_U243_out),
    .out(_U239_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U241 (
    .in(in2_hw_kernel_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U241_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U242 (
    .in(_U241_out),
    .clk(clk),
    .out(_U242_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U243 (
    .in(_U242_out),
    .clk(clk),
    .out(_U243_out)
);
_U244_pt__U245 _U244 (
    .in(_U248_out),
    .out(_U244_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U246 (
    .in(in1_hw_input_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U246_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U247 (
    .in(_U246_out),
    .clk(clk),
    .out(_U247_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U248 (
    .in(_U247_out),
    .clk(clk),
    .out(_U248_out)
);
_U249_pt__U250 _U249 (
    .in(_U254_out),
    .out(_U249_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U251 (
    .in(in2_hw_kernel_global_wrapper_stencil[4]),
    .clk(clk),
    .out(_U251_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U252 (
    .in(_U251_out),
    .clk(clk),
    .out(_U252_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U253 (
    .in(_U252_out),
    .clk(clk),
    .out(_U253_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U254 (
    .in(_U253_out),
    .clk(clk),
    .out(_U254_out)
);
_U255_pt__U256 _U255 (
    .in(_U260_out),
    .out(_U255_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U257 (
    .in(in1_hw_input_global_wrapper_stencil[4]),
    .clk(clk),
    .out(_U257_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U258 (
    .in(_U257_out),
    .clk(clk),
    .out(_U258_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U259 (
    .in(_U258_out),
    .clk(clk),
    .out(_U259_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U260 (
    .in(_U259_out),
    .clk(clk),
    .out(_U260_out)
);
_U261_pt__U262 _U261 (
    .in(_U267_out),
    .out(_U261_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U263 (
    .in(in2_hw_kernel_global_wrapper_stencil[5]),
    .clk(clk),
    .out(_U263_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U264 (
    .in(_U263_out),
    .clk(clk),
    .out(_U264_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U265 (
    .in(_U264_out),
    .clk(clk),
    .out(_U265_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U266 (
    .in(_U265_out),
    .clk(clk),
    .out(_U266_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U267 (
    .in(_U266_out),
    .clk(clk),
    .out(_U267_out)
);
_U268_pt__U269 _U268 (
    .in(_U274_out),
    .out(_U268_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U270 (
    .in(in1_hw_input_global_wrapper_stencil[5]),
    .clk(clk),
    .out(_U270_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U271 (
    .in(_U270_out),
    .clk(clk),
    .out(_U271_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U272 (
    .in(_U271_out),
    .clk(clk),
    .out(_U272_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U273 (
    .in(_U272_out),
    .clk(clk),
    .out(_U273_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U274 (
    .in(_U273_out),
    .clk(clk),
    .out(_U274_out)
);
_U275_pt__U276 _U275 (
    .in(_U282_out),
    .out(_U275_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U277 (
    .in(in2_hw_kernel_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U277_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U278 (
    .in(_U277_out),
    .clk(clk),
    .out(_U278_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U279 (
    .in(_U278_out),
    .clk(clk),
    .out(_U279_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U280 (
    .in(_U279_out),
    .clk(clk),
    .out(_U280_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U281 (
    .in(_U280_out),
    .clk(clk),
    .out(_U281_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U282 (
    .in(_U281_out),
    .clk(clk),
    .out(_U282_out)
);
_U283_pt__U284 _U283 (
    .in(_U290_out),
    .out(_U283_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U285 (
    .in(in1_hw_input_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U285_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U286 (
    .in(_U285_out),
    .clk(clk),
    .out(_U286_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U287 (
    .in(_U286_out),
    .clk(clk),
    .out(_U287_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U288 (
    .in(_U287_out),
    .clk(clk),
    .out(_U288_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U289 (
    .in(_U288_out),
    .clk(clk),
    .out(_U289_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U290 (
    .in(_U289_out),
    .clk(clk),
    .out(_U290_out)
);
_U291_pt__U292 _U291 (
    .in(_U299_out),
    .out(_U291_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U293 (
    .in(in2_hw_kernel_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U293_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U294 (
    .in(_U293_out),
    .clk(clk),
    .out(_U294_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U295 (
    .in(_U294_out),
    .clk(clk),
    .out(_U295_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U296 (
    .in(_U295_out),
    .clk(clk),
    .out(_U296_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U297 (
    .in(_U296_out),
    .clk(clk),
    .out(_U297_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U298 (
    .in(_U297_out),
    .clk(clk),
    .out(_U298_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U299 (
    .in(_U298_out),
    .clk(clk),
    .out(_U299_out)
);
_U300_pt__U301 _U300 (
    .in(_U308_out),
    .out(_U300_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U302 (
    .in(in1_hw_input_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U302_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U303 (
    .in(_U302_out),
    .clk(clk),
    .out(_U303_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U304 (
    .in(_U303_out),
    .clk(clk),
    .out(_U304_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U305 (
    .in(_U304_out),
    .clk(clk),
    .out(_U305_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U306 (
    .in(_U305_out),
    .clk(clk),
    .out(_U306_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U307 (
    .in(_U306_out),
    .clk(clk),
    .out(_U307_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U308 (
    .in(_U307_out),
    .clk(clk),
    .out(_U308_out)
);
_U309_pt__U310 _U309 (
    .in(_U311_out),
    .out(_U309_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U311 (
    .in(add_789_794_795_out),
    .clk(clk),
    .out(_U311_out)
);
_U312_pt__U313 _U312 (
    .in(_U320_out),
    .out(_U312_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U314 (
    .in(mul_hw_kernel_global_wrapper_stencil_13_hw_input_global_wrapper_stencil_13_789_out),
    .clk(clk),
    .out(_U314_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U315 (
    .in(_U314_out),
    .clk(clk),
    .out(_U315_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U316 (
    .in(_U315_out),
    .clk(clk),
    .out(_U316_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U317 (
    .in(_U316_out),
    .clk(clk),
    .out(_U317_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U318 (
    .in(_U317_out),
    .clk(clk),
    .out(_U318_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U319 (
    .in(_U318_out),
    .clk(clk),
    .out(_U319_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U320 (
    .in(_U319_out),
    .clk(clk),
    .out(_U320_out)
);
_U321_pt__U322 _U321 (
    .in(_U323_out),
    .out(_U321_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U323 (
    .in(add_790_793_794_out),
    .clk(clk),
    .out(_U323_out)
);
_U324_pt__U325 _U324 (
    .in(_U330_out),
    .out(_U324_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U326 (
    .in(mul_hw_kernel_global_wrapper_stencil_14_hw_input_global_wrapper_stencil_14_790_out),
    .clk(clk),
    .out(_U326_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U327 (
    .in(_U326_out),
    .clk(clk),
    .out(_U327_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U328 (
    .in(_U327_out),
    .clk(clk),
    .out(_U328_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U329 (
    .in(_U328_out),
    .clk(clk),
    .out(_U329_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U330 (
    .in(_U329_out),
    .clk(clk),
    .out(_U330_out)
);
_U331_pt__U332 _U331 (
    .in(_U333_out),
    .out(_U331_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U333 (
    .in(add_791_792_793_out),
    .clk(clk),
    .out(_U333_out)
);
_U334_pt__U335 _U334 (
    .in(_U338_out),
    .out(_U334_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U336 (
    .in(mul_hw_kernel_global_wrapper_stencil_15_hw_input_global_wrapper_stencil_15_791_out),
    .clk(clk),
    .out(_U336_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U337 (
    .in(_U336_out),
    .clk(clk),
    .out(_U337_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U338 (
    .in(_U337_out),
    .clk(clk),
    .out(_U338_out)
);
_U339_pt__U340 _U339 (
    .in(_U342_out),
    .out(_U339_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U341 (
    .in(mul_hw_kernel_global_wrapper_stencil_16_hw_input_global_wrapper_stencil_16_792_out),
    .clk(clk),
    .out(_U341_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U342 (
    .in(_U341_out),
    .clk(clk),
    .out(_U342_out)
);
_U343_pt__U344 _U343 (
    .in(_U358_out),
    .out(_U343_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U345 (
    .in(in0_conv_stencil[0]),
    .clk(clk),
    .out(_U345_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U346 (
    .in(_U345_out),
    .clk(clk),
    .out(_U346_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U347 (
    .in(_U346_out),
    .clk(clk),
    .out(_U347_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U348 (
    .in(_U347_out),
    .clk(clk),
    .out(_U348_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U349 (
    .in(_U348_out),
    .clk(clk),
    .out(_U349_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U350 (
    .in(_U349_out),
    .clk(clk),
    .out(_U350_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U351 (
    .in(_U350_out),
    .clk(clk),
    .out(_U351_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U352 (
    .in(_U351_out),
    .clk(clk),
    .out(_U352_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U353 (
    .in(_U352_out),
    .clk(clk),
    .out(_U353_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U354 (
    .in(_U353_out),
    .clk(clk),
    .out(_U354_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U355 (
    .in(_U354_out),
    .clk(clk),
    .out(_U355_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U356 (
    .in(_U355_out),
    .clk(clk),
    .out(_U356_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U357 (
    .in(_U356_out),
    .clk(clk),
    .out(_U357_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U358 (
    .in(_U357_out),
    .clk(clk),
    .out(_U358_out)
);
_U359_pt__U360 _U359 (
    .in(in2_hw_kernel_global_wrapper_stencil[0]),
    .out(_U359_out)
);
_U361_pt__U362 _U361 (
    .in(in1_hw_input_global_wrapper_stencil[0]),
    .out(_U361_out)
);
_U363_pt__U364 _U363 (
    .in(_U365_out),
    .out(_U363_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U365 (
    .in(in2_hw_kernel_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U365_out)
);
_U366_pt__U367 _U366 (
    .in(_U368_out),
    .out(_U366_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U368 (
    .in(in1_hw_input_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U368_out)
);
_U369_pt__U370 _U369 (
    .in(_U372_out),
    .out(_U369_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U371 (
    .in(in2_hw_kernel_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U371_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U372 (
    .in(_U371_out),
    .clk(clk),
    .out(_U372_out)
);
_U373_pt__U374 _U373 (
    .in(_U382_out),
    .out(_U373_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U375 (
    .in(mul_hw_kernel_global_wrapper_stencil_9_hw_input_global_wrapper_stencil_9_785_out),
    .clk(clk),
    .out(_U375_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U376 (
    .in(_U375_out),
    .clk(clk),
    .out(_U376_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U377 (
    .in(_U376_out),
    .clk(clk),
    .out(_U377_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U378 (
    .in(_U377_out),
    .clk(clk),
    .out(_U378_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U379 (
    .in(_U378_out),
    .clk(clk),
    .out(_U379_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U380 (
    .in(_U379_out),
    .clk(clk),
    .out(_U380_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U381 (
    .in(_U380_out),
    .clk(clk),
    .out(_U381_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U382 (
    .in(_U381_out),
    .clk(clk),
    .out(_U382_out)
);
_U383_pt__U384 _U383 (
    .in(_U385_out),
    .out(_U383_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U385 (
    .in(add_conv_stencil_2_798_799_out),
    .clk(clk),
    .out(_U385_out)
);
_U386_pt__U387 _U386 (
    .in(add_785_799_800_out),
    .out(out_conv_stencil)
);
_U388_pt__U389 _U388 (
    .in(_U402_out),
    .out(_U388_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U390 (
    .in(mul_hw_kernel_global_wrapper_stencil_10_hw_input_global_wrapper_stencil_10_786_out),
    .clk(clk),
    .out(_U390_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U391 (
    .in(_U390_out),
    .clk(clk),
    .out(_U391_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U392 (
    .in(_U391_out),
    .clk(clk),
    .out(_U392_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U393 (
    .in(_U392_out),
    .clk(clk),
    .out(_U393_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U394 (
    .in(_U393_out),
    .clk(clk),
    .out(_U394_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U395 (
    .in(_U394_out),
    .clk(clk),
    .out(_U395_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U396 (
    .in(_U395_out),
    .clk(clk),
    .out(_U396_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U397 (
    .in(_U396_out),
    .clk(clk),
    .out(_U397_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U398 (
    .in(_U397_out),
    .clk(clk),
    .out(_U398_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U399 (
    .in(_U398_out),
    .clk(clk),
    .out(_U399_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U400 (
    .in(_U399_out),
    .clk(clk),
    .out(_U400_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U401 (
    .in(_U400_out),
    .clk(clk),
    .out(_U401_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U402 (
    .in(_U401_out),
    .clk(clk),
    .out(_U402_out)
);
_U403_pt__U404 _U403 (
    .in(_U405_out),
    .out(_U403_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U405 (
    .in(add_787_796_797_out),
    .clk(clk),
    .out(_U405_out)
);
_U406_pt__U407 _U406 (
    .in(_U408_out),
    .out(_U406_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U408 (
    .in(add_786_797_798_out),
    .clk(clk),
    .out(_U408_out)
);
_U409_pt__U410 _U409 (
    .in(_U421_out),
    .out(_U409_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U411 (
    .in(mul_hw_kernel_global_wrapper_stencil_11_hw_input_global_wrapper_stencil_11_787_out),
    .clk(clk),
    .out(_U411_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U412 (
    .in(_U411_out),
    .clk(clk),
    .out(_U412_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U413 (
    .in(_U412_out),
    .clk(clk),
    .out(_U413_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U414 (
    .in(_U413_out),
    .clk(clk),
    .out(_U414_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U415 (
    .in(_U414_out),
    .clk(clk),
    .out(_U415_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U416 (
    .in(_U415_out),
    .clk(clk),
    .out(_U416_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U417 (
    .in(_U416_out),
    .clk(clk),
    .out(_U417_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U418 (
    .in(_U417_out),
    .clk(clk),
    .out(_U418_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U419 (
    .in(_U418_out),
    .clk(clk),
    .out(_U419_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U420 (
    .in(_U419_out),
    .clk(clk),
    .out(_U420_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U421 (
    .in(_U420_out),
    .clk(clk),
    .out(_U421_out)
);
_U422_pt__U423 _U422 (
    .in(_U424_out),
    .out(_U422_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U424 (
    .in(add_788_795_796_out),
    .clk(clk),
    .out(_U424_out)
);
_U425_pt__U426 _U425 (
    .in(_U435_out),
    .out(_U425_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U427 (
    .in(mul_hw_kernel_global_wrapper_stencil_12_hw_input_global_wrapper_stencil_12_788_out),
    .clk(clk),
    .out(_U427_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U428 (
    .in(_U427_out),
    .clk(clk),
    .out(_U428_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U429 (
    .in(_U428_out),
    .clk(clk),
    .out(_U429_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U430 (
    .in(_U429_out),
    .clk(clk),
    .out(_U430_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U431 (
    .in(_U430_out),
    .clk(clk),
    .out(_U431_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U432 (
    .in(_U431_out),
    .clk(clk),
    .out(_U432_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U433 (
    .in(_U432_out),
    .clk(clk),
    .out(_U433_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U434 (
    .in(_U433_out),
    .clk(clk),
    .out(_U434_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U435 (
    .in(_U434_out),
    .clk(clk),
    .out(_U435_out)
);
assign add_785_799_800_out = 16'(_U373_out + _U383_out);
assign add_786_797_798_out = 16'(_U388_out + _U403_out);
assign add_787_796_797_out = 16'(_U409_out + _U422_out);
assign add_788_795_796_out = 16'(_U425_out + _U309_out);
assign add_789_794_795_out = 16'(_U312_out + _U321_out);
assign add_790_793_794_out = 16'(_U324_out + _U331_out);
assign add_791_792_793_out = 16'(_U334_out + _U339_out);
assign add_conv_stencil_2_798_799_out = 16'(_U343_out + _U406_out);
assign mul_hw_kernel_global_wrapper_stencil_10_hw_input_global_wrapper_stencil_10_786_out = 16'(_U359_out * _U361_out);
assign mul_hw_kernel_global_wrapper_stencil_11_hw_input_global_wrapper_stencil_11_787_out = 16'(_U363_out * _U366_out);
assign mul_hw_kernel_global_wrapper_stencil_12_hw_input_global_wrapper_stencil_12_788_out = 16'(_U369_out * _U235_out);
assign mul_hw_kernel_global_wrapper_stencil_13_hw_input_global_wrapper_stencil_13_789_out = 16'(_U239_out * _U244_out);
assign mul_hw_kernel_global_wrapper_stencil_14_hw_input_global_wrapper_stencil_14_790_out = 16'(_U249_out * _U255_out);
assign mul_hw_kernel_global_wrapper_stencil_15_hw_input_global_wrapper_stencil_15_791_out = 16'(_U261_out * _U268_out);
assign mul_hw_kernel_global_wrapper_stencil_16_hw_input_global_wrapper_stencil_16_792_out = 16'(_U275_out * _U283_out);
assign mul_hw_kernel_global_wrapper_stencil_9_hw_input_global_wrapper_stencil_9_785_out = 16'(_U291_out * _U300_out);
endmodule

module cu_op_hcompute_conv_stencil_9 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_9_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_9_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_9_read[0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[0];
hcompute_conv_stencil_9_pipelined inner_compute (
    .clk(clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_9_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U233_pt__U234 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U230_pt__U231 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U22_pt__U23 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_2_pipelined (
    output [15:0] out_conv_stencil
);
_U22_pt__U23 _U22 (
    .in(16'h0000),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_2 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_2_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U213_pt__U214 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U20_pt__U21 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_1_pipelined (
    output [15:0] out_conv_stencil
);
_U20_pt__U21 _U20 (
    .in(16'h0000),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_1 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_1_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U209_pt__U210 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U205_pt__U206 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U202_pt__U203 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U199_pt__U200 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U197_pt__U198 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U195_pt__U196 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U18_pt__U19 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_pipelined (
    output [15:0] out_conv_stencil
);
_U18_pt__U19 _U18 (
    .in(16'h0000),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U179_pt__U180 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U176_pt__U177 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U172_pt__U173 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U16_pt__U17 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_kernel_global_wrapper_stencil_pipelined (
    output [15:0] out_hw_kernel_global_wrapper_stencil,
    input [15:0] in0_hw_kernel_stencil [0:0]
);
_U16_pt__U17 _U16 (
    .in(in0_hw_kernel_stencil[0]),
    .out(out_hw_kernel_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_kernel_global_wrapper_stencil (
    input clk,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_kernel_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_kernel_stencil [0:0];
assign inner_compute_in0_hw_kernel_stencil[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
hcompute_hw_kernel_global_wrapper_stencil_pipelined inner_compute (
    .out_hw_kernel_global_wrapper_stencil(inner_compute_out_hw_kernel_global_wrapper_stencil),
    .in0_hw_kernel_stencil(inner_compute_in0_hw_kernel_stencil)
);
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = inner_compute_out_hw_kernel_global_wrapper_stencil;
endmodule

module _U169_pt__U170 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1656_pt__U1657 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_7_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
_U1656_pt__U1657 _U1656 (
    .in(in0_conv_stencil[0]),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil_7 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_7_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_7_read[0];
hcompute_hw_output_stencil_7_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1654_pt__U1655 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_6_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
_U1654_pt__U1655 _U1654 (
    .in(in0_conv_stencil[0]),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil_6 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_6_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_6_read[0];
hcompute_hw_output_stencil_6_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1652_pt__U1653 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_5_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
_U1652_pt__U1653 _U1652 (
    .in(in0_conv_stencil[0]),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil_5 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_5_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_5_read[0];
hcompute_hw_output_stencil_5_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1650_pt__U1651 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_4_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
_U1650_pt__U1651 _U1650 (
    .in(in0_conv_stencil[0]),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil_4 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_4_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_4_read[0];
hcompute_hw_output_stencil_4_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1648_pt__U1649 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_3_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
_U1648_pt__U1649 _U1648 (
    .in(in0_conv_stencil[0]),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil_3 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_3_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_3_read[0];
hcompute_hw_output_stencil_3_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1646_pt__U1647 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_2_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
_U1646_pt__U1647 _U1646 (
    .in(in0_conv_stencil[0]),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil_2 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_2_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_2_read[0];
hcompute_hw_output_stencil_2_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1644_pt__U1645 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_1_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
_U1644_pt__U1645 _U1644 (
    .in(in0_conv_stencil[0]),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil_1 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_1_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_1_read[0];
hcompute_hw_output_stencil_1_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1642_pt__U1643 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
_U1642_pt__U1643 _U1642 (
    .in(in0_conv_stencil[0]),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
hcompute_hw_output_stencil_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U163_pt__U164 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1628_pt__U1629 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1626_pt__U1627 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1623_pt__U1624 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U160_pt__U161 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1606_pt__U1607 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1604_pt__U1605 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1588_pt__U1589 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1585_pt__U1586 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1581_pt__U1582 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1578_pt__U1579 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1572_pt__U1573 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1563_pt__U1564 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1554_pt__U1555 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1546_pt__U1547 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1538_pt__U1539 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1535_pt__U1536 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U152_pt__U153 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1527_pt__U1528 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1524_pt__U1525 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1514_pt__U1515 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1511_pt__U1512 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U14_pt__U15 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_7_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
_U14_pt__U15 _U14 (
    .in(in0_hw_input_stencil[0]),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil_7 (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read[0];
hcompute_hw_input_global_wrapper_stencil_7_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U149_pt__U150 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1499_pt__U1500 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1496_pt__U1497 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1493_pt__U1494 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1486_pt__U1487 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1479_pt__U1480 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1473_pt__U1474 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1467_pt__U1468 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1462_pt__U1463 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1457_pt__U1458 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1453_pt__U1454 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1449_pt__U1450 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1446_pt__U1447 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1443_pt__U1444 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1441_pt__U1442 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_15_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U1441_out;
wire [15:0] _U1443_out;
wire [15:0] _U1445_out;
wire [15:0] _U1446_out;
wire [15:0] _U1448_out;
wire [15:0] _U1449_out;
wire [15:0] _U1451_out;
wire [15:0] _U1452_out;
wire [15:0] _U1453_out;
wire [15:0] _U1455_out;
wire [15:0] _U1456_out;
wire [15:0] _U1457_out;
wire [15:0] _U1459_out;
wire [15:0] _U1460_out;
wire [15:0] _U1461_out;
wire [15:0] _U1462_out;
wire [15:0] _U1464_out;
wire [15:0] _U1465_out;
wire [15:0] _U1466_out;
wire [15:0] _U1467_out;
wire [15:0] _U1469_out;
wire [15:0] _U1470_out;
wire [15:0] _U1471_out;
wire [15:0] _U1472_out;
wire [15:0] _U1473_out;
wire [15:0] _U1475_out;
wire [15:0] _U1476_out;
wire [15:0] _U1477_out;
wire [15:0] _U1478_out;
wire [15:0] _U1479_out;
wire [15:0] _U1481_out;
wire [15:0] _U1482_out;
wire [15:0] _U1483_out;
wire [15:0] _U1484_out;
wire [15:0] _U1485_out;
wire [15:0] _U1486_out;
wire [15:0] _U1488_out;
wire [15:0] _U1489_out;
wire [15:0] _U1490_out;
wire [15:0] _U1491_out;
wire [15:0] _U1492_out;
wire [15:0] _U1493_out;
wire [15:0] _U1495_out;
wire [15:0] _U1496_out;
wire [15:0] _U1498_out;
wire [15:0] _U1499_out;
wire [15:0] _U1501_out;
wire [15:0] _U1502_out;
wire [15:0] _U1503_out;
wire [15:0] _U1504_out;
wire [15:0] _U1505_out;
wire [15:0] _U1506_out;
wire [15:0] _U1507_out;
wire [15:0] _U1508_out;
wire [15:0] _U1509_out;
wire [15:0] _U1510_out;
wire [15:0] _U1511_out;
wire [15:0] _U1513_out;
wire [15:0] _U1514_out;
wire [15:0] _U1516_out;
wire [15:0] _U1517_out;
wire [15:0] _U1518_out;
wire [15:0] _U1519_out;
wire [15:0] _U1520_out;
wire [15:0] _U1521_out;
wire [15:0] _U1522_out;
wire [15:0] _U1523_out;
wire [15:0] _U1524_out;
wire [15:0] _U1526_out;
wire [15:0] _U1527_out;
wire [15:0] _U1529_out;
wire [15:0] _U1530_out;
wire [15:0] _U1531_out;
wire [15:0] _U1532_out;
wire [15:0] _U1533_out;
wire [15:0] _U1534_out;
wire [15:0] _U1535_out;
wire [15:0] _U1537_out;
wire [15:0] _U1538_out;
wire [15:0] _U1540_out;
wire [15:0] _U1541_out;
wire [15:0] _U1542_out;
wire [15:0] _U1543_out;
wire [15:0] _U1544_out;
wire [15:0] _U1545_out;
wire [15:0] _U1546_out;
wire [15:0] _U1548_out;
wire [15:0] _U1549_out;
wire [15:0] _U1550_out;
wire [15:0] _U1551_out;
wire [15:0] _U1552_out;
wire [15:0] _U1553_out;
wire [15:0] _U1554_out;
wire [15:0] _U1556_out;
wire [15:0] _U1557_out;
wire [15:0] _U1558_out;
wire [15:0] _U1559_out;
wire [15:0] _U1560_out;
wire [15:0] _U1561_out;
wire [15:0] _U1562_out;
wire [15:0] _U1563_out;
wire [15:0] _U1565_out;
wire [15:0] _U1566_out;
wire [15:0] _U1567_out;
wire [15:0] _U1568_out;
wire [15:0] _U1569_out;
wire [15:0] _U1570_out;
wire [15:0] _U1571_out;
wire [15:0] _U1572_out;
wire [15:0] _U1574_out;
wire [15:0] _U1575_out;
wire [15:0] _U1576_out;
wire [15:0] _U1577_out;
wire [15:0] _U1578_out;
wire [15:0] _U1580_out;
wire [15:0] _U1581_out;
wire [15:0] _U1583_out;
wire [15:0] _U1584_out;
wire [15:0] _U1585_out;
wire [15:0] _U1587_out;
wire [15:0] _U1588_out;
wire [15:0] _U1590_out;
wire [15:0] _U1591_out;
wire [15:0] _U1592_out;
wire [15:0] _U1593_out;
wire [15:0] _U1594_out;
wire [15:0] _U1595_out;
wire [15:0] _U1596_out;
wire [15:0] _U1597_out;
wire [15:0] _U1598_out;
wire [15:0] _U1599_out;
wire [15:0] _U1600_out;
wire [15:0] _U1601_out;
wire [15:0] _U1602_out;
wire [15:0] _U1603_out;
wire [15:0] _U1604_out;
wire [15:0] _U1606_out;
wire [15:0] _U1608_out;
wire [15:0] _U1609_out;
wire [15:0] _U1610_out;
wire [15:0] _U1611_out;
wire [15:0] _U1612_out;
wire [15:0] _U1613_out;
wire [15:0] _U1614_out;
wire [15:0] _U1615_out;
wire [15:0] _U1616_out;
wire [15:0] _U1617_out;
wire [15:0] _U1618_out;
wire [15:0] _U1619_out;
wire [15:0] _U1620_out;
wire [15:0] _U1621_out;
wire [15:0] _U1622_out;
wire [15:0] _U1623_out;
wire [15:0] _U1625_out;
wire [15:0] _U1628_out;
wire [15:0] _U1630_out;
wire [15:0] _U1631_out;
wire [15:0] _U1632_out;
wire [15:0] _U1633_out;
wire [15:0] _U1634_out;
wire [15:0] _U1635_out;
wire [15:0] _U1636_out;
wire [15:0] _U1637_out;
wire [15:0] _U1638_out;
wire [15:0] _U1639_out;
wire [15:0] _U1640_out;
wire [15:0] _U1641_out;
wire [15:0] add_1187_1201_1202_out;
wire [15:0] add_1188_1199_1200_out;
wire [15:0] add_1189_1198_1199_out;
wire [15:0] add_1190_1197_1198_out;
wire [15:0] add_1191_1196_1197_out;
wire [15:0] add_1192_1195_1196_out;
wire [15:0] add_1193_1194_1195_out;
wire [15:0] add_conv_stencil_8_1200_1201_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_57_hw_input_global_wrapper_stencil_57_1187_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_58_hw_input_global_wrapper_stencil_58_1188_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_59_hw_input_global_wrapper_stencil_59_1189_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_60_hw_input_global_wrapper_stencil_60_1190_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_61_hw_input_global_wrapper_stencil_61_1191_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_62_hw_input_global_wrapper_stencil_62_1192_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_63_hw_input_global_wrapper_stencil_63_1193_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_64_hw_input_global_wrapper_stencil_64_1194_out;
_U1441_pt__U1442 _U1441 (
    .in(in1_hw_input_global_wrapper_stencil[0]),
    .out(_U1441_out)
);
_U1443_pt__U1444 _U1443 (
    .in(_U1445_out),
    .out(_U1443_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1445 (
    .in(in2_hw_kernel_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U1445_out)
);
_U1446_pt__U1447 _U1446 (
    .in(_U1448_out),
    .out(_U1446_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1448 (
    .in(in1_hw_input_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U1448_out)
);
_U1449_pt__U1450 _U1449 (
    .in(_U1452_out),
    .out(_U1449_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1451 (
    .in(in2_hw_kernel_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U1451_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1452 (
    .in(_U1451_out),
    .clk(clk),
    .out(_U1452_out)
);
_U1453_pt__U1454 _U1453 (
    .in(_U1456_out),
    .out(_U1453_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1455 (
    .in(in1_hw_input_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U1455_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1456 (
    .in(_U1455_out),
    .clk(clk),
    .out(_U1456_out)
);
_U1457_pt__U1458 _U1457 (
    .in(_U1461_out),
    .out(_U1457_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1459 (
    .in(in2_hw_kernel_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U1459_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1460 (
    .in(_U1459_out),
    .clk(clk),
    .out(_U1460_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1461 (
    .in(_U1460_out),
    .clk(clk),
    .out(_U1461_out)
);
_U1462_pt__U1463 _U1462 (
    .in(_U1466_out),
    .out(_U1462_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1464 (
    .in(in1_hw_input_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U1464_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1465 (
    .in(_U1464_out),
    .clk(clk),
    .out(_U1465_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1466 (
    .in(_U1465_out),
    .clk(clk),
    .out(_U1466_out)
);
_U1467_pt__U1468 _U1467 (
    .in(_U1472_out),
    .out(_U1467_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1469 (
    .in(in2_hw_kernel_global_wrapper_stencil[4]),
    .clk(clk),
    .out(_U1469_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1470 (
    .in(_U1469_out),
    .clk(clk),
    .out(_U1470_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1471 (
    .in(_U1470_out),
    .clk(clk),
    .out(_U1471_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1472 (
    .in(_U1471_out),
    .clk(clk),
    .out(_U1472_out)
);
_U1473_pt__U1474 _U1473 (
    .in(_U1478_out),
    .out(_U1473_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1475 (
    .in(in1_hw_input_global_wrapper_stencil[4]),
    .clk(clk),
    .out(_U1475_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1476 (
    .in(_U1475_out),
    .clk(clk),
    .out(_U1476_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1477 (
    .in(_U1476_out),
    .clk(clk),
    .out(_U1477_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1478 (
    .in(_U1477_out),
    .clk(clk),
    .out(_U1478_out)
);
_U1479_pt__U1480 _U1479 (
    .in(_U1485_out),
    .out(_U1479_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1481 (
    .in(in2_hw_kernel_global_wrapper_stencil[5]),
    .clk(clk),
    .out(_U1481_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1482 (
    .in(_U1481_out),
    .clk(clk),
    .out(_U1482_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1483 (
    .in(_U1482_out),
    .clk(clk),
    .out(_U1483_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1484 (
    .in(_U1483_out),
    .clk(clk),
    .out(_U1484_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1485 (
    .in(_U1484_out),
    .clk(clk),
    .out(_U1485_out)
);
_U1486_pt__U1487 _U1486 (
    .in(_U1492_out),
    .out(_U1486_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1488 (
    .in(in1_hw_input_global_wrapper_stencil[5]),
    .clk(clk),
    .out(_U1488_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1489 (
    .in(_U1488_out),
    .clk(clk),
    .out(_U1489_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1490 (
    .in(_U1489_out),
    .clk(clk),
    .out(_U1490_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1491 (
    .in(_U1490_out),
    .clk(clk),
    .out(_U1491_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1492 (
    .in(_U1491_out),
    .clk(clk),
    .out(_U1492_out)
);
_U1493_pt__U1494 _U1493 (
    .in(_U1495_out),
    .out(_U1493_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1495 (
    .in(add_1189_1198_1199_out),
    .clk(clk),
    .out(_U1495_out)
);
_U1496_pt__U1497 _U1496 (
    .in(_U1498_out),
    .out(_U1496_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1498 (
    .in(add_1188_1199_1200_out),
    .clk(clk),
    .out(_U1498_out)
);
_U1499_pt__U1500 _U1499 (
    .in(_U1510_out),
    .out(_U1499_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1501 (
    .in(mul_hw_kernel_global_wrapper_stencil_59_hw_input_global_wrapper_stencil_59_1189_out),
    .clk(clk),
    .out(_U1501_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1502 (
    .in(_U1501_out),
    .clk(clk),
    .out(_U1502_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1503 (
    .in(_U1502_out),
    .clk(clk),
    .out(_U1503_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1504 (
    .in(_U1503_out),
    .clk(clk),
    .out(_U1504_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1505 (
    .in(_U1504_out),
    .clk(clk),
    .out(_U1505_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1506 (
    .in(_U1505_out),
    .clk(clk),
    .out(_U1506_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1507 (
    .in(_U1506_out),
    .clk(clk),
    .out(_U1507_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1508 (
    .in(_U1507_out),
    .clk(clk),
    .out(_U1508_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1509 (
    .in(_U1508_out),
    .clk(clk),
    .out(_U1509_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1510 (
    .in(_U1509_out),
    .clk(clk),
    .out(_U1510_out)
);
_U1511_pt__U1512 _U1511 (
    .in(_U1513_out),
    .out(_U1511_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1513 (
    .in(add_1190_1197_1198_out),
    .clk(clk),
    .out(_U1513_out)
);
_U1514_pt__U1515 _U1514 (
    .in(_U1523_out),
    .out(_U1514_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1516 (
    .in(mul_hw_kernel_global_wrapper_stencil_60_hw_input_global_wrapper_stencil_60_1190_out),
    .clk(clk),
    .out(_U1516_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1517 (
    .in(_U1516_out),
    .clk(clk),
    .out(_U1517_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1518 (
    .in(_U1517_out),
    .clk(clk),
    .out(_U1518_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1519 (
    .in(_U1518_out),
    .clk(clk),
    .out(_U1519_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1520 (
    .in(_U1519_out),
    .clk(clk),
    .out(_U1520_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1521 (
    .in(_U1520_out),
    .clk(clk),
    .out(_U1521_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1522 (
    .in(_U1521_out),
    .clk(clk),
    .out(_U1522_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1523 (
    .in(_U1522_out),
    .clk(clk),
    .out(_U1523_out)
);
_U1524_pt__U1525 _U1524 (
    .in(_U1526_out),
    .out(_U1524_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1526 (
    .in(add_1191_1196_1197_out),
    .clk(clk),
    .out(_U1526_out)
);
_U1527_pt__U1528 _U1527 (
    .in(_U1534_out),
    .out(_U1527_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1529 (
    .in(mul_hw_kernel_global_wrapper_stencil_61_hw_input_global_wrapper_stencil_61_1191_out),
    .clk(clk),
    .out(_U1529_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1530 (
    .in(_U1529_out),
    .clk(clk),
    .out(_U1530_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1531 (
    .in(_U1530_out),
    .clk(clk),
    .out(_U1531_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1532 (
    .in(_U1531_out),
    .clk(clk),
    .out(_U1532_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1533 (
    .in(_U1532_out),
    .clk(clk),
    .out(_U1533_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1534 (
    .in(_U1533_out),
    .clk(clk),
    .out(_U1534_out)
);
_U1535_pt__U1536 _U1535 (
    .in(_U1537_out),
    .out(_U1535_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1537 (
    .in(add_1192_1195_1196_out),
    .clk(clk),
    .out(_U1537_out)
);
_U1538_pt__U1539 _U1538 (
    .in(_U1545_out),
    .out(_U1538_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1540 (
    .in(in2_hw_kernel_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U1540_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1541 (
    .in(_U1540_out),
    .clk(clk),
    .out(_U1541_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1542 (
    .in(_U1541_out),
    .clk(clk),
    .out(_U1542_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1543 (
    .in(_U1542_out),
    .clk(clk),
    .out(_U1543_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1544 (
    .in(_U1543_out),
    .clk(clk),
    .out(_U1544_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1545 (
    .in(_U1544_out),
    .clk(clk),
    .out(_U1545_out)
);
_U1546_pt__U1547 _U1546 (
    .in(_U1553_out),
    .out(_U1546_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1548 (
    .in(in1_hw_input_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U1548_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1549 (
    .in(_U1548_out),
    .clk(clk),
    .out(_U1549_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1550 (
    .in(_U1549_out),
    .clk(clk),
    .out(_U1550_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1551 (
    .in(_U1550_out),
    .clk(clk),
    .out(_U1551_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1552 (
    .in(_U1551_out),
    .clk(clk),
    .out(_U1552_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1553 (
    .in(_U1552_out),
    .clk(clk),
    .out(_U1553_out)
);
_U1554_pt__U1555 _U1554 (
    .in(_U1562_out),
    .out(_U1554_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1556 (
    .in(in2_hw_kernel_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U1556_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1557 (
    .in(_U1556_out),
    .clk(clk),
    .out(_U1557_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1558 (
    .in(_U1557_out),
    .clk(clk),
    .out(_U1558_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1559 (
    .in(_U1558_out),
    .clk(clk),
    .out(_U1559_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1560 (
    .in(_U1559_out),
    .clk(clk),
    .out(_U1560_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1561 (
    .in(_U1560_out),
    .clk(clk),
    .out(_U1561_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1562 (
    .in(_U1561_out),
    .clk(clk),
    .out(_U1562_out)
);
_U1563_pt__U1564 _U1563 (
    .in(_U1571_out),
    .out(_U1563_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1565 (
    .in(in1_hw_input_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U1565_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1566 (
    .in(_U1565_out),
    .clk(clk),
    .out(_U1566_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1567 (
    .in(_U1566_out),
    .clk(clk),
    .out(_U1567_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1568 (
    .in(_U1567_out),
    .clk(clk),
    .out(_U1568_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1569 (
    .in(_U1568_out),
    .clk(clk),
    .out(_U1569_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1570 (
    .in(_U1569_out),
    .clk(clk),
    .out(_U1570_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1571 (
    .in(_U1570_out),
    .clk(clk),
    .out(_U1571_out)
);
_U1572_pt__U1573 _U1572 (
    .in(_U1577_out),
    .out(_U1572_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1574 (
    .in(mul_hw_kernel_global_wrapper_stencil_62_hw_input_global_wrapper_stencil_62_1192_out),
    .clk(clk),
    .out(_U1574_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1575 (
    .in(_U1574_out),
    .clk(clk),
    .out(_U1575_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1576 (
    .in(_U1575_out),
    .clk(clk),
    .out(_U1576_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1577 (
    .in(_U1576_out),
    .clk(clk),
    .out(_U1577_out)
);
_U1578_pt__U1579 _U1578 (
    .in(_U1580_out),
    .out(_U1578_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1580 (
    .in(add_1193_1194_1195_out),
    .clk(clk),
    .out(_U1580_out)
);
_U1581_pt__U1582 _U1581 (
    .in(_U1584_out),
    .out(_U1581_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1583 (
    .in(mul_hw_kernel_global_wrapper_stencil_63_hw_input_global_wrapper_stencil_63_1193_out),
    .clk(clk),
    .out(_U1583_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1584 (
    .in(_U1583_out),
    .clk(clk),
    .out(_U1584_out)
);
_U1585_pt__U1586 _U1585 (
    .in(_U1587_out),
    .out(_U1585_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1587 (
    .in(mul_hw_kernel_global_wrapper_stencil_64_hw_input_global_wrapper_stencil_64_1194_out),
    .clk(clk),
    .out(_U1587_out)
);
_U1588_pt__U1589 _U1588 (
    .in(_U1603_out),
    .out(_U1588_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1590 (
    .in(in0_conv_stencil[0]),
    .clk(clk),
    .out(_U1590_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1591 (
    .in(_U1590_out),
    .clk(clk),
    .out(_U1591_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1592 (
    .in(_U1591_out),
    .clk(clk),
    .out(_U1592_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1593 (
    .in(_U1592_out),
    .clk(clk),
    .out(_U1593_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1594 (
    .in(_U1593_out),
    .clk(clk),
    .out(_U1594_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1595 (
    .in(_U1594_out),
    .clk(clk),
    .out(_U1595_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1596 (
    .in(_U1595_out),
    .clk(clk),
    .out(_U1596_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1597 (
    .in(_U1596_out),
    .clk(clk),
    .out(_U1597_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1598 (
    .in(_U1597_out),
    .clk(clk),
    .out(_U1598_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1599 (
    .in(_U1598_out),
    .clk(clk),
    .out(_U1599_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1600 (
    .in(_U1599_out),
    .clk(clk),
    .out(_U1600_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1601 (
    .in(_U1600_out),
    .clk(clk),
    .out(_U1601_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1602 (
    .in(_U1601_out),
    .clk(clk),
    .out(_U1602_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1603 (
    .in(_U1602_out),
    .clk(clk),
    .out(_U1603_out)
);
_U1604_pt__U1605 _U1604 (
    .in(in2_hw_kernel_global_wrapper_stencil[0]),
    .out(_U1604_out)
);
_U1606_pt__U1607 _U1606 (
    .in(_U1622_out),
    .out(_U1606_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1608 (
    .in(mul_hw_kernel_global_wrapper_stencil_57_hw_input_global_wrapper_stencil_57_1187_out),
    .clk(clk),
    .out(_U1608_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1609 (
    .in(_U1608_out),
    .clk(clk),
    .out(_U1609_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1610 (
    .in(_U1609_out),
    .clk(clk),
    .out(_U1610_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1611 (
    .in(_U1610_out),
    .clk(clk),
    .out(_U1611_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1612 (
    .in(_U1611_out),
    .clk(clk),
    .out(_U1612_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1613 (
    .in(_U1612_out),
    .clk(clk),
    .out(_U1613_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1614 (
    .in(_U1613_out),
    .clk(clk),
    .out(_U1614_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1615 (
    .in(_U1614_out),
    .clk(clk),
    .out(_U1615_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1616 (
    .in(_U1615_out),
    .clk(clk),
    .out(_U1616_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1617 (
    .in(_U1616_out),
    .clk(clk),
    .out(_U1617_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1618 (
    .in(_U1617_out),
    .clk(clk),
    .out(_U1618_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1619 (
    .in(_U1618_out),
    .clk(clk),
    .out(_U1619_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1620 (
    .in(_U1619_out),
    .clk(clk),
    .out(_U1620_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1621 (
    .in(_U1620_out),
    .clk(clk),
    .out(_U1621_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1622 (
    .in(_U1621_out),
    .clk(clk),
    .out(_U1622_out)
);
_U1623_pt__U1624 _U1623 (
    .in(_U1625_out),
    .out(_U1623_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1625 (
    .in(add_conv_stencil_8_1200_1201_out),
    .clk(clk),
    .out(_U1625_out)
);
_U1626_pt__U1627 _U1626 (
    .in(add_1187_1201_1202_out),
    .out(out_conv_stencil)
);
_U1628_pt__U1629 _U1628 (
    .in(_U1641_out),
    .out(_U1628_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1630 (
    .in(mul_hw_kernel_global_wrapper_stencil_58_hw_input_global_wrapper_stencil_58_1188_out),
    .clk(clk),
    .out(_U1630_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1631 (
    .in(_U1630_out),
    .clk(clk),
    .out(_U1631_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1632 (
    .in(_U1631_out),
    .clk(clk),
    .out(_U1632_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1633 (
    .in(_U1632_out),
    .clk(clk),
    .out(_U1633_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1634 (
    .in(_U1633_out),
    .clk(clk),
    .out(_U1634_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1635 (
    .in(_U1634_out),
    .clk(clk),
    .out(_U1635_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1636 (
    .in(_U1635_out),
    .clk(clk),
    .out(_U1636_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1637 (
    .in(_U1636_out),
    .clk(clk),
    .out(_U1637_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1638 (
    .in(_U1637_out),
    .clk(clk),
    .out(_U1638_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1639 (
    .in(_U1638_out),
    .clk(clk),
    .out(_U1639_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1640 (
    .in(_U1639_out),
    .clk(clk),
    .out(_U1640_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1641 (
    .in(_U1640_out),
    .clk(clk),
    .out(_U1641_out)
);
assign add_1187_1201_1202_out = 16'(_U1606_out + _U1623_out);
assign add_1188_1199_1200_out = 16'(_U1628_out + _U1493_out);
assign add_1189_1198_1199_out = 16'(_U1499_out + _U1511_out);
assign add_1190_1197_1198_out = 16'(_U1514_out + _U1524_out);
assign add_1191_1196_1197_out = 16'(_U1527_out + _U1535_out);
assign add_1192_1195_1196_out = 16'(_U1572_out + _U1578_out);
assign add_1193_1194_1195_out = 16'(_U1581_out + _U1585_out);
assign add_conv_stencil_8_1200_1201_out = 16'(_U1588_out + _U1496_out);
assign mul_hw_kernel_global_wrapper_stencil_57_hw_input_global_wrapper_stencil_57_1187_out = 16'(_U1604_out * _U1441_out);
assign mul_hw_kernel_global_wrapper_stencil_58_hw_input_global_wrapper_stencil_58_1188_out = 16'(_U1443_out * _U1446_out);
assign mul_hw_kernel_global_wrapper_stencil_59_hw_input_global_wrapper_stencil_59_1189_out = 16'(_U1449_out * _U1453_out);
assign mul_hw_kernel_global_wrapper_stencil_60_hw_input_global_wrapper_stencil_60_1190_out = 16'(_U1457_out * _U1462_out);
assign mul_hw_kernel_global_wrapper_stencil_61_hw_input_global_wrapper_stencil_61_1191_out = 16'(_U1467_out * _U1473_out);
assign mul_hw_kernel_global_wrapper_stencil_62_hw_input_global_wrapper_stencil_62_1192_out = 16'(_U1479_out * _U1486_out);
assign mul_hw_kernel_global_wrapper_stencil_63_hw_input_global_wrapper_stencil_63_1193_out = 16'(_U1538_out * _U1546_out);
assign mul_hw_kernel_global_wrapper_stencil_64_hw_input_global_wrapper_stencil_64_1194_out = 16'(_U1554_out * _U1563_out);
endmodule

module cu_op_hcompute_conv_stencil_15 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_15_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_15_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_15_read[0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[0];
hcompute_conv_stencil_15_pipelined inner_compute (
    .clk(clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_15_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U1432_pt__U1433 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1429_pt__U1430 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1426_pt__U1427 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1421_pt__U1422 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1418_pt__U1419 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1415_pt__U1416 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1412_pt__U1413 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1403_pt__U1404 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U139_pt__U140 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1394_pt__U1395 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1386_pt__U1387 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1378_pt__U1379 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1371_pt__U1372 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U136_pt__U137 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1365_pt__U1366 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1359_pt__U1360 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1354_pt__U1355 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1349_pt__U1350 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1336_pt__U1337 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1334_pt__U1335 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1331_pt__U1332 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1314_pt__U1315 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1307_pt__U1308 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1304_pt__U1305 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U12_pt__U13 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_6_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
_U12_pt__U13 _U12 (
    .in(in0_hw_input_stencil[0]),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil_6 (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read[0];
hcompute_hw_input_global_wrapper_stencil_6_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U1295_pt__U1296 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1292_pt__U1293 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1281_pt__U1282 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1278_pt__U1279 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1275_pt__U1276 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1271_pt__U1272 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1267_pt__U1268 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1265_pt__U1266 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1263_pt__U1264 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U124_pt__U125 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1247_pt__U1248 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1240_pt__U1241 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_14_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U1240_out;
wire [15:0] _U1242_out;
wire [15:0] _U1243_out;
wire [15:0] _U1244_out;
wire [15:0] _U1245_out;
wire [15:0] _U1246_out;
wire [15:0] _U1247_out;
wire [15:0] _U1249_out;
wire [15:0] _U1250_out;
wire [15:0] _U1251_out;
wire [15:0] _U1252_out;
wire [15:0] _U1253_out;
wire [15:0] _U1254_out;
wire [15:0] _U1255_out;
wire [15:0] _U1256_out;
wire [15:0] _U1257_out;
wire [15:0] _U1258_out;
wire [15:0] _U1259_out;
wire [15:0] _U1260_out;
wire [15:0] _U1261_out;
wire [15:0] _U1262_out;
wire [15:0] _U1263_out;
wire [15:0] _U1265_out;
wire [15:0] _U1267_out;
wire [15:0] _U1269_out;
wire [15:0] _U1270_out;
wire [15:0] _U1271_out;
wire [15:0] _U1273_out;
wire [15:0] _U1274_out;
wire [15:0] _U1275_out;
wire [15:0] _U1277_out;
wire [15:0] _U1278_out;
wire [15:0] _U1280_out;
wire [15:0] _U1281_out;
wire [15:0] _U1283_out;
wire [15:0] _U1284_out;
wire [15:0] _U1285_out;
wire [15:0] _U1286_out;
wire [15:0] _U1287_out;
wire [15:0] _U1288_out;
wire [15:0] _U1289_out;
wire [15:0] _U1290_out;
wire [15:0] _U1291_out;
wire [15:0] _U1292_out;
wire [15:0] _U1294_out;
wire [15:0] _U1295_out;
wire [15:0] _U1297_out;
wire [15:0] _U1298_out;
wire [15:0] _U1299_out;
wire [15:0] _U1300_out;
wire [15:0] _U1301_out;
wire [15:0] _U1302_out;
wire [15:0] _U1303_out;
wire [15:0] _U1304_out;
wire [15:0] _U1306_out;
wire [15:0] _U1307_out;
wire [15:0] _U1309_out;
wire [15:0] _U1310_out;
wire [15:0] _U1311_out;
wire [15:0] _U1312_out;
wire [15:0] _U1313_out;
wire [15:0] _U1314_out;
wire [15:0] _U1316_out;
wire [15:0] _U1317_out;
wire [15:0] _U1318_out;
wire [15:0] _U1319_out;
wire [15:0] _U1320_out;
wire [15:0] _U1321_out;
wire [15:0] _U1322_out;
wire [15:0] _U1323_out;
wire [15:0] _U1324_out;
wire [15:0] _U1325_out;
wire [15:0] _U1326_out;
wire [15:0] _U1327_out;
wire [15:0] _U1328_out;
wire [15:0] _U1329_out;
wire [15:0] _U1330_out;
wire [15:0] _U1331_out;
wire [15:0] _U1333_out;
wire [15:0] _U1336_out;
wire [15:0] _U1338_out;
wire [15:0] _U1339_out;
wire [15:0] _U1340_out;
wire [15:0] _U1341_out;
wire [15:0] _U1342_out;
wire [15:0] _U1343_out;
wire [15:0] _U1344_out;
wire [15:0] _U1345_out;
wire [15:0] _U1346_out;
wire [15:0] _U1347_out;
wire [15:0] _U1348_out;
wire [15:0] _U1349_out;
wire [15:0] _U1351_out;
wire [15:0] _U1352_out;
wire [15:0] _U1353_out;
wire [15:0] _U1354_out;
wire [15:0] _U1356_out;
wire [15:0] _U1357_out;
wire [15:0] _U1358_out;
wire [15:0] _U1359_out;
wire [15:0] _U1361_out;
wire [15:0] _U1362_out;
wire [15:0] _U1363_out;
wire [15:0] _U1364_out;
wire [15:0] _U1365_out;
wire [15:0] _U1367_out;
wire [15:0] _U1368_out;
wire [15:0] _U1369_out;
wire [15:0] _U1370_out;
wire [15:0] _U1371_out;
wire [15:0] _U1373_out;
wire [15:0] _U1374_out;
wire [15:0] _U1375_out;
wire [15:0] _U1376_out;
wire [15:0] _U1377_out;
wire [15:0] _U1378_out;
wire [15:0] _U1380_out;
wire [15:0] _U1381_out;
wire [15:0] _U1382_out;
wire [15:0] _U1383_out;
wire [15:0] _U1384_out;
wire [15:0] _U1385_out;
wire [15:0] _U1386_out;
wire [15:0] _U1388_out;
wire [15:0] _U1389_out;
wire [15:0] _U1390_out;
wire [15:0] _U1391_out;
wire [15:0] _U1392_out;
wire [15:0] _U1393_out;
wire [15:0] _U1394_out;
wire [15:0] _U1396_out;
wire [15:0] _U1397_out;
wire [15:0] _U1398_out;
wire [15:0] _U1399_out;
wire [15:0] _U1400_out;
wire [15:0] _U1401_out;
wire [15:0] _U1402_out;
wire [15:0] _U1403_out;
wire [15:0] _U1405_out;
wire [15:0] _U1406_out;
wire [15:0] _U1407_out;
wire [15:0] _U1408_out;
wire [15:0] _U1409_out;
wire [15:0] _U1410_out;
wire [15:0] _U1411_out;
wire [15:0] _U1412_out;
wire [15:0] _U1414_out;
wire [15:0] _U1415_out;
wire [15:0] _U1417_out;
wire [15:0] _U1418_out;
wire [15:0] _U1420_out;
wire [15:0] _U1421_out;
wire [15:0] _U1423_out;
wire [15:0] _U1424_out;
wire [15:0] _U1425_out;
wire [15:0] _U1426_out;
wire [15:0] _U1428_out;
wire [15:0] _U1429_out;
wire [15:0] _U1431_out;
wire [15:0] _U1432_out;
wire [15:0] _U1434_out;
wire [15:0] _U1435_out;
wire [15:0] _U1436_out;
wire [15:0] _U1437_out;
wire [15:0] _U1438_out;
wire [15:0] _U1439_out;
wire [15:0] _U1440_out;
wire [15:0] add_1120_1134_1135_out;
wire [15:0] add_1121_1132_1133_out;
wire [15:0] add_1122_1131_1132_out;
wire [15:0] add_1123_1130_1131_out;
wire [15:0] add_1124_1129_1130_out;
wire [15:0] add_1125_1128_1129_out;
wire [15:0] add_1126_1127_1128_out;
wire [15:0] add_conv_stencil_7_1133_1134_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_49_hw_input_global_wrapper_stencil_49_1120_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_50_hw_input_global_wrapper_stencil_50_1121_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_51_hw_input_global_wrapper_stencil_51_1122_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_52_hw_input_global_wrapper_stencil_52_1123_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_53_hw_input_global_wrapper_stencil_53_1124_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_54_hw_input_global_wrapper_stencil_54_1125_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_55_hw_input_global_wrapper_stencil_55_1126_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_56_hw_input_global_wrapper_stencil_56_1127_out;
_U1240_pt__U1241 _U1240 (
    .in(_U1246_out),
    .out(_U1240_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1242 (
    .in(in1_hw_input_global_wrapper_stencil[4]),
    .clk(clk),
    .out(_U1242_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1243 (
    .in(_U1242_out),
    .clk(clk),
    .out(_U1243_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1244 (
    .in(_U1243_out),
    .clk(clk),
    .out(_U1244_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1245 (
    .in(_U1244_out),
    .clk(clk),
    .out(_U1245_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1246 (
    .in(_U1245_out),
    .clk(clk),
    .out(_U1246_out)
);
_U1247_pt__U1248 _U1247 (
    .in(_U1262_out),
    .out(_U1247_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1249 (
    .in(in0_conv_stencil[0]),
    .clk(clk),
    .out(_U1249_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1250 (
    .in(_U1249_out),
    .clk(clk),
    .out(_U1250_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1251 (
    .in(_U1250_out),
    .clk(clk),
    .out(_U1251_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1252 (
    .in(_U1251_out),
    .clk(clk),
    .out(_U1252_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1253 (
    .in(_U1252_out),
    .clk(clk),
    .out(_U1253_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1254 (
    .in(_U1253_out),
    .clk(clk),
    .out(_U1254_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1255 (
    .in(_U1254_out),
    .clk(clk),
    .out(_U1255_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1256 (
    .in(_U1255_out),
    .clk(clk),
    .out(_U1256_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1257 (
    .in(_U1256_out),
    .clk(clk),
    .out(_U1257_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1258 (
    .in(_U1257_out),
    .clk(clk),
    .out(_U1258_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1259 (
    .in(_U1258_out),
    .clk(clk),
    .out(_U1259_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1260 (
    .in(_U1259_out),
    .clk(clk),
    .out(_U1260_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1261 (
    .in(_U1260_out),
    .clk(clk),
    .out(_U1261_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1262 (
    .in(_U1261_out),
    .clk(clk),
    .out(_U1262_out)
);
_U1263_pt__U1264 _U1263 (
    .in(in2_hw_kernel_global_wrapper_stencil[0]),
    .out(_U1263_out)
);
_U1265_pt__U1266 _U1265 (
    .in(in1_hw_input_global_wrapper_stencil[0]),
    .out(_U1265_out)
);
_U1267_pt__U1268 _U1267 (
    .in(_U1270_out),
    .out(_U1267_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1269 (
    .in(in2_hw_kernel_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U1269_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1270 (
    .in(_U1269_out),
    .clk(clk),
    .out(_U1270_out)
);
_U1271_pt__U1272 _U1271 (
    .in(_U1274_out),
    .out(_U1271_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1273 (
    .in(in1_hw_input_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U1273_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1274 (
    .in(_U1273_out),
    .clk(clk),
    .out(_U1274_out)
);
_U1275_pt__U1276 _U1275 (
    .in(_U1277_out),
    .out(_U1275_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1277 (
    .in(add_1122_1131_1132_out),
    .clk(clk),
    .out(_U1277_out)
);
_U1278_pt__U1279 _U1278 (
    .in(_U1280_out),
    .out(_U1278_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1280 (
    .in(add_1121_1132_1133_out),
    .clk(clk),
    .out(_U1280_out)
);
_U1281_pt__U1282 _U1281 (
    .in(_U1291_out),
    .out(_U1281_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1283 (
    .in(mul_hw_kernel_global_wrapper_stencil_51_hw_input_global_wrapper_stencil_51_1122_out),
    .clk(clk),
    .out(_U1283_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1284 (
    .in(_U1283_out),
    .clk(clk),
    .out(_U1284_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1285 (
    .in(_U1284_out),
    .clk(clk),
    .out(_U1285_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1286 (
    .in(_U1285_out),
    .clk(clk),
    .out(_U1286_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1287 (
    .in(_U1286_out),
    .clk(clk),
    .out(_U1287_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1288 (
    .in(_U1287_out),
    .clk(clk),
    .out(_U1288_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1289 (
    .in(_U1288_out),
    .clk(clk),
    .out(_U1289_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1290 (
    .in(_U1289_out),
    .clk(clk),
    .out(_U1290_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1291 (
    .in(_U1290_out),
    .clk(clk),
    .out(_U1291_out)
);
_U1292_pt__U1293 _U1292 (
    .in(_U1294_out),
    .out(_U1292_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1294 (
    .in(add_1123_1130_1131_out),
    .clk(clk),
    .out(_U1294_out)
);
_U1295_pt__U1296 _U1295 (
    .in(_U1303_out),
    .out(_U1295_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1297 (
    .in(mul_hw_kernel_global_wrapper_stencil_52_hw_input_global_wrapper_stencil_52_1123_out),
    .clk(clk),
    .out(_U1297_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1298 (
    .in(_U1297_out),
    .clk(clk),
    .out(_U1298_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1299 (
    .in(_U1298_out),
    .clk(clk),
    .out(_U1299_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1300 (
    .in(_U1299_out),
    .clk(clk),
    .out(_U1300_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1301 (
    .in(_U1300_out),
    .clk(clk),
    .out(_U1301_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1302 (
    .in(_U1301_out),
    .clk(clk),
    .out(_U1302_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1303 (
    .in(_U1302_out),
    .clk(clk),
    .out(_U1303_out)
);
_U1304_pt__U1305 _U1304 (
    .in(_U1306_out),
    .out(_U1304_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1306 (
    .in(add_1124_1129_1130_out),
    .clk(clk),
    .out(_U1306_out)
);
_U1307_pt__U1308 _U1307 (
    .in(_U1313_out),
    .out(_U1307_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1309 (
    .in(mul_hw_kernel_global_wrapper_stencil_53_hw_input_global_wrapper_stencil_53_1124_out),
    .clk(clk),
    .out(_U1309_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1310 (
    .in(_U1309_out),
    .clk(clk),
    .out(_U1310_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1311 (
    .in(_U1310_out),
    .clk(clk),
    .out(_U1311_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1312 (
    .in(_U1311_out),
    .clk(clk),
    .out(_U1312_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1313 (
    .in(_U1312_out),
    .clk(clk),
    .out(_U1313_out)
);
_U1314_pt__U1315 _U1314 (
    .in(_U1330_out),
    .out(_U1314_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1316 (
    .in(mul_hw_kernel_global_wrapper_stencil_49_hw_input_global_wrapper_stencil_49_1120_out),
    .clk(clk),
    .out(_U1316_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1317 (
    .in(_U1316_out),
    .clk(clk),
    .out(_U1317_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1318 (
    .in(_U1317_out),
    .clk(clk),
    .out(_U1318_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1319 (
    .in(_U1318_out),
    .clk(clk),
    .out(_U1319_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1320 (
    .in(_U1319_out),
    .clk(clk),
    .out(_U1320_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1321 (
    .in(_U1320_out),
    .clk(clk),
    .out(_U1321_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1322 (
    .in(_U1321_out),
    .clk(clk),
    .out(_U1322_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1323 (
    .in(_U1322_out),
    .clk(clk),
    .out(_U1323_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1324 (
    .in(_U1323_out),
    .clk(clk),
    .out(_U1324_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1325 (
    .in(_U1324_out),
    .clk(clk),
    .out(_U1325_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1326 (
    .in(_U1325_out),
    .clk(clk),
    .out(_U1326_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1327 (
    .in(_U1326_out),
    .clk(clk),
    .out(_U1327_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1328 (
    .in(_U1327_out),
    .clk(clk),
    .out(_U1328_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1329 (
    .in(_U1328_out),
    .clk(clk),
    .out(_U1329_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1330 (
    .in(_U1329_out),
    .clk(clk),
    .out(_U1330_out)
);
_U1331_pt__U1332 _U1331 (
    .in(_U1333_out),
    .out(_U1331_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1333 (
    .in(add_conv_stencil_7_1133_1134_out),
    .clk(clk),
    .out(_U1333_out)
);
_U1334_pt__U1335 _U1334 (
    .in(add_1120_1134_1135_out),
    .out(out_conv_stencil)
);
_U1336_pt__U1337 _U1336 (
    .in(_U1348_out),
    .out(_U1336_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1338 (
    .in(mul_hw_kernel_global_wrapper_stencil_50_hw_input_global_wrapper_stencil_50_1121_out),
    .clk(clk),
    .out(_U1338_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1339 (
    .in(_U1338_out),
    .clk(clk),
    .out(_U1339_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1340 (
    .in(_U1339_out),
    .clk(clk),
    .out(_U1340_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1341 (
    .in(_U1340_out),
    .clk(clk),
    .out(_U1341_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1342 (
    .in(_U1341_out),
    .clk(clk),
    .out(_U1342_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1343 (
    .in(_U1342_out),
    .clk(clk),
    .out(_U1343_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1344 (
    .in(_U1343_out),
    .clk(clk),
    .out(_U1344_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1345 (
    .in(_U1344_out),
    .clk(clk),
    .out(_U1345_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1346 (
    .in(_U1345_out),
    .clk(clk),
    .out(_U1346_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1347 (
    .in(_U1346_out),
    .clk(clk),
    .out(_U1347_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1348 (
    .in(_U1347_out),
    .clk(clk),
    .out(_U1348_out)
);
_U1349_pt__U1350 _U1349 (
    .in(_U1353_out),
    .out(_U1349_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1351 (
    .in(in2_hw_kernel_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U1351_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1352 (
    .in(_U1351_out),
    .clk(clk),
    .out(_U1352_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1353 (
    .in(_U1352_out),
    .clk(clk),
    .out(_U1353_out)
);
_U1354_pt__U1355 _U1354 (
    .in(_U1358_out),
    .out(_U1354_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1356 (
    .in(in1_hw_input_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U1356_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1357 (
    .in(_U1356_out),
    .clk(clk),
    .out(_U1357_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1358 (
    .in(_U1357_out),
    .clk(clk),
    .out(_U1358_out)
);
_U1359_pt__U1360 _U1359 (
    .in(_U1364_out),
    .out(_U1359_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1361 (
    .in(in2_hw_kernel_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U1361_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1362 (
    .in(_U1361_out),
    .clk(clk),
    .out(_U1362_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1363 (
    .in(_U1362_out),
    .clk(clk),
    .out(_U1363_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1364 (
    .in(_U1363_out),
    .clk(clk),
    .out(_U1364_out)
);
_U1365_pt__U1366 _U1365 (
    .in(_U1370_out),
    .out(_U1365_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1367 (
    .in(in1_hw_input_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U1367_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1368 (
    .in(_U1367_out),
    .clk(clk),
    .out(_U1368_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1369 (
    .in(_U1368_out),
    .clk(clk),
    .out(_U1369_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1370 (
    .in(_U1369_out),
    .clk(clk),
    .out(_U1370_out)
);
_U1371_pt__U1372 _U1371 (
    .in(_U1377_out),
    .out(_U1371_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1373 (
    .in(in2_hw_kernel_global_wrapper_stencil[4]),
    .clk(clk),
    .out(_U1373_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1374 (
    .in(_U1373_out),
    .clk(clk),
    .out(_U1374_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1375 (
    .in(_U1374_out),
    .clk(clk),
    .out(_U1375_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1376 (
    .in(_U1375_out),
    .clk(clk),
    .out(_U1376_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1377 (
    .in(_U1376_out),
    .clk(clk),
    .out(_U1377_out)
);
_U1378_pt__U1379 _U1378 (
    .in(_U1385_out),
    .out(_U1378_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1380 (
    .in(in2_hw_kernel_global_wrapper_stencil[5]),
    .clk(clk),
    .out(_U1380_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1381 (
    .in(_U1380_out),
    .clk(clk),
    .out(_U1381_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1382 (
    .in(_U1381_out),
    .clk(clk),
    .out(_U1382_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1383 (
    .in(_U1382_out),
    .clk(clk),
    .out(_U1383_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1384 (
    .in(_U1383_out),
    .clk(clk),
    .out(_U1384_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1385 (
    .in(_U1384_out),
    .clk(clk),
    .out(_U1385_out)
);
_U1386_pt__U1387 _U1386 (
    .in(_U1393_out),
    .out(_U1386_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1388 (
    .in(in1_hw_input_global_wrapper_stencil[5]),
    .clk(clk),
    .out(_U1388_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1389 (
    .in(_U1388_out),
    .clk(clk),
    .out(_U1389_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1390 (
    .in(_U1389_out),
    .clk(clk),
    .out(_U1390_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1391 (
    .in(_U1390_out),
    .clk(clk),
    .out(_U1391_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1392 (
    .in(_U1391_out),
    .clk(clk),
    .out(_U1392_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1393 (
    .in(_U1392_out),
    .clk(clk),
    .out(_U1393_out)
);
_U1394_pt__U1395 _U1394 (
    .in(_U1402_out),
    .out(_U1394_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1396 (
    .in(in2_hw_kernel_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U1396_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1397 (
    .in(_U1396_out),
    .clk(clk),
    .out(_U1397_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1398 (
    .in(_U1397_out),
    .clk(clk),
    .out(_U1398_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1399 (
    .in(_U1398_out),
    .clk(clk),
    .out(_U1399_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1400 (
    .in(_U1399_out),
    .clk(clk),
    .out(_U1400_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1401 (
    .in(_U1400_out),
    .clk(clk),
    .out(_U1401_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1402 (
    .in(_U1401_out),
    .clk(clk),
    .out(_U1402_out)
);
_U1403_pt__U1404 _U1403 (
    .in(_U1411_out),
    .out(_U1403_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1405 (
    .in(in1_hw_input_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U1405_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1406 (
    .in(_U1405_out),
    .clk(clk),
    .out(_U1406_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1407 (
    .in(_U1406_out),
    .clk(clk),
    .out(_U1407_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1408 (
    .in(_U1407_out),
    .clk(clk),
    .out(_U1408_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1409 (
    .in(_U1408_out),
    .clk(clk),
    .out(_U1409_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1410 (
    .in(_U1409_out),
    .clk(clk),
    .out(_U1410_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1411 (
    .in(_U1410_out),
    .clk(clk),
    .out(_U1411_out)
);
_U1412_pt__U1413 _U1412 (
    .in(_U1414_out),
    .out(_U1412_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1414 (
    .in(in2_hw_kernel_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U1414_out)
);
_U1415_pt__U1416 _U1415 (
    .in(_U1417_out),
    .out(_U1415_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1417 (
    .in(in1_hw_input_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U1417_out)
);
_U1418_pt__U1419 _U1418 (
    .in(_U1420_out),
    .out(_U1418_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1420 (
    .in(add_1125_1128_1129_out),
    .clk(clk),
    .out(_U1420_out)
);
_U1421_pt__U1422 _U1421 (
    .in(_U1425_out),
    .out(_U1421_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1423 (
    .in(mul_hw_kernel_global_wrapper_stencil_54_hw_input_global_wrapper_stencil_54_1125_out),
    .clk(clk),
    .out(_U1423_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1424 (
    .in(_U1423_out),
    .clk(clk),
    .out(_U1424_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1425 (
    .in(_U1424_out),
    .clk(clk),
    .out(_U1425_out)
);
_U1426_pt__U1427 _U1426 (
    .in(_U1428_out),
    .out(_U1426_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1428 (
    .in(add_1126_1127_1128_out),
    .clk(clk),
    .out(_U1428_out)
);
_U1429_pt__U1430 _U1429 (
    .in(_U1431_out),
    .out(_U1429_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1431 (
    .in(mul_hw_kernel_global_wrapper_stencil_55_hw_input_global_wrapper_stencil_55_1126_out),
    .clk(clk),
    .out(_U1431_out)
);
_U1432_pt__U1433 _U1432 (
    .in(_U1440_out),
    .out(_U1432_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1434 (
    .in(mul_hw_kernel_global_wrapper_stencil_56_hw_input_global_wrapper_stencil_56_1127_out),
    .clk(clk),
    .out(_U1434_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1435 (
    .in(_U1434_out),
    .clk(clk),
    .out(_U1435_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1436 (
    .in(_U1435_out),
    .clk(clk),
    .out(_U1436_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1437 (
    .in(_U1436_out),
    .clk(clk),
    .out(_U1437_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1438 (
    .in(_U1437_out),
    .clk(clk),
    .out(_U1438_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1439 (
    .in(_U1438_out),
    .clk(clk),
    .out(_U1439_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1440 (
    .in(_U1439_out),
    .clk(clk),
    .out(_U1440_out)
);
assign add_1120_1134_1135_out = 16'(_U1314_out + _U1331_out);
assign add_1121_1132_1133_out = 16'(_U1336_out + _U1275_out);
assign add_1122_1131_1132_out = 16'(_U1281_out + _U1292_out);
assign add_1123_1130_1131_out = 16'(_U1295_out + _U1304_out);
assign add_1124_1129_1130_out = 16'(_U1307_out + _U1418_out);
assign add_1125_1128_1129_out = 16'(_U1421_out + _U1426_out);
assign add_1126_1127_1128_out = 16'(_U1429_out + _U1432_out);
assign add_conv_stencil_7_1133_1134_out = 16'(_U1247_out + _U1278_out);
assign mul_hw_kernel_global_wrapper_stencil_49_hw_input_global_wrapper_stencil_49_1120_out = 16'(_U1263_out * _U1265_out);
assign mul_hw_kernel_global_wrapper_stencil_50_hw_input_global_wrapper_stencil_50_1121_out = 16'(_U1267_out * _U1271_out);
assign mul_hw_kernel_global_wrapper_stencil_51_hw_input_global_wrapper_stencil_51_1122_out = 16'(_U1349_out * _U1354_out);
assign mul_hw_kernel_global_wrapper_stencil_52_hw_input_global_wrapper_stencil_52_1123_out = 16'(_U1359_out * _U1365_out);
assign mul_hw_kernel_global_wrapper_stencil_53_hw_input_global_wrapper_stencil_53_1124_out = 16'(_U1371_out * _U1240_out);
assign mul_hw_kernel_global_wrapper_stencil_54_hw_input_global_wrapper_stencil_54_1125_out = 16'(_U1378_out * _U1386_out);
assign mul_hw_kernel_global_wrapper_stencil_55_hw_input_global_wrapper_stencil_55_1126_out = 16'(_U1394_out * _U1403_out);
assign mul_hw_kernel_global_wrapper_stencil_56_hw_input_global_wrapper_stencil_56_1127_out = 16'(_U1412_out * _U1415_out);
endmodule

module cu_op_hcompute_conv_stencil_14 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_14_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_14_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_14_read[0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[0];
hcompute_conv_stencil_14_pipelined inner_compute (
    .clk(clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_14_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U1238_pt__U1239 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1229_pt__U1230 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1226_pt__U1227 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1221_pt__U1222 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U121_pt__U122 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1214_pt__U1215 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1208_pt__U1209 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1201_pt__U1202 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1197_pt__U1198 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U118_pt__U119 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1181_pt__U1182 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1176_pt__U1177 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1173_pt__U1174 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1170_pt__U1171 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1168_pt__U1169 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1153_pt__U1154 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1150_pt__U1151 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1148_pt__U1149 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1145_pt__U1146 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1134_pt__U1135 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1127_pt__U1128 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1118_pt__U1119 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1115_pt__U1116 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1112_pt__U1113 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1109_pt__U1110 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U10_pt__U11 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_5_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
_U10_pt__U11 _U10 (
    .in(in0_hw_input_stencil[0]),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil_5 (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read[0];
hcompute_hw_input_global_wrapper_stencil_5_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U1098_pt__U1099 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1089_pt__U1090 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1081_pt__U1082 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1073_pt__U1074 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1066_pt__U1067 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1063_pt__U1064 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1054_pt__U1055 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U104_pt__U105 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_8_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U100_out;
wire [15:0] _U101_out;
wire [15:0] _U102_out;
wire [15:0] _U103_out;
wire [15:0] _U104_out;
wire [15:0] _U106_out;
wire [15:0] _U107_out;
wire [15:0] _U108_out;
wire [15:0] _U109_out;
wire [15:0] _U110_out;
wire [15:0] _U111_out;
wire [15:0] _U112_out;
wire [15:0] _U113_out;
wire [15:0] _U114_out;
wire [15:0] _U115_out;
wire [15:0] _U116_out;
wire [15:0] _U117_out;
wire [15:0] _U118_out;
wire [15:0] _U120_out;
wire [15:0] _U121_out;
wire [15:0] _U123_out;
wire [15:0] _U124_out;
wire [15:0] _U126_out;
wire [15:0] _U127_out;
wire [15:0] _U128_out;
wire [15:0] _U129_out;
wire [15:0] _U130_out;
wire [15:0] _U131_out;
wire [15:0] _U132_out;
wire [15:0] _U133_out;
wire [15:0] _U134_out;
wire [15:0] _U135_out;
wire [15:0] _U136_out;
wire [15:0] _U138_out;
wire [15:0] _U139_out;
wire [15:0] _U141_out;
wire [15:0] _U142_out;
wire [15:0] _U143_out;
wire [15:0] _U144_out;
wire [15:0] _U145_out;
wire [15:0] _U146_out;
wire [15:0] _U147_out;
wire [15:0] _U148_out;
wire [15:0] _U149_out;
wire [15:0] _U151_out;
wire [15:0] _U152_out;
wire [15:0] _U154_out;
wire [15:0] _U155_out;
wire [15:0] _U156_out;
wire [15:0] _U157_out;
wire [15:0] _U158_out;
wire [15:0] _U159_out;
wire [15:0] _U160_out;
wire [15:0] _U162_out;
wire [15:0] _U163_out;
wire [15:0] _U165_out;
wire [15:0] _U166_out;
wire [15:0] _U167_out;
wire [15:0] _U168_out;
wire [15:0] _U169_out;
wire [15:0] _U171_out;
wire [15:0] _U172_out;
wire [15:0] _U174_out;
wire [15:0] _U175_out;
wire [15:0] _U176_out;
wire [15:0] _U178_out;
wire [15:0] _U179_out;
wire [15:0] _U181_out;
wire [15:0] _U182_out;
wire [15:0] _U183_out;
wire [15:0] _U184_out;
wire [15:0] _U185_out;
wire [15:0] _U186_out;
wire [15:0] _U187_out;
wire [15:0] _U188_out;
wire [15:0] _U189_out;
wire [15:0] _U190_out;
wire [15:0] _U191_out;
wire [15:0] _U192_out;
wire [15:0] _U193_out;
wire [15:0] _U194_out;
wire [15:0] _U195_out;
wire [15:0] _U197_out;
wire [15:0] _U199_out;
wire [15:0] _U201_out;
wire [15:0] _U202_out;
wire [15:0] _U204_out;
wire [15:0] _U205_out;
wire [15:0] _U207_out;
wire [15:0] _U208_out;
wire [15:0] _U209_out;
wire [15:0] _U211_out;
wire [15:0] _U212_out;
wire [15:0] _U213_out;
wire [15:0] _U215_out;
wire [15:0] _U216_out;
wire [15:0] _U217_out;
wire [15:0] _U218_out;
wire [15:0] _U219_out;
wire [15:0] _U220_out;
wire [15:0] _U221_out;
wire [15:0] _U222_out;
wire [15:0] _U223_out;
wire [15:0] _U224_out;
wire [15:0] _U225_out;
wire [15:0] _U226_out;
wire [15:0] _U227_out;
wire [15:0] _U228_out;
wire [15:0] _U229_out;
wire [15:0] _U230_out;
wire [15:0] _U232_out;
wire [15:0] _U34_out;
wire [15:0] _U36_out;
wire [15:0] _U37_out;
wire [15:0] _U38_out;
wire [15:0] _U39_out;
wire [15:0] _U41_out;
wire [15:0] _U42_out;
wire [15:0] _U43_out;
wire [15:0] _U44_out;
wire [15:0] _U46_out;
wire [15:0] _U47_out;
wire [15:0] _U48_out;
wire [15:0] _U49_out;
wire [15:0] _U50_out;
wire [15:0] _U52_out;
wire [15:0] _U53_out;
wire [15:0] _U54_out;
wire [15:0] _U55_out;
wire [15:0] _U56_out;
wire [15:0] _U58_out;
wire [15:0] _U59_out;
wire [15:0] _U60_out;
wire [15:0] _U61_out;
wire [15:0] _U62_out;
wire [15:0] _U63_out;
wire [15:0] _U65_out;
wire [15:0] _U66_out;
wire [15:0] _U67_out;
wire [15:0] _U68_out;
wire [15:0] _U69_out;
wire [15:0] _U70_out;
wire [15:0] _U72_out;
wire [15:0] _U73_out;
wire [15:0] _U74_out;
wire [15:0] _U75_out;
wire [15:0] _U76_out;
wire [15:0] _U77_out;
wire [15:0] _U78_out;
wire [15:0] _U80_out;
wire [15:0] _U81_out;
wire [15:0] _U82_out;
wire [15:0] _U83_out;
wire [15:0] _U84_out;
wire [15:0] _U85_out;
wire [15:0] _U86_out;
wire [15:0] _U88_out;
wire [15:0] _U89_out;
wire [15:0] _U90_out;
wire [15:0] _U91_out;
wire [15:0] _U92_out;
wire [15:0] _U93_out;
wire [15:0] _U94_out;
wire [15:0] _U95_out;
wire [15:0] _U97_out;
wire [15:0] _U98_out;
wire [15:0] _U99_out;
wire [15:0] add_718_732_733_out;
wire [15:0] add_719_730_731_out;
wire [15:0] add_720_729_730_out;
wire [15:0] add_721_728_729_out;
wire [15:0] add_722_727_728_out;
wire [15:0] add_723_726_727_out;
wire [15:0] add_724_725_726_out;
wire [15:0] add_conv_stencil_1_731_732_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_1_hw_input_global_wrapper_stencil_1_718_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_2_hw_input_global_wrapper_stencil_2_719_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_3_hw_input_global_wrapper_stencil_3_720_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_4_hw_input_global_wrapper_stencil_4_721_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_5_hw_input_global_wrapper_stencil_5_722_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_6_hw_input_global_wrapper_stencil_6_723_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_7_hw_input_global_wrapper_stencil_7_724_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_8_hw_input_global_wrapper_stencil_8_725_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U100 (
    .in(_U99_out),
    .clk(clk),
    .out(_U100_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U101 (
    .in(_U100_out),
    .clk(clk),
    .out(_U101_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U102 (
    .in(_U101_out),
    .clk(clk),
    .out(_U102_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U103 (
    .in(_U102_out),
    .clk(clk),
    .out(_U103_out)
);
_U104_pt__U105 _U104 (
    .in(_U117_out),
    .out(_U104_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U106 (
    .in(mul_hw_kernel_global_wrapper_stencil_2_hw_input_global_wrapper_stencil_2_719_out),
    .clk(clk),
    .out(_U106_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U107 (
    .in(_U106_out),
    .clk(clk),
    .out(_U107_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U108 (
    .in(_U107_out),
    .clk(clk),
    .out(_U108_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U109 (
    .in(_U108_out),
    .clk(clk),
    .out(_U109_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U110 (
    .in(_U109_out),
    .clk(clk),
    .out(_U110_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U111 (
    .in(_U110_out),
    .clk(clk),
    .out(_U111_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U112 (
    .in(_U111_out),
    .clk(clk),
    .out(_U112_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U113 (
    .in(_U112_out),
    .clk(clk),
    .out(_U113_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U114 (
    .in(_U113_out),
    .clk(clk),
    .out(_U114_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U115 (
    .in(_U114_out),
    .clk(clk),
    .out(_U115_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U116 (
    .in(_U115_out),
    .clk(clk),
    .out(_U116_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U117 (
    .in(_U116_out),
    .clk(clk),
    .out(_U117_out)
);
_U118_pt__U119 _U118 (
    .in(_U120_out),
    .out(_U118_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U120 (
    .in(add_720_729_730_out),
    .clk(clk),
    .out(_U120_out)
);
_U121_pt__U122 _U121 (
    .in(_U123_out),
    .out(_U121_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U123 (
    .in(add_719_730_731_out),
    .clk(clk),
    .out(_U123_out)
);
_U124_pt__U125 _U124 (
    .in(_U135_out),
    .out(_U124_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U126 (
    .in(mul_hw_kernel_global_wrapper_stencil_3_hw_input_global_wrapper_stencil_3_720_out),
    .clk(clk),
    .out(_U126_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U127 (
    .in(_U126_out),
    .clk(clk),
    .out(_U127_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U128 (
    .in(_U127_out),
    .clk(clk),
    .out(_U128_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U129 (
    .in(_U128_out),
    .clk(clk),
    .out(_U129_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U130 (
    .in(_U129_out),
    .clk(clk),
    .out(_U130_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U131 (
    .in(_U130_out),
    .clk(clk),
    .out(_U131_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U132 (
    .in(_U131_out),
    .clk(clk),
    .out(_U132_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U133 (
    .in(_U132_out),
    .clk(clk),
    .out(_U133_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U134 (
    .in(_U133_out),
    .clk(clk),
    .out(_U134_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U135 (
    .in(_U134_out),
    .clk(clk),
    .out(_U135_out)
);
_U136_pt__U137 _U136 (
    .in(_U138_out),
    .out(_U136_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U138 (
    .in(add_721_728_729_out),
    .clk(clk),
    .out(_U138_out)
);
_U139_pt__U140 _U139 (
    .in(_U148_out),
    .out(_U139_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U141 (
    .in(mul_hw_kernel_global_wrapper_stencil_4_hw_input_global_wrapper_stencil_4_721_out),
    .clk(clk),
    .out(_U141_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U142 (
    .in(_U141_out),
    .clk(clk),
    .out(_U142_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U143 (
    .in(_U142_out),
    .clk(clk),
    .out(_U143_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U144 (
    .in(_U143_out),
    .clk(clk),
    .out(_U144_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U145 (
    .in(_U144_out),
    .clk(clk),
    .out(_U145_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U146 (
    .in(_U145_out),
    .clk(clk),
    .out(_U146_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U147 (
    .in(_U146_out),
    .clk(clk),
    .out(_U147_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U148 (
    .in(_U147_out),
    .clk(clk),
    .out(_U148_out)
);
_U149_pt__U150 _U149 (
    .in(_U151_out),
    .out(_U149_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U151 (
    .in(add_722_727_728_out),
    .clk(clk),
    .out(_U151_out)
);
_U152_pt__U153 _U152 (
    .in(_U159_out),
    .out(_U152_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U154 (
    .in(mul_hw_kernel_global_wrapper_stencil_5_hw_input_global_wrapper_stencil_5_722_out),
    .clk(clk),
    .out(_U154_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U155 (
    .in(_U154_out),
    .clk(clk),
    .out(_U155_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U156 (
    .in(_U155_out),
    .clk(clk),
    .out(_U156_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U157 (
    .in(_U156_out),
    .clk(clk),
    .out(_U157_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U158 (
    .in(_U157_out),
    .clk(clk),
    .out(_U158_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U159 (
    .in(_U158_out),
    .clk(clk),
    .out(_U159_out)
);
_U160_pt__U161 _U160 (
    .in(_U162_out),
    .out(_U160_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U162 (
    .in(add_723_726_727_out),
    .clk(clk),
    .out(_U162_out)
);
_U163_pt__U164 _U163 (
    .in(_U168_out),
    .out(_U163_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U165 (
    .in(mul_hw_kernel_global_wrapper_stencil_6_hw_input_global_wrapper_stencil_6_723_out),
    .clk(clk),
    .out(_U165_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U166 (
    .in(_U165_out),
    .clk(clk),
    .out(_U166_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U167 (
    .in(_U166_out),
    .clk(clk),
    .out(_U167_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U168 (
    .in(_U167_out),
    .clk(clk),
    .out(_U168_out)
);
_U169_pt__U170 _U169 (
    .in(_U171_out),
    .out(_U169_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U171 (
    .in(add_724_725_726_out),
    .clk(clk),
    .out(_U171_out)
);
_U172_pt__U173 _U172 (
    .in(_U175_out),
    .out(_U172_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U174 (
    .in(mul_hw_kernel_global_wrapper_stencil_7_hw_input_global_wrapper_stencil_7_724_out),
    .clk(clk),
    .out(_U174_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U175 (
    .in(_U174_out),
    .clk(clk),
    .out(_U175_out)
);
_U176_pt__U177 _U176 (
    .in(_U178_out),
    .out(_U176_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U178 (
    .in(mul_hw_kernel_global_wrapper_stencil_8_hw_input_global_wrapper_stencil_8_725_out),
    .clk(clk),
    .out(_U178_out)
);
_U179_pt__U180 _U179 (
    .in(_U194_out),
    .out(_U179_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U181 (
    .in(in0_conv_stencil[0]),
    .clk(clk),
    .out(_U181_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U182 (
    .in(_U181_out),
    .clk(clk),
    .out(_U182_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U183 (
    .in(_U182_out),
    .clk(clk),
    .out(_U183_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U184 (
    .in(_U183_out),
    .clk(clk),
    .out(_U184_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U185 (
    .in(_U184_out),
    .clk(clk),
    .out(_U185_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U186 (
    .in(_U185_out),
    .clk(clk),
    .out(_U186_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U187 (
    .in(_U186_out),
    .clk(clk),
    .out(_U187_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U188 (
    .in(_U187_out),
    .clk(clk),
    .out(_U188_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U189 (
    .in(_U188_out),
    .clk(clk),
    .out(_U189_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U190 (
    .in(_U189_out),
    .clk(clk),
    .out(_U190_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U191 (
    .in(_U190_out),
    .clk(clk),
    .out(_U191_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U192 (
    .in(_U191_out),
    .clk(clk),
    .out(_U192_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U193 (
    .in(_U192_out),
    .clk(clk),
    .out(_U193_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U194 (
    .in(_U193_out),
    .clk(clk),
    .out(_U194_out)
);
_U195_pt__U196 _U195 (
    .in(in2_hw_kernel_global_wrapper_stencil[0]),
    .out(_U195_out)
);
_U197_pt__U198 _U197 (
    .in(in1_hw_input_global_wrapper_stencil[0]),
    .out(_U197_out)
);
_U199_pt__U200 _U199 (
    .in(_U201_out),
    .out(_U199_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U201 (
    .in(in2_hw_kernel_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U201_out)
);
_U202_pt__U203 _U202 (
    .in(_U204_out),
    .out(_U202_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U204 (
    .in(in1_hw_input_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U204_out)
);
_U205_pt__U206 _U205 (
    .in(_U208_out),
    .out(_U205_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U207 (
    .in(in2_hw_kernel_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U207_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U208 (
    .in(_U207_out),
    .clk(clk),
    .out(_U208_out)
);
_U209_pt__U210 _U209 (
    .in(_U212_out),
    .out(_U209_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U211 (
    .in(in1_hw_input_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U211_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U212 (
    .in(_U211_out),
    .clk(clk),
    .out(_U212_out)
);
_U213_pt__U214 _U213 (
    .in(_U229_out),
    .out(_U213_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U215 (
    .in(mul_hw_kernel_global_wrapper_stencil_1_hw_input_global_wrapper_stencil_1_718_out),
    .clk(clk),
    .out(_U215_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U216 (
    .in(_U215_out),
    .clk(clk),
    .out(_U216_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U217 (
    .in(_U216_out),
    .clk(clk),
    .out(_U217_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U218 (
    .in(_U217_out),
    .clk(clk),
    .out(_U218_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U219 (
    .in(_U218_out),
    .clk(clk),
    .out(_U219_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U220 (
    .in(_U219_out),
    .clk(clk),
    .out(_U220_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U221 (
    .in(_U220_out),
    .clk(clk),
    .out(_U221_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U222 (
    .in(_U221_out),
    .clk(clk),
    .out(_U222_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U223 (
    .in(_U222_out),
    .clk(clk),
    .out(_U223_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U224 (
    .in(_U223_out),
    .clk(clk),
    .out(_U224_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U225 (
    .in(_U224_out),
    .clk(clk),
    .out(_U225_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U226 (
    .in(_U225_out),
    .clk(clk),
    .out(_U226_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U227 (
    .in(_U226_out),
    .clk(clk),
    .out(_U227_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U228 (
    .in(_U227_out),
    .clk(clk),
    .out(_U228_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U229 (
    .in(_U228_out),
    .clk(clk),
    .out(_U229_out)
);
_U230_pt__U231 _U230 (
    .in(_U232_out),
    .out(_U230_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U232 (
    .in(add_conv_stencil_1_731_732_out),
    .clk(clk),
    .out(_U232_out)
);
_U233_pt__U234 _U233 (
    .in(add_718_732_733_out),
    .out(out_conv_stencil)
);
_U34_pt__U35 _U34 (
    .in(_U38_out),
    .out(_U34_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U36 (
    .in(in2_hw_kernel_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U36_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U37 (
    .in(_U36_out),
    .clk(clk),
    .out(_U37_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U38 (
    .in(_U37_out),
    .clk(clk),
    .out(_U38_out)
);
_U39_pt__U40 _U39 (
    .in(_U43_out),
    .out(_U39_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U41 (
    .in(in1_hw_input_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U41_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U42 (
    .in(_U41_out),
    .clk(clk),
    .out(_U42_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U43 (
    .in(_U42_out),
    .clk(clk),
    .out(_U43_out)
);
_U44_pt__U45 _U44 (
    .in(_U49_out),
    .out(_U44_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U46 (
    .in(in2_hw_kernel_global_wrapper_stencil[4]),
    .clk(clk),
    .out(_U46_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U47 (
    .in(_U46_out),
    .clk(clk),
    .out(_U47_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U48 (
    .in(_U47_out),
    .clk(clk),
    .out(_U48_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U49 (
    .in(_U48_out),
    .clk(clk),
    .out(_U49_out)
);
_U50_pt__U51 _U50 (
    .in(_U55_out),
    .out(_U50_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U52 (
    .in(in1_hw_input_global_wrapper_stencil[4]),
    .clk(clk),
    .out(_U52_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U53 (
    .in(_U52_out),
    .clk(clk),
    .out(_U53_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U54 (
    .in(_U53_out),
    .clk(clk),
    .out(_U54_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U55 (
    .in(_U54_out),
    .clk(clk),
    .out(_U55_out)
);
_U56_pt__U57 _U56 (
    .in(_U62_out),
    .out(_U56_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U58 (
    .in(in2_hw_kernel_global_wrapper_stencil[5]),
    .clk(clk),
    .out(_U58_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U59 (
    .in(_U58_out),
    .clk(clk),
    .out(_U59_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U60 (
    .in(_U59_out),
    .clk(clk),
    .out(_U60_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U61 (
    .in(_U60_out),
    .clk(clk),
    .out(_U61_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U62 (
    .in(_U61_out),
    .clk(clk),
    .out(_U62_out)
);
_U63_pt__U64 _U63 (
    .in(_U69_out),
    .out(_U63_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U65 (
    .in(in1_hw_input_global_wrapper_stencil[5]),
    .clk(clk),
    .out(_U65_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U66 (
    .in(_U65_out),
    .clk(clk),
    .out(_U66_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U67 (
    .in(_U66_out),
    .clk(clk),
    .out(_U67_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U68 (
    .in(_U67_out),
    .clk(clk),
    .out(_U68_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U69 (
    .in(_U68_out),
    .clk(clk),
    .out(_U69_out)
);
_U70_pt__U71 _U70 (
    .in(_U77_out),
    .out(_U70_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U72 (
    .in(in2_hw_kernel_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U72_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U73 (
    .in(_U72_out),
    .clk(clk),
    .out(_U73_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U74 (
    .in(_U73_out),
    .clk(clk),
    .out(_U74_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U75 (
    .in(_U74_out),
    .clk(clk),
    .out(_U75_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U76 (
    .in(_U75_out),
    .clk(clk),
    .out(_U76_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U77 (
    .in(_U76_out),
    .clk(clk),
    .out(_U77_out)
);
_U78_pt__U79 _U78 (
    .in(_U85_out),
    .out(_U78_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U80 (
    .in(in1_hw_input_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U80_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U81 (
    .in(_U80_out),
    .clk(clk),
    .out(_U81_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U82 (
    .in(_U81_out),
    .clk(clk),
    .out(_U82_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U83 (
    .in(_U82_out),
    .clk(clk),
    .out(_U83_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U84 (
    .in(_U83_out),
    .clk(clk),
    .out(_U84_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U85 (
    .in(_U84_out),
    .clk(clk),
    .out(_U85_out)
);
_U86_pt__U87 _U86 (
    .in(_U94_out),
    .out(_U86_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U88 (
    .in(in2_hw_kernel_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U88_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U89 (
    .in(_U88_out),
    .clk(clk),
    .out(_U89_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U90 (
    .in(_U89_out),
    .clk(clk),
    .out(_U90_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U91 (
    .in(_U90_out),
    .clk(clk),
    .out(_U91_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U92 (
    .in(_U91_out),
    .clk(clk),
    .out(_U92_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U93 (
    .in(_U92_out),
    .clk(clk),
    .out(_U93_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U94 (
    .in(_U93_out),
    .clk(clk),
    .out(_U94_out)
);
_U95_pt__U96 _U95 (
    .in(_U103_out),
    .out(_U95_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U97 (
    .in(in1_hw_input_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U97_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U98 (
    .in(_U97_out),
    .clk(clk),
    .out(_U98_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U99 (
    .in(_U98_out),
    .clk(clk),
    .out(_U99_out)
);
assign add_718_732_733_out = 16'(_U213_out + _U230_out);
assign add_719_730_731_out = 16'(_U104_out + _U118_out);
assign add_720_729_730_out = 16'(_U124_out + _U136_out);
assign add_721_728_729_out = 16'(_U139_out + _U149_out);
assign add_722_727_728_out = 16'(_U152_out + _U160_out);
assign add_723_726_727_out = 16'(_U163_out + _U169_out);
assign add_724_725_726_out = 16'(_U172_out + _U176_out);
assign add_conv_stencil_1_731_732_out = 16'(_U179_out + _U121_out);
assign mul_hw_kernel_global_wrapper_stencil_1_hw_input_global_wrapper_stencil_1_718_out = 16'(_U195_out * _U197_out);
assign mul_hw_kernel_global_wrapper_stencil_2_hw_input_global_wrapper_stencil_2_719_out = 16'(_U199_out * _U202_out);
assign mul_hw_kernel_global_wrapper_stencil_3_hw_input_global_wrapper_stencil_3_720_out = 16'(_U205_out * _U209_out);
assign mul_hw_kernel_global_wrapper_stencil_4_hw_input_global_wrapper_stencil_4_721_out = 16'(_U34_out * _U39_out);
assign mul_hw_kernel_global_wrapper_stencil_5_hw_input_global_wrapper_stencil_5_722_out = 16'(_U44_out * _U50_out);
assign mul_hw_kernel_global_wrapper_stencil_6_hw_input_global_wrapper_stencil_6_723_out = 16'(_U56_out * _U63_out);
assign mul_hw_kernel_global_wrapper_stencil_7_hw_input_global_wrapper_stencil_7_724_out = 16'(_U70_out * _U78_out);
assign mul_hw_kernel_global_wrapper_stencil_8_hw_input_global_wrapper_stencil_8_725_out = 16'(_U86_out * _U95_out);
endmodule

module cu_op_hcompute_conv_stencil_8 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_8_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_8_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_8_read[0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[0];
hcompute_conv_stencil_8_pipelined inner_compute (
    .clk(clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_8_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U1049_pt__U1050 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1043_pt__U1044 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1039_pt__U1040 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_13_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U1039_out;
wire [15:0] _U1041_out;
wire [15:0] _U1042_out;
wire [15:0] _U1043_out;
wire [15:0] _U1045_out;
wire [15:0] _U1046_out;
wire [15:0] _U1047_out;
wire [15:0] _U1048_out;
wire [15:0] _U1049_out;
wire [15:0] _U1051_out;
wire [15:0] _U1052_out;
wire [15:0] _U1053_out;
wire [15:0] _U1054_out;
wire [15:0] _U1056_out;
wire [15:0] _U1057_out;
wire [15:0] _U1058_out;
wire [15:0] _U1059_out;
wire [15:0] _U1060_out;
wire [15:0] _U1061_out;
wire [15:0] _U1062_out;
wire [15:0] _U1063_out;
wire [15:0] _U1065_out;
wire [15:0] _U1066_out;
wire [15:0] _U1068_out;
wire [15:0] _U1069_out;
wire [15:0] _U1070_out;
wire [15:0] _U1071_out;
wire [15:0] _U1072_out;
wire [15:0] _U1073_out;
wire [15:0] _U1075_out;
wire [15:0] _U1076_out;
wire [15:0] _U1077_out;
wire [15:0] _U1078_out;
wire [15:0] _U1079_out;
wire [15:0] _U1080_out;
wire [15:0] _U1081_out;
wire [15:0] _U1083_out;
wire [15:0] _U1084_out;
wire [15:0] _U1085_out;
wire [15:0] _U1086_out;
wire [15:0] _U1087_out;
wire [15:0] _U1088_out;
wire [15:0] _U1089_out;
wire [15:0] _U1091_out;
wire [15:0] _U1092_out;
wire [15:0] _U1093_out;
wire [15:0] _U1094_out;
wire [15:0] _U1095_out;
wire [15:0] _U1096_out;
wire [15:0] _U1097_out;
wire [15:0] _U1098_out;
wire [15:0] _U1100_out;
wire [15:0] _U1101_out;
wire [15:0] _U1102_out;
wire [15:0] _U1103_out;
wire [15:0] _U1104_out;
wire [15:0] _U1105_out;
wire [15:0] _U1106_out;
wire [15:0] _U1107_out;
wire [15:0] _U1108_out;
wire [15:0] _U1109_out;
wire [15:0] _U1111_out;
wire [15:0] _U1112_out;
wire [15:0] _U1114_out;
wire [15:0] _U1115_out;
wire [15:0] _U1117_out;
wire [15:0] _U1118_out;
wire [15:0] _U1120_out;
wire [15:0] _U1121_out;
wire [15:0] _U1122_out;
wire [15:0] _U1123_out;
wire [15:0] _U1124_out;
wire [15:0] _U1125_out;
wire [15:0] _U1126_out;
wire [15:0] _U1127_out;
wire [15:0] _U1129_out;
wire [15:0] _U1130_out;
wire [15:0] _U1131_out;
wire [15:0] _U1132_out;
wire [15:0] _U1133_out;
wire [15:0] _U1134_out;
wire [15:0] _U1136_out;
wire [15:0] _U1137_out;
wire [15:0] _U1138_out;
wire [15:0] _U1139_out;
wire [15:0] _U1140_out;
wire [15:0] _U1141_out;
wire [15:0] _U1142_out;
wire [15:0] _U1143_out;
wire [15:0] _U1144_out;
wire [15:0] _U1145_out;
wire [15:0] _U1147_out;
wire [15:0] _U1150_out;
wire [15:0] _U1152_out;
wire [15:0] _U1153_out;
wire [15:0] _U1155_out;
wire [15:0] _U1156_out;
wire [15:0] _U1157_out;
wire [15:0] _U1158_out;
wire [15:0] _U1159_out;
wire [15:0] _U1160_out;
wire [15:0] _U1161_out;
wire [15:0] _U1162_out;
wire [15:0] _U1163_out;
wire [15:0] _U1164_out;
wire [15:0] _U1165_out;
wire [15:0] _U1166_out;
wire [15:0] _U1167_out;
wire [15:0] _U1168_out;
wire [15:0] _U1170_out;
wire [15:0] _U1172_out;
wire [15:0] _U1173_out;
wire [15:0] _U1175_out;
wire [15:0] _U1176_out;
wire [15:0] _U1178_out;
wire [15:0] _U1179_out;
wire [15:0] _U1180_out;
wire [15:0] _U1181_out;
wire [15:0] _U1183_out;
wire [15:0] _U1184_out;
wire [15:0] _U1185_out;
wire [15:0] _U1186_out;
wire [15:0] _U1187_out;
wire [15:0] _U1188_out;
wire [15:0] _U1189_out;
wire [15:0] _U1190_out;
wire [15:0] _U1191_out;
wire [15:0] _U1192_out;
wire [15:0] _U1193_out;
wire [15:0] _U1194_out;
wire [15:0] _U1195_out;
wire [15:0] _U1196_out;
wire [15:0] _U1197_out;
wire [15:0] _U1199_out;
wire [15:0] _U1200_out;
wire [15:0] _U1201_out;
wire [15:0] _U1203_out;
wire [15:0] _U1204_out;
wire [15:0] _U1205_out;
wire [15:0] _U1206_out;
wire [15:0] _U1207_out;
wire [15:0] _U1208_out;
wire [15:0] _U1210_out;
wire [15:0] _U1211_out;
wire [15:0] _U1212_out;
wire [15:0] _U1213_out;
wire [15:0] _U1214_out;
wire [15:0] _U1216_out;
wire [15:0] _U1217_out;
wire [15:0] _U1218_out;
wire [15:0] _U1219_out;
wire [15:0] _U1220_out;
wire [15:0] _U1221_out;
wire [15:0] _U1223_out;
wire [15:0] _U1224_out;
wire [15:0] _U1225_out;
wire [15:0] _U1226_out;
wire [15:0] _U1228_out;
wire [15:0] _U1229_out;
wire [15:0] _U1231_out;
wire [15:0] _U1232_out;
wire [15:0] _U1233_out;
wire [15:0] _U1234_out;
wire [15:0] _U1235_out;
wire [15:0] _U1236_out;
wire [15:0] _U1237_out;
wire [15:0] _U1238_out;
wire [15:0] add_1053_1067_1068_out;
wire [15:0] add_1054_1065_1066_out;
wire [15:0] add_1055_1064_1065_out;
wire [15:0] add_1056_1063_1064_out;
wire [15:0] add_1057_1062_1063_out;
wire [15:0] add_1058_1061_1062_out;
wire [15:0] add_1059_1060_1061_out;
wire [15:0] add_conv_stencil_6_1066_1067_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_41_hw_input_global_wrapper_stencil_41_1053_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_42_hw_input_global_wrapper_stencil_42_1054_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_43_hw_input_global_wrapper_stencil_43_1055_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_44_hw_input_global_wrapper_stencil_44_1056_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_45_hw_input_global_wrapper_stencil_45_1057_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_46_hw_input_global_wrapper_stencil_46_1058_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_47_hw_input_global_wrapper_stencil_47_1059_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_48_hw_input_global_wrapper_stencil_48_1060_out;
_U1039_pt__U1040 _U1039 (
    .in(_U1042_out),
    .out(_U1039_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1041 (
    .in(in1_hw_input_global_wrapper_stencil[0]),
    .clk(clk),
    .out(_U1041_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1042 (
    .in(_U1041_out),
    .clk(clk),
    .out(_U1042_out)
);
_U1043_pt__U1044 _U1043 (
    .in(_U1048_out),
    .out(_U1043_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1045 (
    .in(in2_hw_kernel_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U1045_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1046 (
    .in(_U1045_out),
    .clk(clk),
    .out(_U1046_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1047 (
    .in(_U1046_out),
    .clk(clk),
    .out(_U1047_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1048 (
    .in(_U1047_out),
    .clk(clk),
    .out(_U1048_out)
);
_U1049_pt__U1050 _U1049 (
    .in(_U1053_out),
    .out(_U1049_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1051 (
    .in(in1_hw_input_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U1051_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1052 (
    .in(_U1051_out),
    .clk(clk),
    .out(_U1052_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1053 (
    .in(_U1052_out),
    .clk(clk),
    .out(_U1053_out)
);
_U1054_pt__U1055 _U1054 (
    .in(_U1062_out),
    .out(_U1054_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1056 (
    .in(mul_hw_kernel_global_wrapper_stencil_43_hw_input_global_wrapper_stencil_43_1055_out),
    .clk(clk),
    .out(_U1056_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1057 (
    .in(_U1056_out),
    .clk(clk),
    .out(_U1057_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1058 (
    .in(_U1057_out),
    .clk(clk),
    .out(_U1058_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1059 (
    .in(_U1058_out),
    .clk(clk),
    .out(_U1059_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1060 (
    .in(_U1059_out),
    .clk(clk),
    .out(_U1060_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1061 (
    .in(_U1060_out),
    .clk(clk),
    .out(_U1061_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1062 (
    .in(_U1061_out),
    .clk(clk),
    .out(_U1062_out)
);
_U1063_pt__U1064 _U1063 (
    .in(_U1065_out),
    .out(_U1063_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1065 (
    .in(add_1056_1063_1064_out),
    .clk(clk),
    .out(_U1065_out)
);
_U1066_pt__U1067 _U1066 (
    .in(_U1072_out),
    .out(_U1066_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1068 (
    .in(in1_hw_input_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U1068_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1069 (
    .in(_U1068_out),
    .clk(clk),
    .out(_U1069_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1070 (
    .in(_U1069_out),
    .clk(clk),
    .out(_U1070_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1071 (
    .in(_U1070_out),
    .clk(clk),
    .out(_U1071_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1072 (
    .in(_U1071_out),
    .clk(clk),
    .out(_U1072_out)
);
_U1073_pt__U1074 _U1073 (
    .in(_U1080_out),
    .out(_U1073_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1075 (
    .in(in2_hw_kernel_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U1075_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1076 (
    .in(_U1075_out),
    .clk(clk),
    .out(_U1076_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1077 (
    .in(_U1076_out),
    .clk(clk),
    .out(_U1077_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1078 (
    .in(_U1077_out),
    .clk(clk),
    .out(_U1078_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1079 (
    .in(_U1078_out),
    .clk(clk),
    .out(_U1079_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1080 (
    .in(_U1079_out),
    .clk(clk),
    .out(_U1080_out)
);
_U1081_pt__U1082 _U1081 (
    .in(_U1088_out),
    .out(_U1081_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1083 (
    .in(in1_hw_input_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U1083_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1084 (
    .in(_U1083_out),
    .clk(clk),
    .out(_U1084_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1085 (
    .in(_U1084_out),
    .clk(clk),
    .out(_U1085_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1086 (
    .in(_U1085_out),
    .clk(clk),
    .out(_U1086_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1087 (
    .in(_U1086_out),
    .clk(clk),
    .out(_U1087_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1088 (
    .in(_U1087_out),
    .clk(clk),
    .out(_U1088_out)
);
_U1089_pt__U1090 _U1089 (
    .in(_U1097_out),
    .out(_U1089_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1091 (
    .in(in2_hw_kernel_global_wrapper_stencil[4]),
    .clk(clk),
    .out(_U1091_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1092 (
    .in(_U1091_out),
    .clk(clk),
    .out(_U1092_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1093 (
    .in(_U1092_out),
    .clk(clk),
    .out(_U1093_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1094 (
    .in(_U1093_out),
    .clk(clk),
    .out(_U1094_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1095 (
    .in(_U1094_out),
    .clk(clk),
    .out(_U1095_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1096 (
    .in(_U1095_out),
    .clk(clk),
    .out(_U1096_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1097 (
    .in(_U1096_out),
    .clk(clk),
    .out(_U1097_out)
);
_U1098_pt__U1099 _U1098 (
    .in(_U1108_out),
    .out(_U1098_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1100 (
    .in(mul_hw_kernel_global_wrapper_stencil_46_hw_input_global_wrapper_stencil_46_1058_out),
    .clk(clk),
    .out(_U1100_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1101 (
    .in(_U1100_out),
    .clk(clk),
    .out(_U1101_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1102 (
    .in(_U1101_out),
    .clk(clk),
    .out(_U1102_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1103 (
    .in(_U1102_out),
    .clk(clk),
    .out(_U1103_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1104 (
    .in(_U1103_out),
    .clk(clk),
    .out(_U1104_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1105 (
    .in(_U1104_out),
    .clk(clk),
    .out(_U1105_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1106 (
    .in(_U1105_out),
    .clk(clk),
    .out(_U1106_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1107 (
    .in(_U1106_out),
    .clk(clk),
    .out(_U1107_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1108 (
    .in(_U1107_out),
    .clk(clk),
    .out(_U1108_out)
);
_U1109_pt__U1110 _U1109 (
    .in(_U1111_out),
    .out(_U1109_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1111 (
    .in(add_1059_1060_1061_out),
    .clk(clk),
    .out(_U1111_out)
);
_U1112_pt__U1113 _U1112 (
    .in(_U1114_out),
    .out(_U1112_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1114 (
    .in(add_1055_1064_1065_out),
    .clk(clk),
    .out(_U1114_out)
);
_U1115_pt__U1116 _U1115 (
    .in(_U1117_out),
    .out(_U1115_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1117 (
    .in(add_1054_1065_1066_out),
    .clk(clk),
    .out(_U1117_out)
);
_U1118_pt__U1119 _U1118 (
    .in(_U1126_out),
    .out(_U1118_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1120 (
    .in(mul_hw_kernel_global_wrapper_stencil_47_hw_input_global_wrapper_stencil_47_1059_out),
    .clk(clk),
    .out(_U1120_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1121 (
    .in(_U1120_out),
    .clk(clk),
    .out(_U1121_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1122 (
    .in(_U1121_out),
    .clk(clk),
    .out(_U1122_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1123 (
    .in(_U1122_out),
    .clk(clk),
    .out(_U1123_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1124 (
    .in(_U1123_out),
    .clk(clk),
    .out(_U1124_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1125 (
    .in(_U1124_out),
    .clk(clk),
    .out(_U1125_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1126 (
    .in(_U1125_out),
    .clk(clk),
    .out(_U1126_out)
);
_U1127_pt__U1128 _U1127 (
    .in(_U1133_out),
    .out(_U1127_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1129 (
    .in(mul_hw_kernel_global_wrapper_stencil_48_hw_input_global_wrapper_stencil_48_1060_out),
    .clk(clk),
    .out(_U1129_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1130 (
    .in(_U1129_out),
    .clk(clk),
    .out(_U1130_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1131 (
    .in(_U1130_out),
    .clk(clk),
    .out(_U1131_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1132 (
    .in(_U1131_out),
    .clk(clk),
    .out(_U1132_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1133 (
    .in(_U1132_out),
    .clk(clk),
    .out(_U1133_out)
);
_U1134_pt__U1135 _U1134 (
    .in(_U1144_out),
    .out(_U1134_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1136 (
    .in(mul_hw_kernel_global_wrapper_stencil_42_hw_input_global_wrapper_stencil_42_1054_out),
    .clk(clk),
    .out(_U1136_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1137 (
    .in(_U1136_out),
    .clk(clk),
    .out(_U1137_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1138 (
    .in(_U1137_out),
    .clk(clk),
    .out(_U1138_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1139 (
    .in(_U1138_out),
    .clk(clk),
    .out(_U1139_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1140 (
    .in(_U1139_out),
    .clk(clk),
    .out(_U1140_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1141 (
    .in(_U1140_out),
    .clk(clk),
    .out(_U1141_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1142 (
    .in(_U1141_out),
    .clk(clk),
    .out(_U1142_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1143 (
    .in(_U1142_out),
    .clk(clk),
    .out(_U1143_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1144 (
    .in(_U1143_out),
    .clk(clk),
    .out(_U1144_out)
);
_U1145_pt__U1146 _U1145 (
    .in(_U1147_out),
    .out(_U1145_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1147 (
    .in(add_conv_stencil_6_1066_1067_out),
    .clk(clk),
    .out(_U1147_out)
);
_U1148_pt__U1149 _U1148 (
    .in(add_1053_1067_1068_out),
    .out(out_conv_stencil)
);
_U1150_pt__U1151 _U1150 (
    .in(_U1152_out),
    .out(_U1150_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1152 (
    .in(add_1057_1062_1063_out),
    .clk(clk),
    .out(_U1152_out)
);
_U1153_pt__U1154 _U1153 (
    .in(_U1167_out),
    .out(_U1153_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1155 (
    .in(mul_hw_kernel_global_wrapper_stencil_41_hw_input_global_wrapper_stencil_41_1053_out),
    .clk(clk),
    .out(_U1155_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1156 (
    .in(_U1155_out),
    .clk(clk),
    .out(_U1156_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1157 (
    .in(_U1156_out),
    .clk(clk),
    .out(_U1157_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1158 (
    .in(_U1157_out),
    .clk(clk),
    .out(_U1158_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1159 (
    .in(_U1158_out),
    .clk(clk),
    .out(_U1159_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1160 (
    .in(_U1159_out),
    .clk(clk),
    .out(_U1160_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1161 (
    .in(_U1160_out),
    .clk(clk),
    .out(_U1161_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1162 (
    .in(_U1161_out),
    .clk(clk),
    .out(_U1162_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1163 (
    .in(_U1162_out),
    .clk(clk),
    .out(_U1163_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1164 (
    .in(_U1163_out),
    .clk(clk),
    .out(_U1164_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1165 (
    .in(_U1164_out),
    .clk(clk),
    .out(_U1165_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1166 (
    .in(_U1165_out),
    .clk(clk),
    .out(_U1166_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1167 (
    .in(_U1166_out),
    .clk(clk),
    .out(_U1167_out)
);
_U1168_pt__U1169 _U1168 (
    .in(in1_hw_input_global_wrapper_stencil[5]),
    .out(_U1168_out)
);
_U1170_pt__U1171 _U1170 (
    .in(_U1172_out),
    .out(_U1170_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1172 (
    .in(in2_hw_kernel_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U1172_out)
);
_U1173_pt__U1174 _U1173 (
    .in(_U1175_out),
    .out(_U1173_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1175 (
    .in(in1_hw_input_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U1175_out)
);
_U1176_pt__U1177 _U1176 (
    .in(_U1180_out),
    .out(_U1176_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1178 (
    .in(in2_hw_kernel_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U1178_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1179 (
    .in(_U1178_out),
    .clk(clk),
    .out(_U1179_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1180 (
    .in(_U1179_out),
    .clk(clk),
    .out(_U1180_out)
);
_U1181_pt__U1182 _U1181 (
    .in(_U1196_out),
    .out(_U1181_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1183 (
    .in(in0_conv_stencil[0]),
    .clk(clk),
    .out(_U1183_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1184 (
    .in(_U1183_out),
    .clk(clk),
    .out(_U1184_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1185 (
    .in(_U1184_out),
    .clk(clk),
    .out(_U1185_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1186 (
    .in(_U1185_out),
    .clk(clk),
    .out(_U1186_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1187 (
    .in(_U1186_out),
    .clk(clk),
    .out(_U1187_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1188 (
    .in(_U1187_out),
    .clk(clk),
    .out(_U1188_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1189 (
    .in(_U1188_out),
    .clk(clk),
    .out(_U1189_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1190 (
    .in(_U1189_out),
    .clk(clk),
    .out(_U1190_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1191 (
    .in(_U1190_out),
    .clk(clk),
    .out(_U1191_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1192 (
    .in(_U1191_out),
    .clk(clk),
    .out(_U1192_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1193 (
    .in(_U1192_out),
    .clk(clk),
    .out(_U1193_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1194 (
    .in(_U1193_out),
    .clk(clk),
    .out(_U1194_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1195 (
    .in(_U1194_out),
    .clk(clk),
    .out(_U1195_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1196 (
    .in(_U1195_out),
    .clk(clk),
    .out(_U1196_out)
);
_U1197_pt__U1198 _U1197 (
    .in(_U1200_out),
    .out(_U1197_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1199 (
    .in(in2_hw_kernel_global_wrapper_stencil[0]),
    .clk(clk),
    .out(_U1199_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1200 (
    .in(_U1199_out),
    .clk(clk),
    .out(_U1200_out)
);
_U1201_pt__U1202 _U1201 (
    .in(_U1207_out),
    .out(_U1201_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1203 (
    .in(mul_hw_kernel_global_wrapper_stencil_44_hw_input_global_wrapper_stencil_44_1056_out),
    .clk(clk),
    .out(_U1203_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1204 (
    .in(_U1203_out),
    .clk(clk),
    .out(_U1204_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1205 (
    .in(_U1204_out),
    .clk(clk),
    .out(_U1205_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1206 (
    .in(_U1205_out),
    .clk(clk),
    .out(_U1206_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1207 (
    .in(_U1206_out),
    .clk(clk),
    .out(_U1207_out)
);
_U1208_pt__U1209 _U1208 (
    .in(_U1213_out),
    .out(_U1208_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1210 (
    .in(in1_hw_input_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U1210_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1211 (
    .in(_U1210_out),
    .clk(clk),
    .out(_U1211_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1212 (
    .in(_U1211_out),
    .clk(clk),
    .out(_U1212_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1213 (
    .in(_U1212_out),
    .clk(clk),
    .out(_U1213_out)
);
_U1214_pt__U1215 _U1214 (
    .in(_U1220_out),
    .out(_U1214_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1216 (
    .in(in2_hw_kernel_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U1216_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1217 (
    .in(_U1216_out),
    .clk(clk),
    .out(_U1217_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1218 (
    .in(_U1217_out),
    .clk(clk),
    .out(_U1218_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1219 (
    .in(_U1218_out),
    .clk(clk),
    .out(_U1219_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1220 (
    .in(_U1219_out),
    .clk(clk),
    .out(_U1220_out)
);
_U1221_pt__U1222 _U1221 (
    .in(_U1225_out),
    .out(_U1221_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1223 (
    .in(mul_hw_kernel_global_wrapper_stencil_45_hw_input_global_wrapper_stencil_45_1057_out),
    .clk(clk),
    .out(_U1223_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1224 (
    .in(_U1223_out),
    .clk(clk),
    .out(_U1224_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1225 (
    .in(_U1224_out),
    .clk(clk),
    .out(_U1225_out)
);
_U1226_pt__U1227 _U1226 (
    .in(_U1228_out),
    .out(_U1226_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1228 (
    .in(add_1058_1061_1062_out),
    .clk(clk),
    .out(_U1228_out)
);
_U1229_pt__U1230 _U1229 (
    .in(_U1237_out),
    .out(_U1229_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1231 (
    .in(in1_hw_input_global_wrapper_stencil[4]),
    .clk(clk),
    .out(_U1231_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1232 (
    .in(_U1231_out),
    .clk(clk),
    .out(_U1232_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1233 (
    .in(_U1232_out),
    .clk(clk),
    .out(_U1233_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1234 (
    .in(_U1233_out),
    .clk(clk),
    .out(_U1234_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1235 (
    .in(_U1234_out),
    .clk(clk),
    .out(_U1235_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1236 (
    .in(_U1235_out),
    .clk(clk),
    .out(_U1236_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1237 (
    .in(_U1236_out),
    .clk(clk),
    .out(_U1237_out)
);
_U1238_pt__U1239 _U1238 (
    .in(in2_hw_kernel_global_wrapper_stencil[5]),
    .out(_U1238_out)
);
assign add_1053_1067_1068_out = 16'(_U1153_out + _U1145_out);
assign add_1054_1065_1066_out = 16'(_U1134_out + _U1112_out);
assign add_1055_1064_1065_out = 16'(_U1054_out + _U1063_out);
assign add_1056_1063_1064_out = 16'(_U1201_out + _U1150_out);
assign add_1057_1062_1063_out = 16'(_U1221_out + _U1226_out);
assign add_1058_1061_1062_out = 16'(_U1098_out + _U1109_out);
assign add_1059_1060_1061_out = 16'(_U1118_out + _U1127_out);
assign add_conv_stencil_6_1066_1067_out = 16'(_U1181_out + _U1115_out);
assign mul_hw_kernel_global_wrapper_stencil_41_hw_input_global_wrapper_stencil_41_1053_out = 16'(_U1197_out * _U1039_out);
assign mul_hw_kernel_global_wrapper_stencil_42_hw_input_global_wrapper_stencil_42_1054_out = 16'(_U1043_out * _U1208_out);
assign mul_hw_kernel_global_wrapper_stencil_43_hw_input_global_wrapper_stencil_43_1055_out = 16'(_U1214_out * _U1066_out);
assign mul_hw_kernel_global_wrapper_stencil_44_hw_input_global_wrapper_stencil_44_1056_out = 16'(_U1073_out * _U1081_out);
assign mul_hw_kernel_global_wrapper_stencil_45_hw_input_global_wrapper_stencil_45_1057_out = 16'(_U1089_out * _U1229_out);
assign mul_hw_kernel_global_wrapper_stencil_46_hw_input_global_wrapper_stencil_46_1058_out = 16'(_U1238_out * _U1168_out);
assign mul_hw_kernel_global_wrapper_stencil_47_hw_input_global_wrapper_stencil_47_1059_out = 16'(_U1170_out * _U1173_out);
assign mul_hw_kernel_global_wrapper_stencil_48_hw_input_global_wrapper_stencil_48_1060_out = 16'(_U1176_out * _U1049_out);
endmodule

module cu_op_hcompute_conv_stencil_13 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_13_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_13_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_13_read[0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[0];
hcompute_conv_stencil_13_pipelined inner_compute (
    .clk(clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_13_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U1030_pt__U1031 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1028_pt__U1029 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1021_pt__U1022 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1012_pt__U1013 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1010_pt__U1011 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1005_pt__U1006 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1002_pt__U1003 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_12_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U1000_out;
wire [15:0] _U1001_out;
wire [15:0] _U1002_out;
wire [15:0] _U1004_out;
wire [15:0] _U1005_out;
wire [15:0] _U1007_out;
wire [15:0] _U1008_out;
wire [15:0] _U1009_out;
wire [15:0] _U1010_out;
wire [15:0] _U1012_out;
wire [15:0] _U1014_out;
wire [15:0] _U1015_out;
wire [15:0] _U1016_out;
wire [15:0] _U1017_out;
wire [15:0] _U1018_out;
wire [15:0] _U1019_out;
wire [15:0] _U1020_out;
wire [15:0] _U1021_out;
wire [15:0] _U1023_out;
wire [15:0] _U1024_out;
wire [15:0] _U1025_out;
wire [15:0] _U1026_out;
wire [15:0] _U1027_out;
wire [15:0] _U1028_out;
wire [15:0] _U1030_out;
wire [15:0] _U1032_out;
wire [15:0] _U1033_out;
wire [15:0] _U1034_out;
wire [15:0] _U1035_out;
wire [15:0] _U1036_out;
wire [15:0] _U1037_out;
wire [15:0] _U1038_out;
wire [15:0] _U840_out;
wire [15:0] _U842_out;
wire [15:0] _U843_out;
wire [15:0] _U844_out;
wire [15:0] _U845_out;
wire [15:0] _U846_out;
wire [15:0] _U847_out;
wire [15:0] _U848_out;
wire [15:0] _U849_out;
wire [15:0] _U850_out;
wire [15:0] _U851_out;
wire [15:0] _U852_out;
wire [15:0] _U853_out;
wire [15:0] _U854_out;
wire [15:0] _U855_out;
wire [15:0] _U856_out;
wire [15:0] _U858_out;
wire [15:0] _U859_out;
wire [15:0] _U861_out;
wire [15:0] _U862_out;
wire [15:0] _U863_out;
wire [15:0] _U864_out;
wire [15:0] _U866_out;
wire [15:0] _U867_out;
wire [15:0] _U868_out;
wire [15:0] _U869_out;
wire [15:0] _U870_out;
wire [15:0] _U871_out;
wire [15:0] _U872_out;
wire [15:0] _U873_out;
wire [15:0] _U874_out;
wire [15:0] _U875_out;
wire [15:0] _U876_out;
wire [15:0] _U878_out;
wire [15:0] _U879_out;
wire [15:0] _U880_out;
wire [15:0] _U881_out;
wire [15:0] _U882_out;
wire [15:0] _U884_out;
wire [15:0] _U885_out;
wire [15:0] _U887_out;
wire [15:0] _U888_out;
wire [15:0] _U890_out;
wire [15:0] _U891_out;
wire [15:0] _U893_out;
wire [15:0] _U894_out;
wire [15:0] _U895_out;
wire [15:0] _U896_out;
wire [15:0] _U897_out;
wire [15:0] _U898_out;
wire [15:0] _U899_out;
wire [15:0] _U901_out;
wire [15:0] _U902_out;
wire [15:0] _U904_out;
wire [15:0] _U905_out;
wire [15:0] _U907_out;
wire [15:0] _U908_out;
wire [15:0] _U909_out;
wire [15:0] _U910_out;
wire [15:0] _U911_out;
wire [15:0] _U912_out;
wire [15:0] _U913_out;
wire [15:0] _U914_out;
wire [15:0] _U916_out;
wire [15:0] _U917_out;
wire [15:0] _U919_out;
wire [15:0] _U920_out;
wire [15:0] _U921_out;
wire [15:0] _U922_out;
wire [15:0] _U923_out;
wire [15:0] _U924_out;
wire [15:0] _U925_out;
wire [15:0] _U926_out;
wire [15:0] _U927_out;
wire [15:0] _U928_out;
wire [15:0] _U929_out;
wire [15:0] _U930_out;
wire [15:0] _U931_out;
wire [15:0] _U932_out;
wire [15:0] _U934_out;
wire [15:0] _U935_out;
wire [15:0] _U936_out;
wire [15:0] _U937_out;
wire [15:0] _U938_out;
wire [15:0] _U940_out;
wire [15:0] _U941_out;
wire [15:0] _U942_out;
wire [15:0] _U943_out;
wire [15:0] _U944_out;
wire [15:0] _U945_out;
wire [15:0] _U946_out;
wire [15:0] _U948_out;
wire [15:0] _U949_out;
wire [15:0] _U951_out;
wire [15:0] _U952_out;
wire [15:0] _U953_out;
wire [15:0] _U954_out;
wire [15:0] _U955_out;
wire [15:0] _U956_out;
wire [15:0] _U957_out;
wire [15:0] _U959_out;
wire [15:0] _U960_out;
wire [15:0] _U961_out;
wire [15:0] _U963_out;
wire [15:0] _U964_out;
wire [15:0] _U965_out;
wire [15:0] _U967_out;
wire [15:0] _U968_out;
wire [15:0] _U969_out;
wire [15:0] _U970_out;
wire [15:0] _U971_out;
wire [15:0] _U972_out;
wire [15:0] _U973_out;
wire [15:0] _U975_out;
wire [15:0] _U976_out;
wire [15:0] _U977_out;
wire [15:0] _U978_out;
wire [15:0] _U979_out;
wire [15:0] _U980_out;
wire [15:0] _U981_out;
wire [15:0] _U982_out;
wire [15:0] _U983_out;
wire [15:0] _U984_out;
wire [15:0] _U985_out;
wire [15:0] _U986_out;
wire [15:0] _U987_out;
wire [15:0] _U989_out;
wire [15:0] _U990_out;
wire [15:0] _U992_out;
wire [15:0] _U993_out;
wire [15:0] _U994_out;
wire [15:0] _U995_out;
wire [15:0] _U996_out;
wire [15:0] _U997_out;
wire [15:0] _U999_out;
wire [15:0] add_986_1000_1001_out;
wire [15:0] add_987_998_999_out;
wire [15:0] add_988_997_998_out;
wire [15:0] add_989_996_997_out;
wire [15:0] add_990_995_996_out;
wire [15:0] add_991_994_995_out;
wire [15:0] add_992_993_994_out;
wire [15:0] add_conv_stencil_5_999_1000_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_33_hw_input_global_wrapper_stencil_33_986_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_34_hw_input_global_wrapper_stencil_34_987_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_35_hw_input_global_wrapper_stencil_35_988_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_36_hw_input_global_wrapper_stencil_36_989_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_37_hw_input_global_wrapper_stencil_37_990_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_38_hw_input_global_wrapper_stencil_38_991_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_39_hw_input_global_wrapper_stencil_39_992_out;
wire [15:0] mul_hw_kernel_global_wrapper_stencil_40_hw_input_global_wrapper_stencil_40_993_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1000 (
    .in(_U999_out),
    .clk(clk),
    .out(_U1000_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1001 (
    .in(_U1000_out),
    .clk(clk),
    .out(_U1001_out)
);
_U1002_pt__U1003 _U1002 (
    .in(_U1004_out),
    .out(_U1002_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1004 (
    .in(mul_hw_kernel_global_wrapper_stencil_39_hw_input_global_wrapper_stencil_39_992_out),
    .clk(clk),
    .out(_U1004_out)
);
_U1005_pt__U1006 _U1005 (
    .in(_U1009_out),
    .out(_U1005_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1007 (
    .in(in2_hw_kernel_global_wrapper_stencil[5]),
    .clk(clk),
    .out(_U1007_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1008 (
    .in(_U1007_out),
    .clk(clk),
    .out(_U1008_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1009 (
    .in(_U1008_out),
    .clk(clk),
    .out(_U1009_out)
);
_U1010_pt__U1011 _U1010 (
    .in(in2_hw_kernel_global_wrapper_stencil[4]),
    .out(_U1010_out)
);
_U1012_pt__U1013 _U1012 (
    .in(_U1020_out),
    .out(_U1012_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1014 (
    .in(in2_hw_kernel_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U1014_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1015 (
    .in(_U1014_out),
    .clk(clk),
    .out(_U1015_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1016 (
    .in(_U1015_out),
    .clk(clk),
    .out(_U1016_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1017 (
    .in(_U1016_out),
    .clk(clk),
    .out(_U1017_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1018 (
    .in(_U1017_out),
    .clk(clk),
    .out(_U1018_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1019 (
    .in(_U1018_out),
    .clk(clk),
    .out(_U1019_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1020 (
    .in(_U1019_out),
    .clk(clk),
    .out(_U1020_out)
);
_U1021_pt__U1022 _U1021 (
    .in(_U1027_out),
    .out(_U1021_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1023 (
    .in(in1_hw_input_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U1023_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1024 (
    .in(_U1023_out),
    .clk(clk),
    .out(_U1024_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1025 (
    .in(_U1024_out),
    .clk(clk),
    .out(_U1025_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1026 (
    .in(_U1025_out),
    .clk(clk),
    .out(_U1026_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1027 (
    .in(_U1026_out),
    .clk(clk),
    .out(_U1027_out)
);
_U1028_pt__U1029 _U1028 (
    .in(in1_hw_input_global_wrapper_stencil[4]),
    .out(_U1028_out)
);
_U1030_pt__U1031 _U1030 (
    .in(_U1038_out),
    .out(_U1030_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1032 (
    .in(in1_hw_input_global_wrapper_stencil[6]),
    .clk(clk),
    .out(_U1032_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1033 (
    .in(_U1032_out),
    .clk(clk),
    .out(_U1033_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1034 (
    .in(_U1033_out),
    .clk(clk),
    .out(_U1034_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1035 (
    .in(_U1034_out),
    .clk(clk),
    .out(_U1035_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1036 (
    .in(_U1035_out),
    .clk(clk),
    .out(_U1036_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1037 (
    .in(_U1036_out),
    .clk(clk),
    .out(_U1037_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1038 (
    .in(_U1037_out),
    .clk(clk),
    .out(_U1038_out)
);
_U838_pt__U839 _U838 (
    .in(add_986_1000_1001_out),
    .out(out_conv_stencil)
);
_U840_pt__U841 _U840 (
    .in(_U855_out),
    .out(_U840_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U842 (
    .in(in0_conv_stencil[0]),
    .clk(clk),
    .out(_U842_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U843 (
    .in(_U842_out),
    .clk(clk),
    .out(_U843_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U844 (
    .in(_U843_out),
    .clk(clk),
    .out(_U844_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U845 (
    .in(_U844_out),
    .clk(clk),
    .out(_U845_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U846 (
    .in(_U845_out),
    .clk(clk),
    .out(_U846_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U847 (
    .in(_U846_out),
    .clk(clk),
    .out(_U847_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U848 (
    .in(_U847_out),
    .clk(clk),
    .out(_U848_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U849 (
    .in(_U848_out),
    .clk(clk),
    .out(_U849_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U850 (
    .in(_U849_out),
    .clk(clk),
    .out(_U850_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U851 (
    .in(_U850_out),
    .clk(clk),
    .out(_U851_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U852 (
    .in(_U851_out),
    .clk(clk),
    .out(_U852_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U853 (
    .in(_U852_out),
    .clk(clk),
    .out(_U853_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U854 (
    .in(_U853_out),
    .clk(clk),
    .out(_U854_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U855 (
    .in(_U854_out),
    .clk(clk),
    .out(_U855_out)
);
_U856_pt__U857 _U856 (
    .in(_U858_out),
    .out(_U856_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U858 (
    .in(add_989_996_997_out),
    .clk(clk),
    .out(_U858_out)
);
_U859_pt__U860 _U859 (
    .in(_U863_out),
    .out(_U859_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U861 (
    .in(mul_hw_kernel_global_wrapper_stencil_40_hw_input_global_wrapper_stencil_40_993_out),
    .clk(clk),
    .out(_U861_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U862 (
    .in(_U861_out),
    .clk(clk),
    .out(_U862_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U863 (
    .in(_U862_out),
    .clk(clk),
    .out(_U863_out)
);
_U864_pt__U865 _U864 (
    .in(_U875_out),
    .out(_U864_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U866 (
    .in(mul_hw_kernel_global_wrapper_stencil_37_hw_input_global_wrapper_stencil_37_990_out),
    .clk(clk),
    .out(_U866_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U867 (
    .in(_U866_out),
    .clk(clk),
    .out(_U867_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U868 (
    .in(_U867_out),
    .clk(clk),
    .out(_U868_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U869 (
    .in(_U868_out),
    .clk(clk),
    .out(_U869_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U870 (
    .in(_U869_out),
    .clk(clk),
    .out(_U870_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U871 (
    .in(_U870_out),
    .clk(clk),
    .out(_U871_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U872 (
    .in(_U871_out),
    .clk(clk),
    .out(_U872_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U873 (
    .in(_U872_out),
    .clk(clk),
    .out(_U873_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U874 (
    .in(_U873_out),
    .clk(clk),
    .out(_U874_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U875 (
    .in(_U874_out),
    .clk(clk),
    .out(_U875_out)
);
_U876_pt__U877 _U876 (
    .in(_U881_out),
    .out(_U876_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U878 (
    .in(in2_hw_kernel_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U878_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U879 (
    .in(_U878_out),
    .clk(clk),
    .out(_U879_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U880 (
    .in(_U879_out),
    .clk(clk),
    .out(_U880_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U881 (
    .in(_U880_out),
    .clk(clk),
    .out(_U881_out)
);
_U882_pt__U883 _U882 (
    .in(_U884_out),
    .out(_U882_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U884 (
    .in(add_991_994_995_out),
    .clk(clk),
    .out(_U884_out)
);
_U885_pt__U886 _U885 (
    .in(_U887_out),
    .out(_U885_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U887 (
    .in(add_992_993_994_out),
    .clk(clk),
    .out(_U887_out)
);
_U888_pt__U889 _U888 (
    .in(_U890_out),
    .out(_U888_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U890 (
    .in(add_990_995_996_out),
    .clk(clk),
    .out(_U890_out)
);
_U891_pt__U892 _U891 (
    .in(_U898_out),
    .out(_U891_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U893 (
    .in(mul_hw_kernel_global_wrapper_stencil_38_hw_input_global_wrapper_stencil_38_991_out),
    .clk(clk),
    .out(_U893_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U894 (
    .in(_U893_out),
    .clk(clk),
    .out(_U894_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U895 (
    .in(_U894_out),
    .clk(clk),
    .out(_U895_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U896 (
    .in(_U895_out),
    .clk(clk),
    .out(_U896_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U897 (
    .in(_U896_out),
    .clk(clk),
    .out(_U897_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U898 (
    .in(_U897_out),
    .clk(clk),
    .out(_U898_out)
);
_U899_pt__U900 _U899 (
    .in(_U901_out),
    .out(_U899_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U901 (
    .in(add_conv_stencil_5_999_1000_out),
    .clk(clk),
    .out(_U901_out)
);
_U902_pt__U903 _U902 (
    .in(_U904_out),
    .out(_U902_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U904 (
    .in(add_987_998_999_out),
    .clk(clk),
    .out(_U904_out)
);
_U905_pt__U906 _U905 (
    .in(_U913_out),
    .out(_U905_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U907 (
    .in(mul_hw_kernel_global_wrapper_stencil_36_hw_input_global_wrapper_stencil_36_989_out),
    .clk(clk),
    .out(_U907_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U908 (
    .in(_U907_out),
    .clk(clk),
    .out(_U908_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U909 (
    .in(_U908_out),
    .clk(clk),
    .out(_U909_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U910 (
    .in(_U909_out),
    .clk(clk),
    .out(_U910_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U911 (
    .in(_U910_out),
    .clk(clk),
    .out(_U911_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U912 (
    .in(_U911_out),
    .clk(clk),
    .out(_U912_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U913 (
    .in(_U912_out),
    .clk(clk),
    .out(_U913_out)
);
_U914_pt__U915 _U914 (
    .in(_U916_out),
    .out(_U914_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U916 (
    .in(add_988_997_998_out),
    .clk(clk),
    .out(_U916_out)
);
_U917_pt__U918 _U917 (
    .in(_U931_out),
    .out(_U917_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U919 (
    .in(mul_hw_kernel_global_wrapper_stencil_33_hw_input_global_wrapper_stencil_33_986_out),
    .clk(clk),
    .out(_U919_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U920 (
    .in(_U919_out),
    .clk(clk),
    .out(_U920_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U921 (
    .in(_U920_out),
    .clk(clk),
    .out(_U921_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U922 (
    .in(_U921_out),
    .clk(clk),
    .out(_U922_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U923 (
    .in(_U922_out),
    .clk(clk),
    .out(_U923_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U924 (
    .in(_U923_out),
    .clk(clk),
    .out(_U924_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U925 (
    .in(_U924_out),
    .clk(clk),
    .out(_U925_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U926 (
    .in(_U925_out),
    .clk(clk),
    .out(_U926_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U927 (
    .in(_U926_out),
    .clk(clk),
    .out(_U927_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U928 (
    .in(_U927_out),
    .clk(clk),
    .out(_U928_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U929 (
    .in(_U928_out),
    .clk(clk),
    .out(_U929_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U930 (
    .in(_U929_out),
    .clk(clk),
    .out(_U930_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U931 (
    .in(_U930_out),
    .clk(clk),
    .out(_U931_out)
);
_U932_pt__U933 _U932 (
    .in(_U937_out),
    .out(_U932_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U934 (
    .in(in1_hw_input_global_wrapper_stencil[3]),
    .clk(clk),
    .out(_U934_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U935 (
    .in(_U934_out),
    .clk(clk),
    .out(_U935_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U936 (
    .in(_U935_out),
    .clk(clk),
    .out(_U936_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U937 (
    .in(_U936_out),
    .clk(clk),
    .out(_U937_out)
);
_U938_pt__U939 _U938 (
    .in(_U945_out),
    .out(_U938_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U940 (
    .in(in2_hw_kernel_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U940_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U941 (
    .in(_U940_out),
    .clk(clk),
    .out(_U941_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U942 (
    .in(_U941_out),
    .clk(clk),
    .out(_U942_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U943 (
    .in(_U942_out),
    .clk(clk),
    .out(_U943_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U944 (
    .in(_U943_out),
    .clk(clk),
    .out(_U944_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U945 (
    .in(_U944_out),
    .clk(clk),
    .out(_U945_out)
);
_U946_pt__U947 _U946 (
    .in(_U948_out),
    .out(_U946_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U948 (
    .in(in1_hw_input_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U948_out)
);
_U949_pt__U950 _U949 (
    .in(_U956_out),
    .out(_U949_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U951 (
    .in(in1_hw_input_global_wrapper_stencil[2]),
    .clk(clk),
    .out(_U951_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U952 (
    .in(_U951_out),
    .clk(clk),
    .out(_U952_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U953 (
    .in(_U952_out),
    .clk(clk),
    .out(_U953_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U954 (
    .in(_U953_out),
    .clk(clk),
    .out(_U954_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U955 (
    .in(_U954_out),
    .clk(clk),
    .out(_U955_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U956 (
    .in(_U955_out),
    .clk(clk),
    .out(_U956_out)
);
_U957_pt__U958 _U957 (
    .in(_U960_out),
    .out(_U957_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U959 (
    .in(in2_hw_kernel_global_wrapper_stencil[0]),
    .clk(clk),
    .out(_U959_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U960 (
    .in(_U959_out),
    .clk(clk),
    .out(_U960_out)
);
_U961_pt__U962 _U961 (
    .in(_U964_out),
    .out(_U961_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U963 (
    .in(in1_hw_input_global_wrapper_stencil[0]),
    .clk(clk),
    .out(_U963_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U964 (
    .in(_U963_out),
    .clk(clk),
    .out(_U964_out)
);
_U965_pt__U966 _U965 (
    .in(_U972_out),
    .out(_U965_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U967 (
    .in(mul_hw_kernel_global_wrapper_stencil_35_hw_input_global_wrapper_stencil_35_988_out),
    .clk(clk),
    .out(_U967_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U968 (
    .in(_U967_out),
    .clk(clk),
    .out(_U968_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U969 (
    .in(_U968_out),
    .clk(clk),
    .out(_U969_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U970 (
    .in(_U969_out),
    .clk(clk),
    .out(_U970_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U971 (
    .in(_U970_out),
    .clk(clk),
    .out(_U971_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U972 (
    .in(_U971_out),
    .clk(clk),
    .out(_U972_out)
);
_U973_pt__U974 _U973 (
    .in(_U986_out),
    .out(_U973_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U975 (
    .in(mul_hw_kernel_global_wrapper_stencil_34_hw_input_global_wrapper_stencil_34_987_out),
    .clk(clk),
    .out(_U975_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U976 (
    .in(_U975_out),
    .clk(clk),
    .out(_U976_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U977 (
    .in(_U976_out),
    .clk(clk),
    .out(_U977_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U978 (
    .in(_U977_out),
    .clk(clk),
    .out(_U978_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U979 (
    .in(_U978_out),
    .clk(clk),
    .out(_U979_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U980 (
    .in(_U979_out),
    .clk(clk),
    .out(_U980_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U981 (
    .in(_U980_out),
    .clk(clk),
    .out(_U981_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U982 (
    .in(_U981_out),
    .clk(clk),
    .out(_U982_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U983 (
    .in(_U982_out),
    .clk(clk),
    .out(_U983_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U984 (
    .in(_U983_out),
    .clk(clk),
    .out(_U984_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U985 (
    .in(_U984_out),
    .clk(clk),
    .out(_U985_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U986 (
    .in(_U985_out),
    .clk(clk),
    .out(_U986_out)
);
_U987_pt__U988 _U987 (
    .in(_U989_out),
    .out(_U987_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U989 (
    .in(in2_hw_kernel_global_wrapper_stencil[1]),
    .clk(clk),
    .out(_U989_out)
);
_U990_pt__U991 _U990 (
    .in(_U996_out),
    .out(_U990_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U992 (
    .in(in2_hw_kernel_global_wrapper_stencil[7]),
    .clk(clk),
    .out(_U992_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U993 (
    .in(_U992_out),
    .clk(clk),
    .out(_U993_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U994 (
    .in(_U993_out),
    .clk(clk),
    .out(_U994_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U995 (
    .in(_U994_out),
    .clk(clk),
    .out(_U995_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U996 (
    .in(_U995_out),
    .clk(clk),
    .out(_U996_out)
);
_U997_pt__U998 _U997 (
    .in(_U1001_out),
    .out(_U997_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U999 (
    .in(in1_hw_input_global_wrapper_stencil[5]),
    .clk(clk),
    .out(_U999_out)
);
assign add_986_1000_1001_out = 16'(_U917_out + _U899_out);
assign add_987_998_999_out = 16'(_U973_out + _U914_out);
assign add_988_997_998_out = 16'(_U965_out + _U856_out);
assign add_989_996_997_out = 16'(_U905_out + _U888_out);
assign add_990_995_996_out = 16'(_U864_out + _U882_out);
assign add_991_994_995_out = 16'(_U891_out + _U885_out);
assign add_992_993_994_out = 16'(_U1002_out + _U859_out);
assign add_conv_stencil_5_999_1000_out = 16'(_U840_out + _U902_out);
assign mul_hw_kernel_global_wrapper_stencil_33_hw_input_global_wrapper_stencil_33_986_out = 16'(_U957_out * _U961_out);
assign mul_hw_kernel_global_wrapper_stencil_34_hw_input_global_wrapper_stencil_34_987_out = 16'(_U987_out * _U946_out);
assign mul_hw_kernel_global_wrapper_stencil_35_hw_input_global_wrapper_stencil_35_988_out = 16'(_U938_out * _U949_out);
assign mul_hw_kernel_global_wrapper_stencil_36_hw_input_global_wrapper_stencil_36_989_out = 16'(_U876_out * _U932_out);
assign mul_hw_kernel_global_wrapper_stencil_37_hw_input_global_wrapper_stencil_37_990_out = 16'(_U1010_out * _U1028_out);
assign mul_hw_kernel_global_wrapper_stencil_38_hw_input_global_wrapper_stencil_38_991_out = 16'(_U1005_out * _U997_out);
assign mul_hw_kernel_global_wrapper_stencil_39_hw_input_global_wrapper_stencil_39_992_out = 16'(_U1012_out * _U1030_out);
assign mul_hw_kernel_global_wrapper_stencil_40_hw_input_global_wrapper_stencil_40_993_out = 16'(_U990_out * _U1021_out);
endmodule

module cu_op_hcompute_conv_stencil_12 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_12_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_12_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_12_read[0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[0];
hcompute_conv_stencil_12_pipelined inner_compute (
    .clk(clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_12_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U0_pt__U1 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
_U0_pt__U1 _U0 (
    .in(in0_hw_input_stencil[0]),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read[0];
hcompute_hw_input_global_wrapper_stencil_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module resnet88 (
    input clk,
    input rst_n,
    input flush,
    output hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read_en,
    input [15:0] hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read_en,
    input [15:0] hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read [0:0],
    output hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read_en,
    input [15:0] hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read [0:0],
    output hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read_en,
    input [15:0] hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read [0:0],
    output hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read_en,
    input [15:0] hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read [0:0],
    output hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read_en,
    input [15:0] hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read [0:0],
    output hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read_en,
    input [15:0] hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read [0:0],
    output hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read_en,
    input [15:0] hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read [0:0],
    output hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write_valid,
    output [15:0] hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write [0:0],
    output hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write_valid,
    output [15:0] hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write [0:0],
    output hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write_valid,
    output [15:0] hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write [0:0],
    output hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write_valid,
    output [15:0] hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write [0:0],
    output hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write_valid,
    output [15:0] hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write [0:0],
    output hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write_valid,
    output [15:0] hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write [0:0],
    output hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write_valid,
    output [15:0] hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write [0:0],
    output hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write_valid,
    output [15:0] hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write [0:0]
);
wire [15:0] arr__U1004_out [4:0];
wire [15:0] arr__U1011_out [4:0];
wire [15:0] arr__U1037_out [4:0];
wire [15:0] arr__U1044_out [4:0];
wire [15:0] arr__U1051_out [4:0];
wire [15:0] arr__U1058_out [4:0];
wire [15:0] arr__U1065_out [4:0];
wire [15:0] arr__U1072_out [4:0];
wire [15:0] arr__U1079_out [4:0];
wire [15:0] arr__U1086_out [4:0];
wire [15:0] arr__U1093_out [4:0];
wire [15:0] arr__U1100_out [4:0];
wire [15:0] arr__U1107_out [4:0];
wire [15:0] arr__U1114_out [4:0];
wire [15:0] arr__U1121_out [4:0];
wire [15:0] arr__U1128_out [4:0];
wire [15:0] arr__U1135_out [4:0];
wire [15:0] arr__U1142_out [4:0];
wire [15:0] arr__U1149_out [4:0];
wire [15:0] arr__U1192_out [4:0];
wire [15:0] arr__U1199_out [4:0];
wire [15:0] arr__U1225_out [4:0];
wire [15:0] arr__U1232_out [4:0];
wire [15:0] arr__U1239_out [4:0];
wire [15:0] arr__U1246_out [4:0];
wire [15:0] arr__U1253_out [4:0];
wire [15:0] arr__U1260_out [4:0];
wire [15:0] arr__U1267_out [4:0];
wire [15:0] arr__U1274_out [4:0];
wire [15:0] arr__U1281_out [4:0];
wire [15:0] arr__U1288_out [4:0];
wire [15:0] arr__U1295_out [4:0];
wire [15:0] arr__U1302_out [4:0];
wire [15:0] arr__U1309_out [4:0];
wire [15:0] arr__U1316_out [4:0];
wire [15:0] arr__U1323_out [4:0];
wire [15:0] arr__U1330_out [4:0];
wire [15:0] arr__U1337_out [4:0];
wire [15:0] arr__U1380_out [4:0];
wire [15:0] arr__U1387_out [4:0];
wire [15:0] arr__U1413_out [4:0];
wire [15:0] arr__U1420_out [4:0];
wire [15:0] arr__U1427_out [4:0];
wire [15:0] arr__U1434_out [4:0];
wire [15:0] arr__U1441_out [4:0];
wire [15:0] arr__U1448_out [4:0];
wire [15:0] arr__U1455_out [4:0];
wire [15:0] arr__U1462_out [4:0];
wire [15:0] arr__U1469_out [4:0];
wire [15:0] arr__U1476_out [4:0];
wire [15:0] arr__U1483_out [4:0];
wire [15:0] arr__U1490_out [4:0];
wire [15:0] arr__U1497_out [4:0];
wire [15:0] arr__U1504_out [4:0];
wire [15:0] arr__U1511_out [4:0];
wire [15:0] arr__U1518_out [4:0];
wire [15:0] arr__U1525_out [4:0];
wire [15:0] arr__U1568_out [4:0];
wire [15:0] arr__U1575_out [4:0];
wire [15:0] arr__U1601_out [4:0];
wire [15:0] arr__U1608_out [4:0];
wire [15:0] arr__U1615_out [4:0];
wire [15:0] arr__U1622_out [4:0];
wire [15:0] arr__U1629_out [4:0];
wire [15:0] arr__U1636_out [4:0];
wire [15:0] arr__U1643_out [4:0];
wire [15:0] arr__U1650_out [4:0];
wire [15:0] arr__U1657_out [4:0];
wire [15:0] arr__U1664_out [4:0];
wire [15:0] arr__U1671_out [4:0];
wire [15:0] arr__U1678_out [4:0];
wire [15:0] arr__U1685_out [4:0];
wire [15:0] arr__U1692_out [4:0];
wire [15:0] arr__U1699_out [4:0];
wire [15:0] arr__U1706_out [4:0];
wire [15:0] arr__U1713_out [4:0];
wire [15:0] arr__U1756_out [4:0];
wire [15:0] arr__U1763_out [4:0];
wire [15:0] arr__U1789_out [4:0];
wire [15:0] arr__U1796_out [4:0];
wire [15:0] arr__U1803_out [4:0];
wire [15:0] arr__U1810_out [4:0];
wire [15:0] arr__U1817_out [4:0];
wire [15:0] arr__U1824_out [4:0];
wire [15:0] arr__U1831_out [4:0];
wire [15:0] arr__U1838_out [4:0];
wire [15:0] arr__U1845_out [4:0];
wire [15:0] arr__U1852_out [4:0];
wire [15:0] arr__U1859_out [4:0];
wire [15:0] arr__U1866_out [4:0];
wire [15:0] arr__U1873_out [4:0];
wire [15:0] arr__U1880_out [4:0];
wire [15:0] arr__U1887_out [4:0];
wire [15:0] arr__U1894_out [4:0];
wire [15:0] arr__U1901_out [4:0];
wire [15:0] arr__U1931_out [2:0];
wire [15:0] arr__U1936_out [2:0];
wire [15:0] arr__U1945_out [2:0];
wire [15:0] arr__U1950_out [2:0];
wire [15:0] arr__U1978_out [2:0];
wire [15:0] arr__U1983_out [2:0];
wire [15:0] arr__U1992_out [2:0];
wire [15:0] arr__U1997_out [2:0];
wire [15:0] arr__U2025_out [2:0];
wire [15:0] arr__U2030_out [2:0];
wire [15:0] arr__U2039_out [2:0];
wire [15:0] arr__U2044_out [2:0];
wire [15:0] arr__U2072_out [2:0];
wire [15:0] arr__U2077_out [2:0];
wire [15:0] arr__U2086_out [2:0];
wire [15:0] arr__U2091_out [2:0];
wire [15:0] arr__U2119_out [2:0];
wire [15:0] arr__U2124_out [2:0];
wire [15:0] arr__U2133_out [2:0];
wire [15:0] arr__U2138_out [2:0];
wire [15:0] arr__U2166_out [2:0];
wire [15:0] arr__U2171_out [2:0];
wire [15:0] arr__U2180_out [2:0];
wire [15:0] arr__U2185_out [2:0];
wire [15:0] arr__U2213_out [2:0];
wire [15:0] arr__U2218_out [2:0];
wire [15:0] arr__U2227_out [2:0];
wire [15:0] arr__U2232_out [2:0];
wire [15:0] arr__U2260_out [2:0];
wire [15:0] arr__U2265_out [2:0];
wire [15:0] arr__U2274_out [2:0];
wire [15:0] arr__U2279_out [2:0];
wire [15:0] arr__U440_out [4:0];
wire [15:0] arr__U447_out [4:0];
wire [15:0] arr__U473_out [4:0];
wire [15:0] arr__U480_out [4:0];
wire [15:0] arr__U487_out [4:0];
wire [15:0] arr__U494_out [4:0];
wire [15:0] arr__U501_out [4:0];
wire [15:0] arr__U508_out [4:0];
wire [15:0] arr__U515_out [4:0];
wire [15:0] arr__U522_out [4:0];
wire [15:0] arr__U529_out [4:0];
wire [15:0] arr__U536_out [4:0];
wire [15:0] arr__U543_out [4:0];
wire [15:0] arr__U550_out [4:0];
wire [15:0] arr__U557_out [4:0];
wire [15:0] arr__U564_out [4:0];
wire [15:0] arr__U571_out [4:0];
wire [15:0] arr__U578_out [4:0];
wire [15:0] arr__U585_out [4:0];
wire [15:0] arr__U628_out [4:0];
wire [15:0] arr__U635_out [4:0];
wire [15:0] arr__U661_out [4:0];
wire [15:0] arr__U668_out [4:0];
wire [15:0] arr__U675_out [4:0];
wire [15:0] arr__U682_out [4:0];
wire [15:0] arr__U689_out [4:0];
wire [15:0] arr__U696_out [4:0];
wire [15:0] arr__U703_out [4:0];
wire [15:0] arr__U710_out [4:0];
wire [15:0] arr__U717_out [4:0];
wire [15:0] arr__U724_out [4:0];
wire [15:0] arr__U731_out [4:0];
wire [15:0] arr__U738_out [4:0];
wire [15:0] arr__U745_out [4:0];
wire [15:0] arr__U752_out [4:0];
wire [15:0] arr__U759_out [4:0];
wire [15:0] arr__U766_out [4:0];
wire [15:0] arr__U773_out [4:0];
wire [15:0] arr__U816_out [4:0];
wire [15:0] arr__U823_out [4:0];
wire [15:0] arr__U849_out [4:0];
wire [15:0] arr__U856_out [4:0];
wire [15:0] arr__U863_out [4:0];
wire [15:0] arr__U870_out [4:0];
wire [15:0] arr__U877_out [4:0];
wire [15:0] arr__U884_out [4:0];
wire [15:0] arr__U891_out [4:0];
wire [15:0] arr__U898_out [4:0];
wire [15:0] arr__U905_out [4:0];
wire [15:0] arr__U912_out [4:0];
wire [15:0] arr__U919_out [4:0];
wire [15:0] arr__U926_out [4:0];
wire [15:0] arr__U933_out [4:0];
wire [15:0] arr__U940_out [4:0];
wire [15:0] arr__U947_out [4:0];
wire [15:0] arr__U954_out [4:0];
wire [15:0] arr__U961_out [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_10_read [0:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_11_read [0:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_12_read [0:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_13_read [0:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_14_read [0:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_15_read [0:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_8_read [0:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_9_read [0:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_1_read [0:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_2_read [0:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_3_read [0:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_4_read [0:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_5_read [0:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_6_read [0:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_7_read [0:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire delay_reg__U1001_out;
wire delay_reg__U1002_out;
wire delay_reg__U1019_out;
wire delay_reg__U1020_out;
wire delay_reg__U1021_out;
wire delay_reg__U1022_out;
wire delay_reg__U1023_out;
wire delay_reg__U1024_out;
wire delay_reg__U1025_out;
wire delay_reg__U1026_out;
wire delay_reg__U1027_out;
wire delay_reg__U1028_out;
wire delay_reg__U1029_out;
wire delay_reg__U1030_out;
wire delay_reg__U1031_out;
wire delay_reg__U1032_out;
wire delay_reg__U1033_out;
wire delay_reg__U1034_out;
wire delay_reg__U1035_out;
wire delay_reg__U1189_out;
wire delay_reg__U1190_out;
wire delay_reg__U1207_out;
wire delay_reg__U1208_out;
wire delay_reg__U1209_out;
wire delay_reg__U1210_out;
wire delay_reg__U1211_out;
wire delay_reg__U1212_out;
wire delay_reg__U1213_out;
wire delay_reg__U1214_out;
wire delay_reg__U1215_out;
wire delay_reg__U1216_out;
wire delay_reg__U1217_out;
wire delay_reg__U1218_out;
wire delay_reg__U1219_out;
wire delay_reg__U1220_out;
wire delay_reg__U1221_out;
wire delay_reg__U1222_out;
wire delay_reg__U1223_out;
wire delay_reg__U1377_out;
wire delay_reg__U1378_out;
wire delay_reg__U1395_out;
wire delay_reg__U1396_out;
wire delay_reg__U1397_out;
wire delay_reg__U1398_out;
wire delay_reg__U1399_out;
wire delay_reg__U1400_out;
wire delay_reg__U1401_out;
wire delay_reg__U1402_out;
wire delay_reg__U1403_out;
wire delay_reg__U1404_out;
wire delay_reg__U1405_out;
wire delay_reg__U1406_out;
wire delay_reg__U1407_out;
wire delay_reg__U1408_out;
wire delay_reg__U1409_out;
wire delay_reg__U1410_out;
wire delay_reg__U1411_out;
wire delay_reg__U1565_out;
wire delay_reg__U1566_out;
wire delay_reg__U1583_out;
wire delay_reg__U1584_out;
wire delay_reg__U1585_out;
wire delay_reg__U1586_out;
wire delay_reg__U1587_out;
wire delay_reg__U1588_out;
wire delay_reg__U1589_out;
wire delay_reg__U1590_out;
wire delay_reg__U1591_out;
wire delay_reg__U1592_out;
wire delay_reg__U1593_out;
wire delay_reg__U1594_out;
wire delay_reg__U1595_out;
wire delay_reg__U1596_out;
wire delay_reg__U1597_out;
wire delay_reg__U1598_out;
wire delay_reg__U1599_out;
wire delay_reg__U1753_out;
wire delay_reg__U1754_out;
wire delay_reg__U1771_out;
wire delay_reg__U1772_out;
wire delay_reg__U1773_out;
wire delay_reg__U1774_out;
wire delay_reg__U1775_out;
wire delay_reg__U1776_out;
wire delay_reg__U1777_out;
wire delay_reg__U1778_out;
wire delay_reg__U1779_out;
wire delay_reg__U1780_out;
wire delay_reg__U1781_out;
wire delay_reg__U1782_out;
wire delay_reg__U1783_out;
wire delay_reg__U1784_out;
wire delay_reg__U1785_out;
wire delay_reg__U1786_out;
wire delay_reg__U1787_out;
wire delay_reg__U1928_out;
wire delay_reg__U1929_out;
wire delay_reg__U1942_out;
wire delay_reg__U1943_out;
wire delay_reg__U1975_out;
wire delay_reg__U1976_out;
wire delay_reg__U1989_out;
wire delay_reg__U1990_out;
wire delay_reg__U2022_out;
wire delay_reg__U2023_out;
wire delay_reg__U2036_out;
wire delay_reg__U2037_out;
wire delay_reg__U2069_out;
wire delay_reg__U2070_out;
wire delay_reg__U2083_out;
wire delay_reg__U2084_out;
wire delay_reg__U2116_out;
wire delay_reg__U2117_out;
wire delay_reg__U2130_out;
wire delay_reg__U2131_out;
wire delay_reg__U2163_out;
wire delay_reg__U2164_out;
wire delay_reg__U2177_out;
wire delay_reg__U2178_out;
wire delay_reg__U2210_out;
wire delay_reg__U2211_out;
wire delay_reg__U2224_out;
wire delay_reg__U2225_out;
wire delay_reg__U2257_out;
wire delay_reg__U2258_out;
wire delay_reg__U2271_out;
wire delay_reg__U2272_out;
wire delay_reg__U437_out;
wire delay_reg__U438_out;
wire delay_reg__U455_out;
wire delay_reg__U456_out;
wire delay_reg__U457_out;
wire delay_reg__U458_out;
wire delay_reg__U459_out;
wire delay_reg__U460_out;
wire delay_reg__U461_out;
wire delay_reg__U462_out;
wire delay_reg__U463_out;
wire delay_reg__U464_out;
wire delay_reg__U465_out;
wire delay_reg__U466_out;
wire delay_reg__U467_out;
wire delay_reg__U468_out;
wire delay_reg__U469_out;
wire delay_reg__U470_out;
wire delay_reg__U471_out;
wire delay_reg__U625_out;
wire delay_reg__U626_out;
wire delay_reg__U643_out;
wire delay_reg__U644_out;
wire delay_reg__U645_out;
wire delay_reg__U646_out;
wire delay_reg__U647_out;
wire delay_reg__U648_out;
wire delay_reg__U649_out;
wire delay_reg__U650_out;
wire delay_reg__U651_out;
wire delay_reg__U652_out;
wire delay_reg__U653_out;
wire delay_reg__U654_out;
wire delay_reg__U655_out;
wire delay_reg__U656_out;
wire delay_reg__U657_out;
wire delay_reg__U658_out;
wire delay_reg__U659_out;
wire delay_reg__U813_out;
wire delay_reg__U814_out;
wire delay_reg__U831_out;
wire delay_reg__U832_out;
wire delay_reg__U833_out;
wire delay_reg__U834_out;
wire delay_reg__U835_out;
wire delay_reg__U836_out;
wire delay_reg__U837_out;
wire delay_reg__U838_out;
wire delay_reg__U839_out;
wire delay_reg__U840_out;
wire delay_reg__U841_out;
wire delay_reg__U842_out;
wire delay_reg__U843_out;
wire delay_reg__U844_out;
wire delay_reg__U845_out;
wire delay_reg__U846_out;
wire delay_reg__U847_out;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read [7:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read [7:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read [7:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read [7:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read [7:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read [7:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read [7:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read [7:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read [7:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read [7:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read [7:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read [7:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read [7:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read [7:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read [7:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read [7:0];
wire [15:0] op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire [15:0] op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire [15:0] op_hcompute_conv_stencil_10_conv_stencil_op_hcompute_conv_stencil_10_write [0:0];
wire op_hcompute_conv_stencil_10_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_10_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_10_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_10_port_controller_d [4:0];
wire op_hcompute_conv_stencil_10_read_start_out;
wire [15:0] op_hcompute_conv_stencil_10_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_10_write_start_out;
wire [15:0] op_hcompute_conv_stencil_10_write_start_control_vars_out [4:0];
wire [15:0] op_hcompute_conv_stencil_11_conv_stencil_op_hcompute_conv_stencil_11_write [0:0];
wire op_hcompute_conv_stencil_11_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_11_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_11_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_11_port_controller_d [4:0];
wire op_hcompute_conv_stencil_11_read_start_out;
wire [15:0] op_hcompute_conv_stencil_11_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_11_write_start_out;
wire [15:0] op_hcompute_conv_stencil_11_write_start_control_vars_out [4:0];
wire [15:0] op_hcompute_conv_stencil_12_conv_stencil_op_hcompute_conv_stencil_12_write [0:0];
wire op_hcompute_conv_stencil_12_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_12_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_12_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_12_port_controller_d [4:0];
wire op_hcompute_conv_stencil_12_read_start_out;
wire [15:0] op_hcompute_conv_stencil_12_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_12_write_start_out;
wire [15:0] op_hcompute_conv_stencil_12_write_start_control_vars_out [4:0];
wire [15:0] op_hcompute_conv_stencil_13_conv_stencil_op_hcompute_conv_stencil_13_write [0:0];
wire op_hcompute_conv_stencil_13_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_13_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_13_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_13_port_controller_d [4:0];
wire op_hcompute_conv_stencil_13_read_start_out;
wire [15:0] op_hcompute_conv_stencil_13_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_13_write_start_out;
wire [15:0] op_hcompute_conv_stencil_13_write_start_control_vars_out [4:0];
wire [15:0] op_hcompute_conv_stencil_14_conv_stencil_op_hcompute_conv_stencil_14_write [0:0];
wire op_hcompute_conv_stencil_14_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_14_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_14_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_14_port_controller_d [4:0];
wire op_hcompute_conv_stencil_14_read_start_out;
wire [15:0] op_hcompute_conv_stencil_14_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_14_write_start_out;
wire [15:0] op_hcompute_conv_stencil_14_write_start_control_vars_out [4:0];
wire [15:0] op_hcompute_conv_stencil_15_conv_stencil_op_hcompute_conv_stencil_15_write [0:0];
wire op_hcompute_conv_stencil_15_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_15_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_15_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_15_port_controller_d [4:0];
wire op_hcompute_conv_stencil_15_read_start_out;
wire [15:0] op_hcompute_conv_stencil_15_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_15_write_start_out;
wire [15:0] op_hcompute_conv_stencil_15_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_1_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_1_port_controller_d [2:0];
wire op_hcompute_conv_stencil_1_read_start_out;
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_write_start_out;
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire op_hcompute_conv_stencil_2_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_2_port_controller_d [2:0];
wire op_hcompute_conv_stencil_2_read_start_out;
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_write_start_out;
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire op_hcompute_conv_stencil_3_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_3_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_3_port_controller_d [2:0];
wire op_hcompute_conv_stencil_3_read_start_out;
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_3_write_start_out;
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire op_hcompute_conv_stencil_4_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_4_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_4_port_controller_d [2:0];
wire op_hcompute_conv_stencil_4_read_start_out;
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_4_write_start_out;
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire op_hcompute_conv_stencil_5_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_5_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_5_port_controller_d [2:0];
wire op_hcompute_conv_stencil_5_read_start_out;
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_5_write_start_out;
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_conv_stencil_6_conv_stencil_op_hcompute_conv_stencil_6_write [0:0];
wire op_hcompute_conv_stencil_6_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_6_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_6_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_6_port_controller_d [2:0];
wire op_hcompute_conv_stencil_6_read_start_out;
wire [15:0] op_hcompute_conv_stencil_6_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_6_write_start_out;
wire [15:0] op_hcompute_conv_stencil_6_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_conv_stencil_7_conv_stencil_op_hcompute_conv_stencil_7_write [0:0];
wire op_hcompute_conv_stencil_7_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_7_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_7_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_7_port_controller_d [2:0];
wire op_hcompute_conv_stencil_7_read_start_out;
wire [15:0] op_hcompute_conv_stencil_7_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_7_write_start_out;
wire [15:0] op_hcompute_conv_stencil_7_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_conv_stencil_8_conv_stencil_op_hcompute_conv_stencil_8_write [0:0];
wire op_hcompute_conv_stencil_8_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_8_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_8_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_8_port_controller_d [4:0];
wire op_hcompute_conv_stencil_8_read_start_out;
wire [15:0] op_hcompute_conv_stencil_8_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_8_write_start_out;
wire [15:0] op_hcompute_conv_stencil_8_write_start_control_vars_out [4:0];
wire [15:0] op_hcompute_conv_stencil_9_conv_stencil_op_hcompute_conv_stencil_9_write [0:0];
wire op_hcompute_conv_stencil_9_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_9_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_9_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_9_port_controller_d [4:0];
wire op_hcompute_conv_stencil_9_read_start_out;
wire [15:0] op_hcompute_conv_stencil_9_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_9_write_start_out;
wire [15:0] op_hcompute_conv_stencil_9_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_port_controller_d [2:0];
wire op_hcompute_conv_stencil_read_start_out;
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_write_start_out;
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_1_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_2_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_3_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_4_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_5_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_6_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_7_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_port_controller_d [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out [4:0];
wire [15:0] op_hcompute_hw_output_stencil_hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write [0:0];
wire [15:0] op_hcompute_hw_output_stencil_1_hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write [0:0];
wire op_hcompute_hw_output_stencil_1_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_1_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_1_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_1_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_1_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_1_read_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_output_stencil_1_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_output_stencil_2_hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write [0:0];
wire op_hcompute_hw_output_stencil_2_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_2_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_2_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_2_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_2_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_2_read_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_output_stencil_2_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_output_stencil_3_hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write [0:0];
wire op_hcompute_hw_output_stencil_3_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_3_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_3_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_3_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_3_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_3_read_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_output_stencil_3_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_output_stencil_4_hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write [0:0];
wire op_hcompute_hw_output_stencil_4_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_4_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_4_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_4_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_4_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_4_read_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_output_stencil_4_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_output_stencil_5_hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write [0:0];
wire op_hcompute_hw_output_stencil_5_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_5_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_5_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_5_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_5_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_5_read_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_output_stencil_5_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_output_stencil_6_hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write [0:0];
wire op_hcompute_hw_output_stencil_6_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_6_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_6_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_6_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_6_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_6_read_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_output_stencil_6_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_output_stencil_7_hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write [0:0];
wire op_hcompute_hw_output_stencil_7_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_7_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_7_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_7_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_7_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_7_read_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_output_stencil_7_write_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_out [2:0];
wire [15:0] arr__U1004_in [4:0];
assign arr__U1004_in[4] = op_hcompute_conv_stencil_11_port_controller_d[4];
assign arr__U1004_in[3] = op_hcompute_conv_stencil_11_port_controller_d[3];
assign arr__U1004_in[2] = op_hcompute_conv_stencil_11_port_controller_d[2];
assign arr__U1004_in[1] = op_hcompute_conv_stencil_11_port_controller_d[1];
assign arr__U1004_in[0] = op_hcompute_conv_stencil_11_port_controller_d[0];
array_delay_U1005 arr__U1004 (
    .clk(clk),
    .in(arr__U1004_in),
    .out(arr__U1004_out)
);
wire [15:0] arr__U1011_in [4:0];
assign arr__U1011_in[4] = arr__U1004_out[4];
assign arr__U1011_in[3] = arr__U1004_out[3];
assign arr__U1011_in[2] = arr__U1004_out[2];
assign arr__U1011_in[1] = arr__U1004_out[1];
assign arr__U1011_in[0] = arr__U1004_out[0];
array_delay_U1012 arr__U1011 (
    .clk(clk),
    .in(arr__U1011_in),
    .out(arr__U1011_out)
);
wire [15:0] arr__U1037_in [4:0];
assign arr__U1037_in[4] = op_hcompute_conv_stencil_11_port_controller_d[4];
assign arr__U1037_in[3] = op_hcompute_conv_stencil_11_port_controller_d[3];
assign arr__U1037_in[2] = op_hcompute_conv_stencil_11_port_controller_d[2];
assign arr__U1037_in[1] = op_hcompute_conv_stencil_11_port_controller_d[1];
assign arr__U1037_in[0] = op_hcompute_conv_stencil_11_port_controller_d[0];
array_delay_U1038 arr__U1037 (
    .clk(clk),
    .in(arr__U1037_in),
    .out(arr__U1037_out)
);
wire [15:0] arr__U1044_in [4:0];
assign arr__U1044_in[4] = arr__U1037_out[4];
assign arr__U1044_in[3] = arr__U1037_out[3];
assign arr__U1044_in[2] = arr__U1037_out[2];
assign arr__U1044_in[1] = arr__U1037_out[1];
assign arr__U1044_in[0] = arr__U1037_out[0];
array_delay_U1045 arr__U1044 (
    .clk(clk),
    .in(arr__U1044_in),
    .out(arr__U1044_out)
);
wire [15:0] arr__U1051_in [4:0];
assign arr__U1051_in[4] = arr__U1044_out[4];
assign arr__U1051_in[3] = arr__U1044_out[3];
assign arr__U1051_in[2] = arr__U1044_out[2];
assign arr__U1051_in[1] = arr__U1044_out[1];
assign arr__U1051_in[0] = arr__U1044_out[0];
array_delay_U1052 arr__U1051 (
    .clk(clk),
    .in(arr__U1051_in),
    .out(arr__U1051_out)
);
wire [15:0] arr__U1058_in [4:0];
assign arr__U1058_in[4] = arr__U1051_out[4];
assign arr__U1058_in[3] = arr__U1051_out[3];
assign arr__U1058_in[2] = arr__U1051_out[2];
assign arr__U1058_in[1] = arr__U1051_out[1];
assign arr__U1058_in[0] = arr__U1051_out[0];
array_delay_U1059 arr__U1058 (
    .clk(clk),
    .in(arr__U1058_in),
    .out(arr__U1058_out)
);
wire [15:0] arr__U1065_in [4:0];
assign arr__U1065_in[4] = arr__U1058_out[4];
assign arr__U1065_in[3] = arr__U1058_out[3];
assign arr__U1065_in[2] = arr__U1058_out[2];
assign arr__U1065_in[1] = arr__U1058_out[1];
assign arr__U1065_in[0] = arr__U1058_out[0];
array_delay_U1066 arr__U1065 (
    .clk(clk),
    .in(arr__U1065_in),
    .out(arr__U1065_out)
);
wire [15:0] arr__U1072_in [4:0];
assign arr__U1072_in[4] = arr__U1065_out[4];
assign arr__U1072_in[3] = arr__U1065_out[3];
assign arr__U1072_in[2] = arr__U1065_out[2];
assign arr__U1072_in[1] = arr__U1065_out[1];
assign arr__U1072_in[0] = arr__U1065_out[0];
array_delay_U1073 arr__U1072 (
    .clk(clk),
    .in(arr__U1072_in),
    .out(arr__U1072_out)
);
wire [15:0] arr__U1079_in [4:0];
assign arr__U1079_in[4] = arr__U1072_out[4];
assign arr__U1079_in[3] = arr__U1072_out[3];
assign arr__U1079_in[2] = arr__U1072_out[2];
assign arr__U1079_in[1] = arr__U1072_out[1];
assign arr__U1079_in[0] = arr__U1072_out[0];
array_delay_U1080 arr__U1079 (
    .clk(clk),
    .in(arr__U1079_in),
    .out(arr__U1079_out)
);
wire [15:0] arr__U1086_in [4:0];
assign arr__U1086_in[4] = arr__U1079_out[4];
assign arr__U1086_in[3] = arr__U1079_out[3];
assign arr__U1086_in[2] = arr__U1079_out[2];
assign arr__U1086_in[1] = arr__U1079_out[1];
assign arr__U1086_in[0] = arr__U1079_out[0];
array_delay_U1087 arr__U1086 (
    .clk(clk),
    .in(arr__U1086_in),
    .out(arr__U1086_out)
);
wire [15:0] arr__U1093_in [4:0];
assign arr__U1093_in[4] = arr__U1086_out[4];
assign arr__U1093_in[3] = arr__U1086_out[3];
assign arr__U1093_in[2] = arr__U1086_out[2];
assign arr__U1093_in[1] = arr__U1086_out[1];
assign arr__U1093_in[0] = arr__U1086_out[0];
array_delay_U1094 arr__U1093 (
    .clk(clk),
    .in(arr__U1093_in),
    .out(arr__U1093_out)
);
wire [15:0] arr__U1100_in [4:0];
assign arr__U1100_in[4] = arr__U1093_out[4];
assign arr__U1100_in[3] = arr__U1093_out[3];
assign arr__U1100_in[2] = arr__U1093_out[2];
assign arr__U1100_in[1] = arr__U1093_out[1];
assign arr__U1100_in[0] = arr__U1093_out[0];
array_delay_U1101 arr__U1100 (
    .clk(clk),
    .in(arr__U1100_in),
    .out(arr__U1100_out)
);
wire [15:0] arr__U1107_in [4:0];
assign arr__U1107_in[4] = arr__U1100_out[4];
assign arr__U1107_in[3] = arr__U1100_out[3];
assign arr__U1107_in[2] = arr__U1100_out[2];
assign arr__U1107_in[1] = arr__U1100_out[1];
assign arr__U1107_in[0] = arr__U1100_out[0];
array_delay_U1108 arr__U1107 (
    .clk(clk),
    .in(arr__U1107_in),
    .out(arr__U1107_out)
);
wire [15:0] arr__U1114_in [4:0];
assign arr__U1114_in[4] = arr__U1107_out[4];
assign arr__U1114_in[3] = arr__U1107_out[3];
assign arr__U1114_in[2] = arr__U1107_out[2];
assign arr__U1114_in[1] = arr__U1107_out[1];
assign arr__U1114_in[0] = arr__U1107_out[0];
array_delay_U1115 arr__U1114 (
    .clk(clk),
    .in(arr__U1114_in),
    .out(arr__U1114_out)
);
wire [15:0] arr__U1121_in [4:0];
assign arr__U1121_in[4] = arr__U1114_out[4];
assign arr__U1121_in[3] = arr__U1114_out[3];
assign arr__U1121_in[2] = arr__U1114_out[2];
assign arr__U1121_in[1] = arr__U1114_out[1];
assign arr__U1121_in[0] = arr__U1114_out[0];
array_delay_U1122 arr__U1121 (
    .clk(clk),
    .in(arr__U1121_in),
    .out(arr__U1121_out)
);
wire [15:0] arr__U1128_in [4:0];
assign arr__U1128_in[4] = arr__U1121_out[4];
assign arr__U1128_in[3] = arr__U1121_out[3];
assign arr__U1128_in[2] = arr__U1121_out[2];
assign arr__U1128_in[1] = arr__U1121_out[1];
assign arr__U1128_in[0] = arr__U1121_out[0];
array_delay_U1129 arr__U1128 (
    .clk(clk),
    .in(arr__U1128_in),
    .out(arr__U1128_out)
);
wire [15:0] arr__U1135_in [4:0];
assign arr__U1135_in[4] = arr__U1128_out[4];
assign arr__U1135_in[3] = arr__U1128_out[3];
assign arr__U1135_in[2] = arr__U1128_out[2];
assign arr__U1135_in[1] = arr__U1128_out[1];
assign arr__U1135_in[0] = arr__U1128_out[0];
array_delay_U1136 arr__U1135 (
    .clk(clk),
    .in(arr__U1135_in),
    .out(arr__U1135_out)
);
wire [15:0] arr__U1142_in [4:0];
assign arr__U1142_in[4] = arr__U1135_out[4];
assign arr__U1142_in[3] = arr__U1135_out[3];
assign arr__U1142_in[2] = arr__U1135_out[2];
assign arr__U1142_in[1] = arr__U1135_out[1];
assign arr__U1142_in[0] = arr__U1135_out[0];
array_delay_U1143 arr__U1142 (
    .clk(clk),
    .in(arr__U1142_in),
    .out(arr__U1142_out)
);
wire [15:0] arr__U1149_in [4:0];
assign arr__U1149_in[4] = arr__U1142_out[4];
assign arr__U1149_in[3] = arr__U1142_out[3];
assign arr__U1149_in[2] = arr__U1142_out[2];
assign arr__U1149_in[1] = arr__U1142_out[1];
assign arr__U1149_in[0] = arr__U1142_out[0];
array_delay_U1150 arr__U1149 (
    .clk(clk),
    .in(arr__U1149_in),
    .out(arr__U1149_out)
);
wire [15:0] arr__U1192_in [4:0];
assign arr__U1192_in[4] = op_hcompute_conv_stencil_12_port_controller_d[4];
assign arr__U1192_in[3] = op_hcompute_conv_stencil_12_port_controller_d[3];
assign arr__U1192_in[2] = op_hcompute_conv_stencil_12_port_controller_d[2];
assign arr__U1192_in[1] = op_hcompute_conv_stencil_12_port_controller_d[1];
assign arr__U1192_in[0] = op_hcompute_conv_stencil_12_port_controller_d[0];
array_delay_U1193 arr__U1192 (
    .clk(clk),
    .in(arr__U1192_in),
    .out(arr__U1192_out)
);
wire [15:0] arr__U1199_in [4:0];
assign arr__U1199_in[4] = arr__U1192_out[4];
assign arr__U1199_in[3] = arr__U1192_out[3];
assign arr__U1199_in[2] = arr__U1192_out[2];
assign arr__U1199_in[1] = arr__U1192_out[1];
assign arr__U1199_in[0] = arr__U1192_out[0];
array_delay_U1200 arr__U1199 (
    .clk(clk),
    .in(arr__U1199_in),
    .out(arr__U1199_out)
);
wire [15:0] arr__U1225_in [4:0];
assign arr__U1225_in[4] = op_hcompute_conv_stencil_12_port_controller_d[4];
assign arr__U1225_in[3] = op_hcompute_conv_stencil_12_port_controller_d[3];
assign arr__U1225_in[2] = op_hcompute_conv_stencil_12_port_controller_d[2];
assign arr__U1225_in[1] = op_hcompute_conv_stencil_12_port_controller_d[1];
assign arr__U1225_in[0] = op_hcompute_conv_stencil_12_port_controller_d[0];
array_delay_U1226 arr__U1225 (
    .clk(clk),
    .in(arr__U1225_in),
    .out(arr__U1225_out)
);
wire [15:0] arr__U1232_in [4:0];
assign arr__U1232_in[4] = arr__U1225_out[4];
assign arr__U1232_in[3] = arr__U1225_out[3];
assign arr__U1232_in[2] = arr__U1225_out[2];
assign arr__U1232_in[1] = arr__U1225_out[1];
assign arr__U1232_in[0] = arr__U1225_out[0];
array_delay_U1233 arr__U1232 (
    .clk(clk),
    .in(arr__U1232_in),
    .out(arr__U1232_out)
);
wire [15:0] arr__U1239_in [4:0];
assign arr__U1239_in[4] = arr__U1232_out[4];
assign arr__U1239_in[3] = arr__U1232_out[3];
assign arr__U1239_in[2] = arr__U1232_out[2];
assign arr__U1239_in[1] = arr__U1232_out[1];
assign arr__U1239_in[0] = arr__U1232_out[0];
array_delay_U1240 arr__U1239 (
    .clk(clk),
    .in(arr__U1239_in),
    .out(arr__U1239_out)
);
wire [15:0] arr__U1246_in [4:0];
assign arr__U1246_in[4] = arr__U1239_out[4];
assign arr__U1246_in[3] = arr__U1239_out[3];
assign arr__U1246_in[2] = arr__U1239_out[2];
assign arr__U1246_in[1] = arr__U1239_out[1];
assign arr__U1246_in[0] = arr__U1239_out[0];
array_delay_U1247 arr__U1246 (
    .clk(clk),
    .in(arr__U1246_in),
    .out(arr__U1246_out)
);
wire [15:0] arr__U1253_in [4:0];
assign arr__U1253_in[4] = arr__U1246_out[4];
assign arr__U1253_in[3] = arr__U1246_out[3];
assign arr__U1253_in[2] = arr__U1246_out[2];
assign arr__U1253_in[1] = arr__U1246_out[1];
assign arr__U1253_in[0] = arr__U1246_out[0];
array_delay_U1254 arr__U1253 (
    .clk(clk),
    .in(arr__U1253_in),
    .out(arr__U1253_out)
);
wire [15:0] arr__U1260_in [4:0];
assign arr__U1260_in[4] = arr__U1253_out[4];
assign arr__U1260_in[3] = arr__U1253_out[3];
assign arr__U1260_in[2] = arr__U1253_out[2];
assign arr__U1260_in[1] = arr__U1253_out[1];
assign arr__U1260_in[0] = arr__U1253_out[0];
array_delay_U1261 arr__U1260 (
    .clk(clk),
    .in(arr__U1260_in),
    .out(arr__U1260_out)
);
wire [15:0] arr__U1267_in [4:0];
assign arr__U1267_in[4] = arr__U1260_out[4];
assign arr__U1267_in[3] = arr__U1260_out[3];
assign arr__U1267_in[2] = arr__U1260_out[2];
assign arr__U1267_in[1] = arr__U1260_out[1];
assign arr__U1267_in[0] = arr__U1260_out[0];
array_delay_U1268 arr__U1267 (
    .clk(clk),
    .in(arr__U1267_in),
    .out(arr__U1267_out)
);
wire [15:0] arr__U1274_in [4:0];
assign arr__U1274_in[4] = arr__U1267_out[4];
assign arr__U1274_in[3] = arr__U1267_out[3];
assign arr__U1274_in[2] = arr__U1267_out[2];
assign arr__U1274_in[1] = arr__U1267_out[1];
assign arr__U1274_in[0] = arr__U1267_out[0];
array_delay_U1275 arr__U1274 (
    .clk(clk),
    .in(arr__U1274_in),
    .out(arr__U1274_out)
);
wire [15:0] arr__U1281_in [4:0];
assign arr__U1281_in[4] = arr__U1274_out[4];
assign arr__U1281_in[3] = arr__U1274_out[3];
assign arr__U1281_in[2] = arr__U1274_out[2];
assign arr__U1281_in[1] = arr__U1274_out[1];
assign arr__U1281_in[0] = arr__U1274_out[0];
array_delay_U1282 arr__U1281 (
    .clk(clk),
    .in(arr__U1281_in),
    .out(arr__U1281_out)
);
wire [15:0] arr__U1288_in [4:0];
assign arr__U1288_in[4] = arr__U1281_out[4];
assign arr__U1288_in[3] = arr__U1281_out[3];
assign arr__U1288_in[2] = arr__U1281_out[2];
assign arr__U1288_in[1] = arr__U1281_out[1];
assign arr__U1288_in[0] = arr__U1281_out[0];
array_delay_U1289 arr__U1288 (
    .clk(clk),
    .in(arr__U1288_in),
    .out(arr__U1288_out)
);
wire [15:0] arr__U1295_in [4:0];
assign arr__U1295_in[4] = arr__U1288_out[4];
assign arr__U1295_in[3] = arr__U1288_out[3];
assign arr__U1295_in[2] = arr__U1288_out[2];
assign arr__U1295_in[1] = arr__U1288_out[1];
assign arr__U1295_in[0] = arr__U1288_out[0];
array_delay_U1296 arr__U1295 (
    .clk(clk),
    .in(arr__U1295_in),
    .out(arr__U1295_out)
);
wire [15:0] arr__U1302_in [4:0];
assign arr__U1302_in[4] = arr__U1295_out[4];
assign arr__U1302_in[3] = arr__U1295_out[3];
assign arr__U1302_in[2] = arr__U1295_out[2];
assign arr__U1302_in[1] = arr__U1295_out[1];
assign arr__U1302_in[0] = arr__U1295_out[0];
array_delay_U1303 arr__U1302 (
    .clk(clk),
    .in(arr__U1302_in),
    .out(arr__U1302_out)
);
wire [15:0] arr__U1309_in [4:0];
assign arr__U1309_in[4] = arr__U1302_out[4];
assign arr__U1309_in[3] = arr__U1302_out[3];
assign arr__U1309_in[2] = arr__U1302_out[2];
assign arr__U1309_in[1] = arr__U1302_out[1];
assign arr__U1309_in[0] = arr__U1302_out[0];
array_delay_U1310 arr__U1309 (
    .clk(clk),
    .in(arr__U1309_in),
    .out(arr__U1309_out)
);
wire [15:0] arr__U1316_in [4:0];
assign arr__U1316_in[4] = arr__U1309_out[4];
assign arr__U1316_in[3] = arr__U1309_out[3];
assign arr__U1316_in[2] = arr__U1309_out[2];
assign arr__U1316_in[1] = arr__U1309_out[1];
assign arr__U1316_in[0] = arr__U1309_out[0];
array_delay_U1317 arr__U1316 (
    .clk(clk),
    .in(arr__U1316_in),
    .out(arr__U1316_out)
);
wire [15:0] arr__U1323_in [4:0];
assign arr__U1323_in[4] = arr__U1316_out[4];
assign arr__U1323_in[3] = arr__U1316_out[3];
assign arr__U1323_in[2] = arr__U1316_out[2];
assign arr__U1323_in[1] = arr__U1316_out[1];
assign arr__U1323_in[0] = arr__U1316_out[0];
array_delay_U1324 arr__U1323 (
    .clk(clk),
    .in(arr__U1323_in),
    .out(arr__U1323_out)
);
wire [15:0] arr__U1330_in [4:0];
assign arr__U1330_in[4] = arr__U1323_out[4];
assign arr__U1330_in[3] = arr__U1323_out[3];
assign arr__U1330_in[2] = arr__U1323_out[2];
assign arr__U1330_in[1] = arr__U1323_out[1];
assign arr__U1330_in[0] = arr__U1323_out[0];
array_delay_U1331 arr__U1330 (
    .clk(clk),
    .in(arr__U1330_in),
    .out(arr__U1330_out)
);
wire [15:0] arr__U1337_in [4:0];
assign arr__U1337_in[4] = arr__U1330_out[4];
assign arr__U1337_in[3] = arr__U1330_out[3];
assign arr__U1337_in[2] = arr__U1330_out[2];
assign arr__U1337_in[1] = arr__U1330_out[1];
assign arr__U1337_in[0] = arr__U1330_out[0];
array_delay_U1338 arr__U1337 (
    .clk(clk),
    .in(arr__U1337_in),
    .out(arr__U1337_out)
);
wire [15:0] arr__U1380_in [4:0];
assign arr__U1380_in[4] = op_hcompute_conv_stencil_13_port_controller_d[4];
assign arr__U1380_in[3] = op_hcompute_conv_stencil_13_port_controller_d[3];
assign arr__U1380_in[2] = op_hcompute_conv_stencil_13_port_controller_d[2];
assign arr__U1380_in[1] = op_hcompute_conv_stencil_13_port_controller_d[1];
assign arr__U1380_in[0] = op_hcompute_conv_stencil_13_port_controller_d[0];
array_delay_U1381 arr__U1380 (
    .clk(clk),
    .in(arr__U1380_in),
    .out(arr__U1380_out)
);
wire [15:0] arr__U1387_in [4:0];
assign arr__U1387_in[4] = arr__U1380_out[4];
assign arr__U1387_in[3] = arr__U1380_out[3];
assign arr__U1387_in[2] = arr__U1380_out[2];
assign arr__U1387_in[1] = arr__U1380_out[1];
assign arr__U1387_in[0] = arr__U1380_out[0];
array_delay_U1388 arr__U1387 (
    .clk(clk),
    .in(arr__U1387_in),
    .out(arr__U1387_out)
);
wire [15:0] arr__U1413_in [4:0];
assign arr__U1413_in[4] = op_hcompute_conv_stencil_13_port_controller_d[4];
assign arr__U1413_in[3] = op_hcompute_conv_stencil_13_port_controller_d[3];
assign arr__U1413_in[2] = op_hcompute_conv_stencil_13_port_controller_d[2];
assign arr__U1413_in[1] = op_hcompute_conv_stencil_13_port_controller_d[1];
assign arr__U1413_in[0] = op_hcompute_conv_stencil_13_port_controller_d[0];
array_delay_U1414 arr__U1413 (
    .clk(clk),
    .in(arr__U1413_in),
    .out(arr__U1413_out)
);
wire [15:0] arr__U1420_in [4:0];
assign arr__U1420_in[4] = arr__U1413_out[4];
assign arr__U1420_in[3] = arr__U1413_out[3];
assign arr__U1420_in[2] = arr__U1413_out[2];
assign arr__U1420_in[1] = arr__U1413_out[1];
assign arr__U1420_in[0] = arr__U1413_out[0];
array_delay_U1421 arr__U1420 (
    .clk(clk),
    .in(arr__U1420_in),
    .out(arr__U1420_out)
);
wire [15:0] arr__U1427_in [4:0];
assign arr__U1427_in[4] = arr__U1420_out[4];
assign arr__U1427_in[3] = arr__U1420_out[3];
assign arr__U1427_in[2] = arr__U1420_out[2];
assign arr__U1427_in[1] = arr__U1420_out[1];
assign arr__U1427_in[0] = arr__U1420_out[0];
array_delay_U1428 arr__U1427 (
    .clk(clk),
    .in(arr__U1427_in),
    .out(arr__U1427_out)
);
wire [15:0] arr__U1434_in [4:0];
assign arr__U1434_in[4] = arr__U1427_out[4];
assign arr__U1434_in[3] = arr__U1427_out[3];
assign arr__U1434_in[2] = arr__U1427_out[2];
assign arr__U1434_in[1] = arr__U1427_out[1];
assign arr__U1434_in[0] = arr__U1427_out[0];
array_delay_U1435 arr__U1434 (
    .clk(clk),
    .in(arr__U1434_in),
    .out(arr__U1434_out)
);
wire [15:0] arr__U1441_in [4:0];
assign arr__U1441_in[4] = arr__U1434_out[4];
assign arr__U1441_in[3] = arr__U1434_out[3];
assign arr__U1441_in[2] = arr__U1434_out[2];
assign arr__U1441_in[1] = arr__U1434_out[1];
assign arr__U1441_in[0] = arr__U1434_out[0];
array_delay_U1442 arr__U1441 (
    .clk(clk),
    .in(arr__U1441_in),
    .out(arr__U1441_out)
);
wire [15:0] arr__U1448_in [4:0];
assign arr__U1448_in[4] = arr__U1441_out[4];
assign arr__U1448_in[3] = arr__U1441_out[3];
assign arr__U1448_in[2] = arr__U1441_out[2];
assign arr__U1448_in[1] = arr__U1441_out[1];
assign arr__U1448_in[0] = arr__U1441_out[0];
array_delay_U1449 arr__U1448 (
    .clk(clk),
    .in(arr__U1448_in),
    .out(arr__U1448_out)
);
wire [15:0] arr__U1455_in [4:0];
assign arr__U1455_in[4] = arr__U1448_out[4];
assign arr__U1455_in[3] = arr__U1448_out[3];
assign arr__U1455_in[2] = arr__U1448_out[2];
assign arr__U1455_in[1] = arr__U1448_out[1];
assign arr__U1455_in[0] = arr__U1448_out[0];
array_delay_U1456 arr__U1455 (
    .clk(clk),
    .in(arr__U1455_in),
    .out(arr__U1455_out)
);
wire [15:0] arr__U1462_in [4:0];
assign arr__U1462_in[4] = arr__U1455_out[4];
assign arr__U1462_in[3] = arr__U1455_out[3];
assign arr__U1462_in[2] = arr__U1455_out[2];
assign arr__U1462_in[1] = arr__U1455_out[1];
assign arr__U1462_in[0] = arr__U1455_out[0];
array_delay_U1463 arr__U1462 (
    .clk(clk),
    .in(arr__U1462_in),
    .out(arr__U1462_out)
);
wire [15:0] arr__U1469_in [4:0];
assign arr__U1469_in[4] = arr__U1462_out[4];
assign arr__U1469_in[3] = arr__U1462_out[3];
assign arr__U1469_in[2] = arr__U1462_out[2];
assign arr__U1469_in[1] = arr__U1462_out[1];
assign arr__U1469_in[0] = arr__U1462_out[0];
array_delay_U1470 arr__U1469 (
    .clk(clk),
    .in(arr__U1469_in),
    .out(arr__U1469_out)
);
wire [15:0] arr__U1476_in [4:0];
assign arr__U1476_in[4] = arr__U1469_out[4];
assign arr__U1476_in[3] = arr__U1469_out[3];
assign arr__U1476_in[2] = arr__U1469_out[2];
assign arr__U1476_in[1] = arr__U1469_out[1];
assign arr__U1476_in[0] = arr__U1469_out[0];
array_delay_U1477 arr__U1476 (
    .clk(clk),
    .in(arr__U1476_in),
    .out(arr__U1476_out)
);
wire [15:0] arr__U1483_in [4:0];
assign arr__U1483_in[4] = arr__U1476_out[4];
assign arr__U1483_in[3] = arr__U1476_out[3];
assign arr__U1483_in[2] = arr__U1476_out[2];
assign arr__U1483_in[1] = arr__U1476_out[1];
assign arr__U1483_in[0] = arr__U1476_out[0];
array_delay_U1484 arr__U1483 (
    .clk(clk),
    .in(arr__U1483_in),
    .out(arr__U1483_out)
);
wire [15:0] arr__U1490_in [4:0];
assign arr__U1490_in[4] = arr__U1483_out[4];
assign arr__U1490_in[3] = arr__U1483_out[3];
assign arr__U1490_in[2] = arr__U1483_out[2];
assign arr__U1490_in[1] = arr__U1483_out[1];
assign arr__U1490_in[0] = arr__U1483_out[0];
array_delay_U1491 arr__U1490 (
    .clk(clk),
    .in(arr__U1490_in),
    .out(arr__U1490_out)
);
wire [15:0] arr__U1497_in [4:0];
assign arr__U1497_in[4] = arr__U1490_out[4];
assign arr__U1497_in[3] = arr__U1490_out[3];
assign arr__U1497_in[2] = arr__U1490_out[2];
assign arr__U1497_in[1] = arr__U1490_out[1];
assign arr__U1497_in[0] = arr__U1490_out[0];
array_delay_U1498 arr__U1497 (
    .clk(clk),
    .in(arr__U1497_in),
    .out(arr__U1497_out)
);
wire [15:0] arr__U1504_in [4:0];
assign arr__U1504_in[4] = arr__U1497_out[4];
assign arr__U1504_in[3] = arr__U1497_out[3];
assign arr__U1504_in[2] = arr__U1497_out[2];
assign arr__U1504_in[1] = arr__U1497_out[1];
assign arr__U1504_in[0] = arr__U1497_out[0];
array_delay_U1505 arr__U1504 (
    .clk(clk),
    .in(arr__U1504_in),
    .out(arr__U1504_out)
);
wire [15:0] arr__U1511_in [4:0];
assign arr__U1511_in[4] = arr__U1504_out[4];
assign arr__U1511_in[3] = arr__U1504_out[3];
assign arr__U1511_in[2] = arr__U1504_out[2];
assign arr__U1511_in[1] = arr__U1504_out[1];
assign arr__U1511_in[0] = arr__U1504_out[0];
array_delay_U1512 arr__U1511 (
    .clk(clk),
    .in(arr__U1511_in),
    .out(arr__U1511_out)
);
wire [15:0] arr__U1518_in [4:0];
assign arr__U1518_in[4] = arr__U1511_out[4];
assign arr__U1518_in[3] = arr__U1511_out[3];
assign arr__U1518_in[2] = arr__U1511_out[2];
assign arr__U1518_in[1] = arr__U1511_out[1];
assign arr__U1518_in[0] = arr__U1511_out[0];
array_delay_U1519 arr__U1518 (
    .clk(clk),
    .in(arr__U1518_in),
    .out(arr__U1518_out)
);
wire [15:0] arr__U1525_in [4:0];
assign arr__U1525_in[4] = arr__U1518_out[4];
assign arr__U1525_in[3] = arr__U1518_out[3];
assign arr__U1525_in[2] = arr__U1518_out[2];
assign arr__U1525_in[1] = arr__U1518_out[1];
assign arr__U1525_in[0] = arr__U1518_out[0];
array_delay_U1526 arr__U1525 (
    .clk(clk),
    .in(arr__U1525_in),
    .out(arr__U1525_out)
);
wire [15:0] arr__U1568_in [4:0];
assign arr__U1568_in[4] = op_hcompute_conv_stencil_14_port_controller_d[4];
assign arr__U1568_in[3] = op_hcompute_conv_stencil_14_port_controller_d[3];
assign arr__U1568_in[2] = op_hcompute_conv_stencil_14_port_controller_d[2];
assign arr__U1568_in[1] = op_hcompute_conv_stencil_14_port_controller_d[1];
assign arr__U1568_in[0] = op_hcompute_conv_stencil_14_port_controller_d[0];
array_delay_U1569 arr__U1568 (
    .clk(clk),
    .in(arr__U1568_in),
    .out(arr__U1568_out)
);
wire [15:0] arr__U1575_in [4:0];
assign arr__U1575_in[4] = arr__U1568_out[4];
assign arr__U1575_in[3] = arr__U1568_out[3];
assign arr__U1575_in[2] = arr__U1568_out[2];
assign arr__U1575_in[1] = arr__U1568_out[1];
assign arr__U1575_in[0] = arr__U1568_out[0];
array_delay_U1576 arr__U1575 (
    .clk(clk),
    .in(arr__U1575_in),
    .out(arr__U1575_out)
);
wire [15:0] arr__U1601_in [4:0];
assign arr__U1601_in[4] = op_hcompute_conv_stencil_14_port_controller_d[4];
assign arr__U1601_in[3] = op_hcompute_conv_stencil_14_port_controller_d[3];
assign arr__U1601_in[2] = op_hcompute_conv_stencil_14_port_controller_d[2];
assign arr__U1601_in[1] = op_hcompute_conv_stencil_14_port_controller_d[1];
assign arr__U1601_in[0] = op_hcompute_conv_stencil_14_port_controller_d[0];
array_delay_U1602 arr__U1601 (
    .clk(clk),
    .in(arr__U1601_in),
    .out(arr__U1601_out)
);
wire [15:0] arr__U1608_in [4:0];
assign arr__U1608_in[4] = arr__U1601_out[4];
assign arr__U1608_in[3] = arr__U1601_out[3];
assign arr__U1608_in[2] = arr__U1601_out[2];
assign arr__U1608_in[1] = arr__U1601_out[1];
assign arr__U1608_in[0] = arr__U1601_out[0];
array_delay_U1609 arr__U1608 (
    .clk(clk),
    .in(arr__U1608_in),
    .out(arr__U1608_out)
);
wire [15:0] arr__U1615_in [4:0];
assign arr__U1615_in[4] = arr__U1608_out[4];
assign arr__U1615_in[3] = arr__U1608_out[3];
assign arr__U1615_in[2] = arr__U1608_out[2];
assign arr__U1615_in[1] = arr__U1608_out[1];
assign arr__U1615_in[0] = arr__U1608_out[0];
array_delay_U1616 arr__U1615 (
    .clk(clk),
    .in(arr__U1615_in),
    .out(arr__U1615_out)
);
wire [15:0] arr__U1622_in [4:0];
assign arr__U1622_in[4] = arr__U1615_out[4];
assign arr__U1622_in[3] = arr__U1615_out[3];
assign arr__U1622_in[2] = arr__U1615_out[2];
assign arr__U1622_in[1] = arr__U1615_out[1];
assign arr__U1622_in[0] = arr__U1615_out[0];
array_delay_U1623 arr__U1622 (
    .clk(clk),
    .in(arr__U1622_in),
    .out(arr__U1622_out)
);
wire [15:0] arr__U1629_in [4:0];
assign arr__U1629_in[4] = arr__U1622_out[4];
assign arr__U1629_in[3] = arr__U1622_out[3];
assign arr__U1629_in[2] = arr__U1622_out[2];
assign arr__U1629_in[1] = arr__U1622_out[1];
assign arr__U1629_in[0] = arr__U1622_out[0];
array_delay_U1630 arr__U1629 (
    .clk(clk),
    .in(arr__U1629_in),
    .out(arr__U1629_out)
);
wire [15:0] arr__U1636_in [4:0];
assign arr__U1636_in[4] = arr__U1629_out[4];
assign arr__U1636_in[3] = arr__U1629_out[3];
assign arr__U1636_in[2] = arr__U1629_out[2];
assign arr__U1636_in[1] = arr__U1629_out[1];
assign arr__U1636_in[0] = arr__U1629_out[0];
array_delay_U1637 arr__U1636 (
    .clk(clk),
    .in(arr__U1636_in),
    .out(arr__U1636_out)
);
wire [15:0] arr__U1643_in [4:0];
assign arr__U1643_in[4] = arr__U1636_out[4];
assign arr__U1643_in[3] = arr__U1636_out[3];
assign arr__U1643_in[2] = arr__U1636_out[2];
assign arr__U1643_in[1] = arr__U1636_out[1];
assign arr__U1643_in[0] = arr__U1636_out[0];
array_delay_U1644 arr__U1643 (
    .clk(clk),
    .in(arr__U1643_in),
    .out(arr__U1643_out)
);
wire [15:0] arr__U1650_in [4:0];
assign arr__U1650_in[4] = arr__U1643_out[4];
assign arr__U1650_in[3] = arr__U1643_out[3];
assign arr__U1650_in[2] = arr__U1643_out[2];
assign arr__U1650_in[1] = arr__U1643_out[1];
assign arr__U1650_in[0] = arr__U1643_out[0];
array_delay_U1651 arr__U1650 (
    .clk(clk),
    .in(arr__U1650_in),
    .out(arr__U1650_out)
);
wire [15:0] arr__U1657_in [4:0];
assign arr__U1657_in[4] = arr__U1650_out[4];
assign arr__U1657_in[3] = arr__U1650_out[3];
assign arr__U1657_in[2] = arr__U1650_out[2];
assign arr__U1657_in[1] = arr__U1650_out[1];
assign arr__U1657_in[0] = arr__U1650_out[0];
array_delay_U1658 arr__U1657 (
    .clk(clk),
    .in(arr__U1657_in),
    .out(arr__U1657_out)
);
wire [15:0] arr__U1664_in [4:0];
assign arr__U1664_in[4] = arr__U1657_out[4];
assign arr__U1664_in[3] = arr__U1657_out[3];
assign arr__U1664_in[2] = arr__U1657_out[2];
assign arr__U1664_in[1] = arr__U1657_out[1];
assign arr__U1664_in[0] = arr__U1657_out[0];
array_delay_U1665 arr__U1664 (
    .clk(clk),
    .in(arr__U1664_in),
    .out(arr__U1664_out)
);
wire [15:0] arr__U1671_in [4:0];
assign arr__U1671_in[4] = arr__U1664_out[4];
assign arr__U1671_in[3] = arr__U1664_out[3];
assign arr__U1671_in[2] = arr__U1664_out[2];
assign arr__U1671_in[1] = arr__U1664_out[1];
assign arr__U1671_in[0] = arr__U1664_out[0];
array_delay_U1672 arr__U1671 (
    .clk(clk),
    .in(arr__U1671_in),
    .out(arr__U1671_out)
);
wire [15:0] arr__U1678_in [4:0];
assign arr__U1678_in[4] = arr__U1671_out[4];
assign arr__U1678_in[3] = arr__U1671_out[3];
assign arr__U1678_in[2] = arr__U1671_out[2];
assign arr__U1678_in[1] = arr__U1671_out[1];
assign arr__U1678_in[0] = arr__U1671_out[0];
array_delay_U1679 arr__U1678 (
    .clk(clk),
    .in(arr__U1678_in),
    .out(arr__U1678_out)
);
wire [15:0] arr__U1685_in [4:0];
assign arr__U1685_in[4] = arr__U1678_out[4];
assign arr__U1685_in[3] = arr__U1678_out[3];
assign arr__U1685_in[2] = arr__U1678_out[2];
assign arr__U1685_in[1] = arr__U1678_out[1];
assign arr__U1685_in[0] = arr__U1678_out[0];
array_delay_U1686 arr__U1685 (
    .clk(clk),
    .in(arr__U1685_in),
    .out(arr__U1685_out)
);
wire [15:0] arr__U1692_in [4:0];
assign arr__U1692_in[4] = arr__U1685_out[4];
assign arr__U1692_in[3] = arr__U1685_out[3];
assign arr__U1692_in[2] = arr__U1685_out[2];
assign arr__U1692_in[1] = arr__U1685_out[1];
assign arr__U1692_in[0] = arr__U1685_out[0];
array_delay_U1693 arr__U1692 (
    .clk(clk),
    .in(arr__U1692_in),
    .out(arr__U1692_out)
);
wire [15:0] arr__U1699_in [4:0];
assign arr__U1699_in[4] = arr__U1692_out[4];
assign arr__U1699_in[3] = arr__U1692_out[3];
assign arr__U1699_in[2] = arr__U1692_out[2];
assign arr__U1699_in[1] = arr__U1692_out[1];
assign arr__U1699_in[0] = arr__U1692_out[0];
array_delay_U1700 arr__U1699 (
    .clk(clk),
    .in(arr__U1699_in),
    .out(arr__U1699_out)
);
wire [15:0] arr__U1706_in [4:0];
assign arr__U1706_in[4] = arr__U1699_out[4];
assign arr__U1706_in[3] = arr__U1699_out[3];
assign arr__U1706_in[2] = arr__U1699_out[2];
assign arr__U1706_in[1] = arr__U1699_out[1];
assign arr__U1706_in[0] = arr__U1699_out[0];
array_delay_U1707 arr__U1706 (
    .clk(clk),
    .in(arr__U1706_in),
    .out(arr__U1706_out)
);
wire [15:0] arr__U1713_in [4:0];
assign arr__U1713_in[4] = arr__U1706_out[4];
assign arr__U1713_in[3] = arr__U1706_out[3];
assign arr__U1713_in[2] = arr__U1706_out[2];
assign arr__U1713_in[1] = arr__U1706_out[1];
assign arr__U1713_in[0] = arr__U1706_out[0];
array_delay_U1714 arr__U1713 (
    .clk(clk),
    .in(arr__U1713_in),
    .out(arr__U1713_out)
);
wire [15:0] arr__U1756_in [4:0];
assign arr__U1756_in[4] = op_hcompute_conv_stencil_15_port_controller_d[4];
assign arr__U1756_in[3] = op_hcompute_conv_stencil_15_port_controller_d[3];
assign arr__U1756_in[2] = op_hcompute_conv_stencil_15_port_controller_d[2];
assign arr__U1756_in[1] = op_hcompute_conv_stencil_15_port_controller_d[1];
assign arr__U1756_in[0] = op_hcompute_conv_stencil_15_port_controller_d[0];
array_delay_U1757 arr__U1756 (
    .clk(clk),
    .in(arr__U1756_in),
    .out(arr__U1756_out)
);
wire [15:0] arr__U1763_in [4:0];
assign arr__U1763_in[4] = arr__U1756_out[4];
assign arr__U1763_in[3] = arr__U1756_out[3];
assign arr__U1763_in[2] = arr__U1756_out[2];
assign arr__U1763_in[1] = arr__U1756_out[1];
assign arr__U1763_in[0] = arr__U1756_out[0];
array_delay_U1764 arr__U1763 (
    .clk(clk),
    .in(arr__U1763_in),
    .out(arr__U1763_out)
);
wire [15:0] arr__U1789_in [4:0];
assign arr__U1789_in[4] = op_hcompute_conv_stencil_15_port_controller_d[4];
assign arr__U1789_in[3] = op_hcompute_conv_stencil_15_port_controller_d[3];
assign arr__U1789_in[2] = op_hcompute_conv_stencil_15_port_controller_d[2];
assign arr__U1789_in[1] = op_hcompute_conv_stencil_15_port_controller_d[1];
assign arr__U1789_in[0] = op_hcompute_conv_stencil_15_port_controller_d[0];
array_delay_U1790 arr__U1789 (
    .clk(clk),
    .in(arr__U1789_in),
    .out(arr__U1789_out)
);
wire [15:0] arr__U1796_in [4:0];
assign arr__U1796_in[4] = arr__U1789_out[4];
assign arr__U1796_in[3] = arr__U1789_out[3];
assign arr__U1796_in[2] = arr__U1789_out[2];
assign arr__U1796_in[1] = arr__U1789_out[1];
assign arr__U1796_in[0] = arr__U1789_out[0];
array_delay_U1797 arr__U1796 (
    .clk(clk),
    .in(arr__U1796_in),
    .out(arr__U1796_out)
);
wire [15:0] arr__U1803_in [4:0];
assign arr__U1803_in[4] = arr__U1796_out[4];
assign arr__U1803_in[3] = arr__U1796_out[3];
assign arr__U1803_in[2] = arr__U1796_out[2];
assign arr__U1803_in[1] = arr__U1796_out[1];
assign arr__U1803_in[0] = arr__U1796_out[0];
array_delay_U1804 arr__U1803 (
    .clk(clk),
    .in(arr__U1803_in),
    .out(arr__U1803_out)
);
wire [15:0] arr__U1810_in [4:0];
assign arr__U1810_in[4] = arr__U1803_out[4];
assign arr__U1810_in[3] = arr__U1803_out[3];
assign arr__U1810_in[2] = arr__U1803_out[2];
assign arr__U1810_in[1] = arr__U1803_out[1];
assign arr__U1810_in[0] = arr__U1803_out[0];
array_delay_U1811 arr__U1810 (
    .clk(clk),
    .in(arr__U1810_in),
    .out(arr__U1810_out)
);
wire [15:0] arr__U1817_in [4:0];
assign arr__U1817_in[4] = arr__U1810_out[4];
assign arr__U1817_in[3] = arr__U1810_out[3];
assign arr__U1817_in[2] = arr__U1810_out[2];
assign arr__U1817_in[1] = arr__U1810_out[1];
assign arr__U1817_in[0] = arr__U1810_out[0];
array_delay_U1818 arr__U1817 (
    .clk(clk),
    .in(arr__U1817_in),
    .out(arr__U1817_out)
);
wire [15:0] arr__U1824_in [4:0];
assign arr__U1824_in[4] = arr__U1817_out[4];
assign arr__U1824_in[3] = arr__U1817_out[3];
assign arr__U1824_in[2] = arr__U1817_out[2];
assign arr__U1824_in[1] = arr__U1817_out[1];
assign arr__U1824_in[0] = arr__U1817_out[0];
array_delay_U1825 arr__U1824 (
    .clk(clk),
    .in(arr__U1824_in),
    .out(arr__U1824_out)
);
wire [15:0] arr__U1831_in [4:0];
assign arr__U1831_in[4] = arr__U1824_out[4];
assign arr__U1831_in[3] = arr__U1824_out[3];
assign arr__U1831_in[2] = arr__U1824_out[2];
assign arr__U1831_in[1] = arr__U1824_out[1];
assign arr__U1831_in[0] = arr__U1824_out[0];
array_delay_U1832 arr__U1831 (
    .clk(clk),
    .in(arr__U1831_in),
    .out(arr__U1831_out)
);
wire [15:0] arr__U1838_in [4:0];
assign arr__U1838_in[4] = arr__U1831_out[4];
assign arr__U1838_in[3] = arr__U1831_out[3];
assign arr__U1838_in[2] = arr__U1831_out[2];
assign arr__U1838_in[1] = arr__U1831_out[1];
assign arr__U1838_in[0] = arr__U1831_out[0];
array_delay_U1839 arr__U1838 (
    .clk(clk),
    .in(arr__U1838_in),
    .out(arr__U1838_out)
);
wire [15:0] arr__U1845_in [4:0];
assign arr__U1845_in[4] = arr__U1838_out[4];
assign arr__U1845_in[3] = arr__U1838_out[3];
assign arr__U1845_in[2] = arr__U1838_out[2];
assign arr__U1845_in[1] = arr__U1838_out[1];
assign arr__U1845_in[0] = arr__U1838_out[0];
array_delay_U1846 arr__U1845 (
    .clk(clk),
    .in(arr__U1845_in),
    .out(arr__U1845_out)
);
wire [15:0] arr__U1852_in [4:0];
assign arr__U1852_in[4] = arr__U1845_out[4];
assign arr__U1852_in[3] = arr__U1845_out[3];
assign arr__U1852_in[2] = arr__U1845_out[2];
assign arr__U1852_in[1] = arr__U1845_out[1];
assign arr__U1852_in[0] = arr__U1845_out[0];
array_delay_U1853 arr__U1852 (
    .clk(clk),
    .in(arr__U1852_in),
    .out(arr__U1852_out)
);
wire [15:0] arr__U1859_in [4:0];
assign arr__U1859_in[4] = arr__U1852_out[4];
assign arr__U1859_in[3] = arr__U1852_out[3];
assign arr__U1859_in[2] = arr__U1852_out[2];
assign arr__U1859_in[1] = arr__U1852_out[1];
assign arr__U1859_in[0] = arr__U1852_out[0];
array_delay_U1860 arr__U1859 (
    .clk(clk),
    .in(arr__U1859_in),
    .out(arr__U1859_out)
);
wire [15:0] arr__U1866_in [4:0];
assign arr__U1866_in[4] = arr__U1859_out[4];
assign arr__U1866_in[3] = arr__U1859_out[3];
assign arr__U1866_in[2] = arr__U1859_out[2];
assign arr__U1866_in[1] = arr__U1859_out[1];
assign arr__U1866_in[0] = arr__U1859_out[0];
array_delay_U1867 arr__U1866 (
    .clk(clk),
    .in(arr__U1866_in),
    .out(arr__U1866_out)
);
wire [15:0] arr__U1873_in [4:0];
assign arr__U1873_in[4] = arr__U1866_out[4];
assign arr__U1873_in[3] = arr__U1866_out[3];
assign arr__U1873_in[2] = arr__U1866_out[2];
assign arr__U1873_in[1] = arr__U1866_out[1];
assign arr__U1873_in[0] = arr__U1866_out[0];
array_delay_U1874 arr__U1873 (
    .clk(clk),
    .in(arr__U1873_in),
    .out(arr__U1873_out)
);
wire [15:0] arr__U1880_in [4:0];
assign arr__U1880_in[4] = arr__U1873_out[4];
assign arr__U1880_in[3] = arr__U1873_out[3];
assign arr__U1880_in[2] = arr__U1873_out[2];
assign arr__U1880_in[1] = arr__U1873_out[1];
assign arr__U1880_in[0] = arr__U1873_out[0];
array_delay_U1881 arr__U1880 (
    .clk(clk),
    .in(arr__U1880_in),
    .out(arr__U1880_out)
);
wire [15:0] arr__U1887_in [4:0];
assign arr__U1887_in[4] = arr__U1880_out[4];
assign arr__U1887_in[3] = arr__U1880_out[3];
assign arr__U1887_in[2] = arr__U1880_out[2];
assign arr__U1887_in[1] = arr__U1880_out[1];
assign arr__U1887_in[0] = arr__U1880_out[0];
array_delay_U1888 arr__U1887 (
    .clk(clk),
    .in(arr__U1887_in),
    .out(arr__U1887_out)
);
wire [15:0] arr__U1894_in [4:0];
assign arr__U1894_in[4] = arr__U1887_out[4];
assign arr__U1894_in[3] = arr__U1887_out[3];
assign arr__U1894_in[2] = arr__U1887_out[2];
assign arr__U1894_in[1] = arr__U1887_out[1];
assign arr__U1894_in[0] = arr__U1887_out[0];
array_delay_U1895 arr__U1894 (
    .clk(clk),
    .in(arr__U1894_in),
    .out(arr__U1894_out)
);
wire [15:0] arr__U1901_in [4:0];
assign arr__U1901_in[4] = arr__U1894_out[4];
assign arr__U1901_in[3] = arr__U1894_out[3];
assign arr__U1901_in[2] = arr__U1894_out[2];
assign arr__U1901_in[1] = arr__U1894_out[1];
assign arr__U1901_in[0] = arr__U1894_out[0];
array_delay_U1902 arr__U1901 (
    .clk(clk),
    .in(arr__U1901_in),
    .out(arr__U1901_out)
);
wire [15:0] arr__U1931_in [2:0];
assign arr__U1931_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U1931_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U1931_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U1932 arr__U1931 (
    .clk(clk),
    .in(arr__U1931_in),
    .out(arr__U1931_out)
);
wire [15:0] arr__U1936_in [2:0];
assign arr__U1936_in[2] = arr__U1931_out[2];
assign arr__U1936_in[1] = arr__U1931_out[1];
assign arr__U1936_in[0] = arr__U1931_out[0];
array_delay_U1937 arr__U1936 (
    .clk(clk),
    .in(arr__U1936_in),
    .out(arr__U1936_out)
);
wire [15:0] arr__U1945_in [2:0];
assign arr__U1945_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U1945_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U1945_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U1946 arr__U1945 (
    .clk(clk),
    .in(arr__U1945_in),
    .out(arr__U1945_out)
);
wire [15:0] arr__U1950_in [2:0];
assign arr__U1950_in[2] = arr__U1945_out[2];
assign arr__U1950_in[1] = arr__U1945_out[1];
assign arr__U1950_in[0] = arr__U1945_out[0];
array_delay_U1951 arr__U1950 (
    .clk(clk),
    .in(arr__U1950_in),
    .out(arr__U1950_out)
);
wire [15:0] arr__U1978_in [2:0];
assign arr__U1978_in[2] = op_hcompute_hw_output_stencil_1_port_controller_d[2];
assign arr__U1978_in[1] = op_hcompute_hw_output_stencil_1_port_controller_d[1];
assign arr__U1978_in[0] = op_hcompute_hw_output_stencil_1_port_controller_d[0];
array_delay_U1979 arr__U1978 (
    .clk(clk),
    .in(arr__U1978_in),
    .out(arr__U1978_out)
);
wire [15:0] arr__U1983_in [2:0];
assign arr__U1983_in[2] = arr__U1978_out[2];
assign arr__U1983_in[1] = arr__U1978_out[1];
assign arr__U1983_in[0] = arr__U1978_out[0];
array_delay_U1984 arr__U1983 (
    .clk(clk),
    .in(arr__U1983_in),
    .out(arr__U1983_out)
);
wire [15:0] arr__U1992_in [2:0];
assign arr__U1992_in[2] = op_hcompute_hw_output_stencil_1_port_controller_d[2];
assign arr__U1992_in[1] = op_hcompute_hw_output_stencil_1_port_controller_d[1];
assign arr__U1992_in[0] = op_hcompute_hw_output_stencil_1_port_controller_d[0];
array_delay_U1993 arr__U1992 (
    .clk(clk),
    .in(arr__U1992_in),
    .out(arr__U1992_out)
);
wire [15:0] arr__U1997_in [2:0];
assign arr__U1997_in[2] = arr__U1992_out[2];
assign arr__U1997_in[1] = arr__U1992_out[1];
assign arr__U1997_in[0] = arr__U1992_out[0];
array_delay_U1998 arr__U1997 (
    .clk(clk),
    .in(arr__U1997_in),
    .out(arr__U1997_out)
);
wire [15:0] arr__U2025_in [2:0];
assign arr__U2025_in[2] = op_hcompute_hw_output_stencil_2_port_controller_d[2];
assign arr__U2025_in[1] = op_hcompute_hw_output_stencil_2_port_controller_d[1];
assign arr__U2025_in[0] = op_hcompute_hw_output_stencil_2_port_controller_d[0];
array_delay_U2026 arr__U2025 (
    .clk(clk),
    .in(arr__U2025_in),
    .out(arr__U2025_out)
);
wire [15:0] arr__U2030_in [2:0];
assign arr__U2030_in[2] = arr__U2025_out[2];
assign arr__U2030_in[1] = arr__U2025_out[1];
assign arr__U2030_in[0] = arr__U2025_out[0];
array_delay_U2031 arr__U2030 (
    .clk(clk),
    .in(arr__U2030_in),
    .out(arr__U2030_out)
);
wire [15:0] arr__U2039_in [2:0];
assign arr__U2039_in[2] = op_hcompute_hw_output_stencil_2_port_controller_d[2];
assign arr__U2039_in[1] = op_hcompute_hw_output_stencil_2_port_controller_d[1];
assign arr__U2039_in[0] = op_hcompute_hw_output_stencil_2_port_controller_d[0];
array_delay_U2040 arr__U2039 (
    .clk(clk),
    .in(arr__U2039_in),
    .out(arr__U2039_out)
);
wire [15:0] arr__U2044_in [2:0];
assign arr__U2044_in[2] = arr__U2039_out[2];
assign arr__U2044_in[1] = arr__U2039_out[1];
assign arr__U2044_in[0] = arr__U2039_out[0];
array_delay_U2045 arr__U2044 (
    .clk(clk),
    .in(arr__U2044_in),
    .out(arr__U2044_out)
);
wire [15:0] arr__U2072_in [2:0];
assign arr__U2072_in[2] = op_hcompute_hw_output_stencil_3_port_controller_d[2];
assign arr__U2072_in[1] = op_hcompute_hw_output_stencil_3_port_controller_d[1];
assign arr__U2072_in[0] = op_hcompute_hw_output_stencil_3_port_controller_d[0];
array_delay_U2073 arr__U2072 (
    .clk(clk),
    .in(arr__U2072_in),
    .out(arr__U2072_out)
);
wire [15:0] arr__U2077_in [2:0];
assign arr__U2077_in[2] = arr__U2072_out[2];
assign arr__U2077_in[1] = arr__U2072_out[1];
assign arr__U2077_in[0] = arr__U2072_out[0];
array_delay_U2078 arr__U2077 (
    .clk(clk),
    .in(arr__U2077_in),
    .out(arr__U2077_out)
);
wire [15:0] arr__U2086_in [2:0];
assign arr__U2086_in[2] = op_hcompute_hw_output_stencil_3_port_controller_d[2];
assign arr__U2086_in[1] = op_hcompute_hw_output_stencil_3_port_controller_d[1];
assign arr__U2086_in[0] = op_hcompute_hw_output_stencil_3_port_controller_d[0];
array_delay_U2087 arr__U2086 (
    .clk(clk),
    .in(arr__U2086_in),
    .out(arr__U2086_out)
);
wire [15:0] arr__U2091_in [2:0];
assign arr__U2091_in[2] = arr__U2086_out[2];
assign arr__U2091_in[1] = arr__U2086_out[1];
assign arr__U2091_in[0] = arr__U2086_out[0];
array_delay_U2092 arr__U2091 (
    .clk(clk),
    .in(arr__U2091_in),
    .out(arr__U2091_out)
);
wire [15:0] arr__U2119_in [2:0];
assign arr__U2119_in[2] = op_hcompute_hw_output_stencil_4_port_controller_d[2];
assign arr__U2119_in[1] = op_hcompute_hw_output_stencil_4_port_controller_d[1];
assign arr__U2119_in[0] = op_hcompute_hw_output_stencil_4_port_controller_d[0];
array_delay_U2120 arr__U2119 (
    .clk(clk),
    .in(arr__U2119_in),
    .out(arr__U2119_out)
);
wire [15:0] arr__U2124_in [2:0];
assign arr__U2124_in[2] = arr__U2119_out[2];
assign arr__U2124_in[1] = arr__U2119_out[1];
assign arr__U2124_in[0] = arr__U2119_out[0];
array_delay_U2125 arr__U2124 (
    .clk(clk),
    .in(arr__U2124_in),
    .out(arr__U2124_out)
);
wire [15:0] arr__U2133_in [2:0];
assign arr__U2133_in[2] = op_hcompute_hw_output_stencil_4_port_controller_d[2];
assign arr__U2133_in[1] = op_hcompute_hw_output_stencil_4_port_controller_d[1];
assign arr__U2133_in[0] = op_hcompute_hw_output_stencil_4_port_controller_d[0];
array_delay_U2134 arr__U2133 (
    .clk(clk),
    .in(arr__U2133_in),
    .out(arr__U2133_out)
);
wire [15:0] arr__U2138_in [2:0];
assign arr__U2138_in[2] = arr__U2133_out[2];
assign arr__U2138_in[1] = arr__U2133_out[1];
assign arr__U2138_in[0] = arr__U2133_out[0];
array_delay_U2139 arr__U2138 (
    .clk(clk),
    .in(arr__U2138_in),
    .out(arr__U2138_out)
);
wire [15:0] arr__U2166_in [2:0];
assign arr__U2166_in[2] = op_hcompute_hw_output_stencil_5_port_controller_d[2];
assign arr__U2166_in[1] = op_hcompute_hw_output_stencil_5_port_controller_d[1];
assign arr__U2166_in[0] = op_hcompute_hw_output_stencil_5_port_controller_d[0];
array_delay_U2167 arr__U2166 (
    .clk(clk),
    .in(arr__U2166_in),
    .out(arr__U2166_out)
);
wire [15:0] arr__U2171_in [2:0];
assign arr__U2171_in[2] = arr__U2166_out[2];
assign arr__U2171_in[1] = arr__U2166_out[1];
assign arr__U2171_in[0] = arr__U2166_out[0];
array_delay_U2172 arr__U2171 (
    .clk(clk),
    .in(arr__U2171_in),
    .out(arr__U2171_out)
);
wire [15:0] arr__U2180_in [2:0];
assign arr__U2180_in[2] = op_hcompute_hw_output_stencil_5_port_controller_d[2];
assign arr__U2180_in[1] = op_hcompute_hw_output_stencil_5_port_controller_d[1];
assign arr__U2180_in[0] = op_hcompute_hw_output_stencil_5_port_controller_d[0];
array_delay_U2181 arr__U2180 (
    .clk(clk),
    .in(arr__U2180_in),
    .out(arr__U2180_out)
);
wire [15:0] arr__U2185_in [2:0];
assign arr__U2185_in[2] = arr__U2180_out[2];
assign arr__U2185_in[1] = arr__U2180_out[1];
assign arr__U2185_in[0] = arr__U2180_out[0];
array_delay_U2186 arr__U2185 (
    .clk(clk),
    .in(arr__U2185_in),
    .out(arr__U2185_out)
);
wire [15:0] arr__U2213_in [2:0];
assign arr__U2213_in[2] = op_hcompute_hw_output_stencil_6_port_controller_d[2];
assign arr__U2213_in[1] = op_hcompute_hw_output_stencil_6_port_controller_d[1];
assign arr__U2213_in[0] = op_hcompute_hw_output_stencil_6_port_controller_d[0];
array_delay_U2214 arr__U2213 (
    .clk(clk),
    .in(arr__U2213_in),
    .out(arr__U2213_out)
);
wire [15:0] arr__U2218_in [2:0];
assign arr__U2218_in[2] = arr__U2213_out[2];
assign arr__U2218_in[1] = arr__U2213_out[1];
assign arr__U2218_in[0] = arr__U2213_out[0];
array_delay_U2219 arr__U2218 (
    .clk(clk),
    .in(arr__U2218_in),
    .out(arr__U2218_out)
);
wire [15:0] arr__U2227_in [2:0];
assign arr__U2227_in[2] = op_hcompute_hw_output_stencil_6_port_controller_d[2];
assign arr__U2227_in[1] = op_hcompute_hw_output_stencil_6_port_controller_d[1];
assign arr__U2227_in[0] = op_hcompute_hw_output_stencil_6_port_controller_d[0];
array_delay_U2228 arr__U2227 (
    .clk(clk),
    .in(arr__U2227_in),
    .out(arr__U2227_out)
);
wire [15:0] arr__U2232_in [2:0];
assign arr__U2232_in[2] = arr__U2227_out[2];
assign arr__U2232_in[1] = arr__U2227_out[1];
assign arr__U2232_in[0] = arr__U2227_out[0];
array_delay_U2233 arr__U2232 (
    .clk(clk),
    .in(arr__U2232_in),
    .out(arr__U2232_out)
);
wire [15:0] arr__U2260_in [2:0];
assign arr__U2260_in[2] = op_hcompute_hw_output_stencil_7_port_controller_d[2];
assign arr__U2260_in[1] = op_hcompute_hw_output_stencil_7_port_controller_d[1];
assign arr__U2260_in[0] = op_hcompute_hw_output_stencil_7_port_controller_d[0];
array_delay_U2261 arr__U2260 (
    .clk(clk),
    .in(arr__U2260_in),
    .out(arr__U2260_out)
);
wire [15:0] arr__U2265_in [2:0];
assign arr__U2265_in[2] = arr__U2260_out[2];
assign arr__U2265_in[1] = arr__U2260_out[1];
assign arr__U2265_in[0] = arr__U2260_out[0];
array_delay_U2266 arr__U2265 (
    .clk(clk),
    .in(arr__U2265_in),
    .out(arr__U2265_out)
);
wire [15:0] arr__U2274_in [2:0];
assign arr__U2274_in[2] = op_hcompute_hw_output_stencil_7_port_controller_d[2];
assign arr__U2274_in[1] = op_hcompute_hw_output_stencil_7_port_controller_d[1];
assign arr__U2274_in[0] = op_hcompute_hw_output_stencil_7_port_controller_d[0];
array_delay_U2275 arr__U2274 (
    .clk(clk),
    .in(arr__U2274_in),
    .out(arr__U2274_out)
);
wire [15:0] arr__U2279_in [2:0];
assign arr__U2279_in[2] = arr__U2274_out[2];
assign arr__U2279_in[1] = arr__U2274_out[1];
assign arr__U2279_in[0] = arr__U2274_out[0];
array_delay_U2280 arr__U2279 (
    .clk(clk),
    .in(arr__U2279_in),
    .out(arr__U2279_out)
);
wire [15:0] arr__U440_in [4:0];
assign arr__U440_in[4] = op_hcompute_conv_stencil_8_port_controller_d[4];
assign arr__U440_in[3] = op_hcompute_conv_stencil_8_port_controller_d[3];
assign arr__U440_in[2] = op_hcompute_conv_stencil_8_port_controller_d[2];
assign arr__U440_in[1] = op_hcompute_conv_stencil_8_port_controller_d[1];
assign arr__U440_in[0] = op_hcompute_conv_stencil_8_port_controller_d[0];
array_delay_U441 arr__U440 (
    .clk(clk),
    .in(arr__U440_in),
    .out(arr__U440_out)
);
wire [15:0] arr__U447_in [4:0];
assign arr__U447_in[4] = arr__U440_out[4];
assign arr__U447_in[3] = arr__U440_out[3];
assign arr__U447_in[2] = arr__U440_out[2];
assign arr__U447_in[1] = arr__U440_out[1];
assign arr__U447_in[0] = arr__U440_out[0];
array_delay_U448 arr__U447 (
    .clk(clk),
    .in(arr__U447_in),
    .out(arr__U447_out)
);
wire [15:0] arr__U473_in [4:0];
assign arr__U473_in[4] = op_hcompute_conv_stencil_8_port_controller_d[4];
assign arr__U473_in[3] = op_hcompute_conv_stencil_8_port_controller_d[3];
assign arr__U473_in[2] = op_hcompute_conv_stencil_8_port_controller_d[2];
assign arr__U473_in[1] = op_hcompute_conv_stencil_8_port_controller_d[1];
assign arr__U473_in[0] = op_hcompute_conv_stencil_8_port_controller_d[0];
array_delay_U474 arr__U473 (
    .clk(clk),
    .in(arr__U473_in),
    .out(arr__U473_out)
);
wire [15:0] arr__U480_in [4:0];
assign arr__U480_in[4] = arr__U473_out[4];
assign arr__U480_in[3] = arr__U473_out[3];
assign arr__U480_in[2] = arr__U473_out[2];
assign arr__U480_in[1] = arr__U473_out[1];
assign arr__U480_in[0] = arr__U473_out[0];
array_delay_U481 arr__U480 (
    .clk(clk),
    .in(arr__U480_in),
    .out(arr__U480_out)
);
wire [15:0] arr__U487_in [4:0];
assign arr__U487_in[4] = arr__U480_out[4];
assign arr__U487_in[3] = arr__U480_out[3];
assign arr__U487_in[2] = arr__U480_out[2];
assign arr__U487_in[1] = arr__U480_out[1];
assign arr__U487_in[0] = arr__U480_out[0];
array_delay_U488 arr__U487 (
    .clk(clk),
    .in(arr__U487_in),
    .out(arr__U487_out)
);
wire [15:0] arr__U494_in [4:0];
assign arr__U494_in[4] = arr__U487_out[4];
assign arr__U494_in[3] = arr__U487_out[3];
assign arr__U494_in[2] = arr__U487_out[2];
assign arr__U494_in[1] = arr__U487_out[1];
assign arr__U494_in[0] = arr__U487_out[0];
array_delay_U495 arr__U494 (
    .clk(clk),
    .in(arr__U494_in),
    .out(arr__U494_out)
);
wire [15:0] arr__U501_in [4:0];
assign arr__U501_in[4] = arr__U494_out[4];
assign arr__U501_in[3] = arr__U494_out[3];
assign arr__U501_in[2] = arr__U494_out[2];
assign arr__U501_in[1] = arr__U494_out[1];
assign arr__U501_in[0] = arr__U494_out[0];
array_delay_U502 arr__U501 (
    .clk(clk),
    .in(arr__U501_in),
    .out(arr__U501_out)
);
wire [15:0] arr__U508_in [4:0];
assign arr__U508_in[4] = arr__U501_out[4];
assign arr__U508_in[3] = arr__U501_out[3];
assign arr__U508_in[2] = arr__U501_out[2];
assign arr__U508_in[1] = arr__U501_out[1];
assign arr__U508_in[0] = arr__U501_out[0];
array_delay_U509 arr__U508 (
    .clk(clk),
    .in(arr__U508_in),
    .out(arr__U508_out)
);
wire [15:0] arr__U515_in [4:0];
assign arr__U515_in[4] = arr__U508_out[4];
assign arr__U515_in[3] = arr__U508_out[3];
assign arr__U515_in[2] = arr__U508_out[2];
assign arr__U515_in[1] = arr__U508_out[1];
assign arr__U515_in[0] = arr__U508_out[0];
array_delay_U516 arr__U515 (
    .clk(clk),
    .in(arr__U515_in),
    .out(arr__U515_out)
);
wire [15:0] arr__U522_in [4:0];
assign arr__U522_in[4] = arr__U515_out[4];
assign arr__U522_in[3] = arr__U515_out[3];
assign arr__U522_in[2] = arr__U515_out[2];
assign arr__U522_in[1] = arr__U515_out[1];
assign arr__U522_in[0] = arr__U515_out[0];
array_delay_U523 arr__U522 (
    .clk(clk),
    .in(arr__U522_in),
    .out(arr__U522_out)
);
wire [15:0] arr__U529_in [4:0];
assign arr__U529_in[4] = arr__U522_out[4];
assign arr__U529_in[3] = arr__U522_out[3];
assign arr__U529_in[2] = arr__U522_out[2];
assign arr__U529_in[1] = arr__U522_out[1];
assign arr__U529_in[0] = arr__U522_out[0];
array_delay_U530 arr__U529 (
    .clk(clk),
    .in(arr__U529_in),
    .out(arr__U529_out)
);
wire [15:0] arr__U536_in [4:0];
assign arr__U536_in[4] = arr__U529_out[4];
assign arr__U536_in[3] = arr__U529_out[3];
assign arr__U536_in[2] = arr__U529_out[2];
assign arr__U536_in[1] = arr__U529_out[1];
assign arr__U536_in[0] = arr__U529_out[0];
array_delay_U537 arr__U536 (
    .clk(clk),
    .in(arr__U536_in),
    .out(arr__U536_out)
);
wire [15:0] arr__U543_in [4:0];
assign arr__U543_in[4] = arr__U536_out[4];
assign arr__U543_in[3] = arr__U536_out[3];
assign arr__U543_in[2] = arr__U536_out[2];
assign arr__U543_in[1] = arr__U536_out[1];
assign arr__U543_in[0] = arr__U536_out[0];
array_delay_U544 arr__U543 (
    .clk(clk),
    .in(arr__U543_in),
    .out(arr__U543_out)
);
wire [15:0] arr__U550_in [4:0];
assign arr__U550_in[4] = arr__U543_out[4];
assign arr__U550_in[3] = arr__U543_out[3];
assign arr__U550_in[2] = arr__U543_out[2];
assign arr__U550_in[1] = arr__U543_out[1];
assign arr__U550_in[0] = arr__U543_out[0];
array_delay_U551 arr__U550 (
    .clk(clk),
    .in(arr__U550_in),
    .out(arr__U550_out)
);
wire [15:0] arr__U557_in [4:0];
assign arr__U557_in[4] = arr__U550_out[4];
assign arr__U557_in[3] = arr__U550_out[3];
assign arr__U557_in[2] = arr__U550_out[2];
assign arr__U557_in[1] = arr__U550_out[1];
assign arr__U557_in[0] = arr__U550_out[0];
array_delay_U558 arr__U557 (
    .clk(clk),
    .in(arr__U557_in),
    .out(arr__U557_out)
);
wire [15:0] arr__U564_in [4:0];
assign arr__U564_in[4] = arr__U557_out[4];
assign arr__U564_in[3] = arr__U557_out[3];
assign arr__U564_in[2] = arr__U557_out[2];
assign arr__U564_in[1] = arr__U557_out[1];
assign arr__U564_in[0] = arr__U557_out[0];
array_delay_U565 arr__U564 (
    .clk(clk),
    .in(arr__U564_in),
    .out(arr__U564_out)
);
wire [15:0] arr__U571_in [4:0];
assign arr__U571_in[4] = arr__U564_out[4];
assign arr__U571_in[3] = arr__U564_out[3];
assign arr__U571_in[2] = arr__U564_out[2];
assign arr__U571_in[1] = arr__U564_out[1];
assign arr__U571_in[0] = arr__U564_out[0];
array_delay_U572 arr__U571 (
    .clk(clk),
    .in(arr__U571_in),
    .out(arr__U571_out)
);
wire [15:0] arr__U578_in [4:0];
assign arr__U578_in[4] = arr__U571_out[4];
assign arr__U578_in[3] = arr__U571_out[3];
assign arr__U578_in[2] = arr__U571_out[2];
assign arr__U578_in[1] = arr__U571_out[1];
assign arr__U578_in[0] = arr__U571_out[0];
array_delay_U579 arr__U578 (
    .clk(clk),
    .in(arr__U578_in),
    .out(arr__U578_out)
);
wire [15:0] arr__U585_in [4:0];
assign arr__U585_in[4] = arr__U578_out[4];
assign arr__U585_in[3] = arr__U578_out[3];
assign arr__U585_in[2] = arr__U578_out[2];
assign arr__U585_in[1] = arr__U578_out[1];
assign arr__U585_in[0] = arr__U578_out[0];
array_delay_U586 arr__U585 (
    .clk(clk),
    .in(arr__U585_in),
    .out(arr__U585_out)
);
wire [15:0] arr__U628_in [4:0];
assign arr__U628_in[4] = op_hcompute_conv_stencil_9_port_controller_d[4];
assign arr__U628_in[3] = op_hcompute_conv_stencil_9_port_controller_d[3];
assign arr__U628_in[2] = op_hcompute_conv_stencil_9_port_controller_d[2];
assign arr__U628_in[1] = op_hcompute_conv_stencil_9_port_controller_d[1];
assign arr__U628_in[0] = op_hcompute_conv_stencil_9_port_controller_d[0];
array_delay_U629 arr__U628 (
    .clk(clk),
    .in(arr__U628_in),
    .out(arr__U628_out)
);
wire [15:0] arr__U635_in [4:0];
assign arr__U635_in[4] = arr__U628_out[4];
assign arr__U635_in[3] = arr__U628_out[3];
assign arr__U635_in[2] = arr__U628_out[2];
assign arr__U635_in[1] = arr__U628_out[1];
assign arr__U635_in[0] = arr__U628_out[0];
array_delay_U636 arr__U635 (
    .clk(clk),
    .in(arr__U635_in),
    .out(arr__U635_out)
);
wire [15:0] arr__U661_in [4:0];
assign arr__U661_in[4] = op_hcompute_conv_stencil_9_port_controller_d[4];
assign arr__U661_in[3] = op_hcompute_conv_stencil_9_port_controller_d[3];
assign arr__U661_in[2] = op_hcompute_conv_stencil_9_port_controller_d[2];
assign arr__U661_in[1] = op_hcompute_conv_stencil_9_port_controller_d[1];
assign arr__U661_in[0] = op_hcompute_conv_stencil_9_port_controller_d[0];
array_delay_U662 arr__U661 (
    .clk(clk),
    .in(arr__U661_in),
    .out(arr__U661_out)
);
wire [15:0] arr__U668_in [4:0];
assign arr__U668_in[4] = arr__U661_out[4];
assign arr__U668_in[3] = arr__U661_out[3];
assign arr__U668_in[2] = arr__U661_out[2];
assign arr__U668_in[1] = arr__U661_out[1];
assign arr__U668_in[0] = arr__U661_out[0];
array_delay_U669 arr__U668 (
    .clk(clk),
    .in(arr__U668_in),
    .out(arr__U668_out)
);
wire [15:0] arr__U675_in [4:0];
assign arr__U675_in[4] = arr__U668_out[4];
assign arr__U675_in[3] = arr__U668_out[3];
assign arr__U675_in[2] = arr__U668_out[2];
assign arr__U675_in[1] = arr__U668_out[1];
assign arr__U675_in[0] = arr__U668_out[0];
array_delay_U676 arr__U675 (
    .clk(clk),
    .in(arr__U675_in),
    .out(arr__U675_out)
);
wire [15:0] arr__U682_in [4:0];
assign arr__U682_in[4] = arr__U675_out[4];
assign arr__U682_in[3] = arr__U675_out[3];
assign arr__U682_in[2] = arr__U675_out[2];
assign arr__U682_in[1] = arr__U675_out[1];
assign arr__U682_in[0] = arr__U675_out[0];
array_delay_U683 arr__U682 (
    .clk(clk),
    .in(arr__U682_in),
    .out(arr__U682_out)
);
wire [15:0] arr__U689_in [4:0];
assign arr__U689_in[4] = arr__U682_out[4];
assign arr__U689_in[3] = arr__U682_out[3];
assign arr__U689_in[2] = arr__U682_out[2];
assign arr__U689_in[1] = arr__U682_out[1];
assign arr__U689_in[0] = arr__U682_out[0];
array_delay_U690 arr__U689 (
    .clk(clk),
    .in(arr__U689_in),
    .out(arr__U689_out)
);
wire [15:0] arr__U696_in [4:0];
assign arr__U696_in[4] = arr__U689_out[4];
assign arr__U696_in[3] = arr__U689_out[3];
assign arr__U696_in[2] = arr__U689_out[2];
assign arr__U696_in[1] = arr__U689_out[1];
assign arr__U696_in[0] = arr__U689_out[0];
array_delay_U697 arr__U696 (
    .clk(clk),
    .in(arr__U696_in),
    .out(arr__U696_out)
);
wire [15:0] arr__U703_in [4:0];
assign arr__U703_in[4] = arr__U696_out[4];
assign arr__U703_in[3] = arr__U696_out[3];
assign arr__U703_in[2] = arr__U696_out[2];
assign arr__U703_in[1] = arr__U696_out[1];
assign arr__U703_in[0] = arr__U696_out[0];
array_delay_U704 arr__U703 (
    .clk(clk),
    .in(arr__U703_in),
    .out(arr__U703_out)
);
wire [15:0] arr__U710_in [4:0];
assign arr__U710_in[4] = arr__U703_out[4];
assign arr__U710_in[3] = arr__U703_out[3];
assign arr__U710_in[2] = arr__U703_out[2];
assign arr__U710_in[1] = arr__U703_out[1];
assign arr__U710_in[0] = arr__U703_out[0];
array_delay_U711 arr__U710 (
    .clk(clk),
    .in(arr__U710_in),
    .out(arr__U710_out)
);
wire [15:0] arr__U717_in [4:0];
assign arr__U717_in[4] = arr__U710_out[4];
assign arr__U717_in[3] = arr__U710_out[3];
assign arr__U717_in[2] = arr__U710_out[2];
assign arr__U717_in[1] = arr__U710_out[1];
assign arr__U717_in[0] = arr__U710_out[0];
array_delay_U718 arr__U717 (
    .clk(clk),
    .in(arr__U717_in),
    .out(arr__U717_out)
);
wire [15:0] arr__U724_in [4:0];
assign arr__U724_in[4] = arr__U717_out[4];
assign arr__U724_in[3] = arr__U717_out[3];
assign arr__U724_in[2] = arr__U717_out[2];
assign arr__U724_in[1] = arr__U717_out[1];
assign arr__U724_in[0] = arr__U717_out[0];
array_delay_U725 arr__U724 (
    .clk(clk),
    .in(arr__U724_in),
    .out(arr__U724_out)
);
wire [15:0] arr__U731_in [4:0];
assign arr__U731_in[4] = arr__U724_out[4];
assign arr__U731_in[3] = arr__U724_out[3];
assign arr__U731_in[2] = arr__U724_out[2];
assign arr__U731_in[1] = arr__U724_out[1];
assign arr__U731_in[0] = arr__U724_out[0];
array_delay_U732 arr__U731 (
    .clk(clk),
    .in(arr__U731_in),
    .out(arr__U731_out)
);
wire [15:0] arr__U738_in [4:0];
assign arr__U738_in[4] = arr__U731_out[4];
assign arr__U738_in[3] = arr__U731_out[3];
assign arr__U738_in[2] = arr__U731_out[2];
assign arr__U738_in[1] = arr__U731_out[1];
assign arr__U738_in[0] = arr__U731_out[0];
array_delay_U739 arr__U738 (
    .clk(clk),
    .in(arr__U738_in),
    .out(arr__U738_out)
);
wire [15:0] arr__U745_in [4:0];
assign arr__U745_in[4] = arr__U738_out[4];
assign arr__U745_in[3] = arr__U738_out[3];
assign arr__U745_in[2] = arr__U738_out[2];
assign arr__U745_in[1] = arr__U738_out[1];
assign arr__U745_in[0] = arr__U738_out[0];
array_delay_U746 arr__U745 (
    .clk(clk),
    .in(arr__U745_in),
    .out(arr__U745_out)
);
wire [15:0] arr__U752_in [4:0];
assign arr__U752_in[4] = arr__U745_out[4];
assign arr__U752_in[3] = arr__U745_out[3];
assign arr__U752_in[2] = arr__U745_out[2];
assign arr__U752_in[1] = arr__U745_out[1];
assign arr__U752_in[0] = arr__U745_out[0];
array_delay_U753 arr__U752 (
    .clk(clk),
    .in(arr__U752_in),
    .out(arr__U752_out)
);
wire [15:0] arr__U759_in [4:0];
assign arr__U759_in[4] = arr__U752_out[4];
assign arr__U759_in[3] = arr__U752_out[3];
assign arr__U759_in[2] = arr__U752_out[2];
assign arr__U759_in[1] = arr__U752_out[1];
assign arr__U759_in[0] = arr__U752_out[0];
array_delay_U760 arr__U759 (
    .clk(clk),
    .in(arr__U759_in),
    .out(arr__U759_out)
);
wire [15:0] arr__U766_in [4:0];
assign arr__U766_in[4] = arr__U759_out[4];
assign arr__U766_in[3] = arr__U759_out[3];
assign arr__U766_in[2] = arr__U759_out[2];
assign arr__U766_in[1] = arr__U759_out[1];
assign arr__U766_in[0] = arr__U759_out[0];
array_delay_U767 arr__U766 (
    .clk(clk),
    .in(arr__U766_in),
    .out(arr__U766_out)
);
wire [15:0] arr__U773_in [4:0];
assign arr__U773_in[4] = arr__U766_out[4];
assign arr__U773_in[3] = arr__U766_out[3];
assign arr__U773_in[2] = arr__U766_out[2];
assign arr__U773_in[1] = arr__U766_out[1];
assign arr__U773_in[0] = arr__U766_out[0];
array_delay_U774 arr__U773 (
    .clk(clk),
    .in(arr__U773_in),
    .out(arr__U773_out)
);
wire [15:0] arr__U816_in [4:0];
assign arr__U816_in[4] = op_hcompute_conv_stencil_10_port_controller_d[4];
assign arr__U816_in[3] = op_hcompute_conv_stencil_10_port_controller_d[3];
assign arr__U816_in[2] = op_hcompute_conv_stencil_10_port_controller_d[2];
assign arr__U816_in[1] = op_hcompute_conv_stencil_10_port_controller_d[1];
assign arr__U816_in[0] = op_hcompute_conv_stencil_10_port_controller_d[0];
array_delay_U817 arr__U816 (
    .clk(clk),
    .in(arr__U816_in),
    .out(arr__U816_out)
);
wire [15:0] arr__U823_in [4:0];
assign arr__U823_in[4] = arr__U816_out[4];
assign arr__U823_in[3] = arr__U816_out[3];
assign arr__U823_in[2] = arr__U816_out[2];
assign arr__U823_in[1] = arr__U816_out[1];
assign arr__U823_in[0] = arr__U816_out[0];
array_delay_U824 arr__U823 (
    .clk(clk),
    .in(arr__U823_in),
    .out(arr__U823_out)
);
wire [15:0] arr__U849_in [4:0];
assign arr__U849_in[4] = op_hcompute_conv_stencil_10_port_controller_d[4];
assign arr__U849_in[3] = op_hcompute_conv_stencil_10_port_controller_d[3];
assign arr__U849_in[2] = op_hcompute_conv_stencil_10_port_controller_d[2];
assign arr__U849_in[1] = op_hcompute_conv_stencil_10_port_controller_d[1];
assign arr__U849_in[0] = op_hcompute_conv_stencil_10_port_controller_d[0];
array_delay_U850 arr__U849 (
    .clk(clk),
    .in(arr__U849_in),
    .out(arr__U849_out)
);
wire [15:0] arr__U856_in [4:0];
assign arr__U856_in[4] = arr__U849_out[4];
assign arr__U856_in[3] = arr__U849_out[3];
assign arr__U856_in[2] = arr__U849_out[2];
assign arr__U856_in[1] = arr__U849_out[1];
assign arr__U856_in[0] = arr__U849_out[0];
array_delay_U857 arr__U856 (
    .clk(clk),
    .in(arr__U856_in),
    .out(arr__U856_out)
);
wire [15:0] arr__U863_in [4:0];
assign arr__U863_in[4] = arr__U856_out[4];
assign arr__U863_in[3] = arr__U856_out[3];
assign arr__U863_in[2] = arr__U856_out[2];
assign arr__U863_in[1] = arr__U856_out[1];
assign arr__U863_in[0] = arr__U856_out[0];
array_delay_U864 arr__U863 (
    .clk(clk),
    .in(arr__U863_in),
    .out(arr__U863_out)
);
wire [15:0] arr__U870_in [4:0];
assign arr__U870_in[4] = arr__U863_out[4];
assign arr__U870_in[3] = arr__U863_out[3];
assign arr__U870_in[2] = arr__U863_out[2];
assign arr__U870_in[1] = arr__U863_out[1];
assign arr__U870_in[0] = arr__U863_out[0];
array_delay_U871 arr__U870 (
    .clk(clk),
    .in(arr__U870_in),
    .out(arr__U870_out)
);
wire [15:0] arr__U877_in [4:0];
assign arr__U877_in[4] = arr__U870_out[4];
assign arr__U877_in[3] = arr__U870_out[3];
assign arr__U877_in[2] = arr__U870_out[2];
assign arr__U877_in[1] = arr__U870_out[1];
assign arr__U877_in[0] = arr__U870_out[0];
array_delay_U878 arr__U877 (
    .clk(clk),
    .in(arr__U877_in),
    .out(arr__U877_out)
);
wire [15:0] arr__U884_in [4:0];
assign arr__U884_in[4] = arr__U877_out[4];
assign arr__U884_in[3] = arr__U877_out[3];
assign arr__U884_in[2] = arr__U877_out[2];
assign arr__U884_in[1] = arr__U877_out[1];
assign arr__U884_in[0] = arr__U877_out[0];
array_delay_U885 arr__U884 (
    .clk(clk),
    .in(arr__U884_in),
    .out(arr__U884_out)
);
wire [15:0] arr__U891_in [4:0];
assign arr__U891_in[4] = arr__U884_out[4];
assign arr__U891_in[3] = arr__U884_out[3];
assign arr__U891_in[2] = arr__U884_out[2];
assign arr__U891_in[1] = arr__U884_out[1];
assign arr__U891_in[0] = arr__U884_out[0];
array_delay_U892 arr__U891 (
    .clk(clk),
    .in(arr__U891_in),
    .out(arr__U891_out)
);
wire [15:0] arr__U898_in [4:0];
assign arr__U898_in[4] = arr__U891_out[4];
assign arr__U898_in[3] = arr__U891_out[3];
assign arr__U898_in[2] = arr__U891_out[2];
assign arr__U898_in[1] = arr__U891_out[1];
assign arr__U898_in[0] = arr__U891_out[0];
array_delay_U899 arr__U898 (
    .clk(clk),
    .in(arr__U898_in),
    .out(arr__U898_out)
);
wire [15:0] arr__U905_in [4:0];
assign arr__U905_in[4] = arr__U898_out[4];
assign arr__U905_in[3] = arr__U898_out[3];
assign arr__U905_in[2] = arr__U898_out[2];
assign arr__U905_in[1] = arr__U898_out[1];
assign arr__U905_in[0] = arr__U898_out[0];
array_delay_U906 arr__U905 (
    .clk(clk),
    .in(arr__U905_in),
    .out(arr__U905_out)
);
wire [15:0] arr__U912_in [4:0];
assign arr__U912_in[4] = arr__U905_out[4];
assign arr__U912_in[3] = arr__U905_out[3];
assign arr__U912_in[2] = arr__U905_out[2];
assign arr__U912_in[1] = arr__U905_out[1];
assign arr__U912_in[0] = arr__U905_out[0];
array_delay_U913 arr__U912 (
    .clk(clk),
    .in(arr__U912_in),
    .out(arr__U912_out)
);
wire [15:0] arr__U919_in [4:0];
assign arr__U919_in[4] = arr__U912_out[4];
assign arr__U919_in[3] = arr__U912_out[3];
assign arr__U919_in[2] = arr__U912_out[2];
assign arr__U919_in[1] = arr__U912_out[1];
assign arr__U919_in[0] = arr__U912_out[0];
array_delay_U920 arr__U919 (
    .clk(clk),
    .in(arr__U919_in),
    .out(arr__U919_out)
);
wire [15:0] arr__U926_in [4:0];
assign arr__U926_in[4] = arr__U919_out[4];
assign arr__U926_in[3] = arr__U919_out[3];
assign arr__U926_in[2] = arr__U919_out[2];
assign arr__U926_in[1] = arr__U919_out[1];
assign arr__U926_in[0] = arr__U919_out[0];
array_delay_U927 arr__U926 (
    .clk(clk),
    .in(arr__U926_in),
    .out(arr__U926_out)
);
wire [15:0] arr__U933_in [4:0];
assign arr__U933_in[4] = arr__U926_out[4];
assign arr__U933_in[3] = arr__U926_out[3];
assign arr__U933_in[2] = arr__U926_out[2];
assign arr__U933_in[1] = arr__U926_out[1];
assign arr__U933_in[0] = arr__U926_out[0];
array_delay_U934 arr__U933 (
    .clk(clk),
    .in(arr__U933_in),
    .out(arr__U933_out)
);
wire [15:0] arr__U940_in [4:0];
assign arr__U940_in[4] = arr__U933_out[4];
assign arr__U940_in[3] = arr__U933_out[3];
assign arr__U940_in[2] = arr__U933_out[2];
assign arr__U940_in[1] = arr__U933_out[1];
assign arr__U940_in[0] = arr__U933_out[0];
array_delay_U941 arr__U940 (
    .clk(clk),
    .in(arr__U940_in),
    .out(arr__U940_out)
);
wire [15:0] arr__U947_in [4:0];
assign arr__U947_in[4] = arr__U940_out[4];
assign arr__U947_in[3] = arr__U940_out[3];
assign arr__U947_in[2] = arr__U940_out[2];
assign arr__U947_in[1] = arr__U940_out[1];
assign arr__U947_in[0] = arr__U940_out[0];
array_delay_U948 arr__U947 (
    .clk(clk),
    .in(arr__U947_in),
    .out(arr__U947_out)
);
wire [15:0] arr__U954_in [4:0];
assign arr__U954_in[4] = arr__U947_out[4];
assign arr__U954_in[3] = arr__U947_out[3];
assign arr__U954_in[2] = arr__U947_out[2];
assign arr__U954_in[1] = arr__U947_out[1];
assign arr__U954_in[0] = arr__U947_out[0];
array_delay_U955 arr__U954 (
    .clk(clk),
    .in(arr__U954_in),
    .out(arr__U954_out)
);
wire [15:0] arr__U961_in [4:0];
assign arr__U961_in[4] = arr__U954_out[4];
assign arr__U961_in[3] = arr__U954_out[3];
assign arr__U961_in[2] = arr__U954_out[2];
assign arr__U961_in[1] = arr__U954_out[1];
assign arr__U961_in[0] = arr__U954_out[0];
array_delay_U962 arr__U961 (
    .clk(clk),
    .in(arr__U961_in),
    .out(arr__U961_out)
);
wire [15:0] conv_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[4] = op_hcompute_conv_stencil_10_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[3] = op_hcompute_conv_stencil_10_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[2] = op_hcompute_conv_stencil_10_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[1] = op_hcompute_conv_stencil_10_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[0] = op_hcompute_conv_stencil_10_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_10_write_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_10_write_ctrl_vars[4] = op_hcompute_conv_stencil_10_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_10_write_ctrl_vars[3] = op_hcompute_conv_stencil_10_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_10_write_ctrl_vars[2] = op_hcompute_conv_stencil_10_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_10_write_ctrl_vars[1] = op_hcompute_conv_stencil_10_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_10_write_ctrl_vars[0] = op_hcompute_conv_stencil_10_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_10_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_10_write[0] = op_hcompute_conv_stencil_10_conv_stencil_op_hcompute_conv_stencil_10_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[4] = op_hcompute_conv_stencil_11_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[3] = op_hcompute_conv_stencil_11_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[2] = op_hcompute_conv_stencil_11_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[1] = op_hcompute_conv_stencil_11_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[0] = op_hcompute_conv_stencil_11_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_11_write_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_11_write_ctrl_vars[4] = op_hcompute_conv_stencil_11_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_11_write_ctrl_vars[3] = op_hcompute_conv_stencil_11_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_11_write_ctrl_vars[2] = op_hcompute_conv_stencil_11_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_11_write_ctrl_vars[1] = op_hcompute_conv_stencil_11_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_11_write_ctrl_vars[0] = op_hcompute_conv_stencil_11_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_11_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_11_write[0] = op_hcompute_conv_stencil_11_conv_stencil_op_hcompute_conv_stencil_11_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[4] = op_hcompute_conv_stencil_12_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[3] = op_hcompute_conv_stencil_12_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[2] = op_hcompute_conv_stencil_12_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[1] = op_hcompute_conv_stencil_12_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[0] = op_hcompute_conv_stencil_12_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_12_write_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_12_write_ctrl_vars[4] = op_hcompute_conv_stencil_12_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_12_write_ctrl_vars[3] = op_hcompute_conv_stencil_12_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_12_write_ctrl_vars[2] = op_hcompute_conv_stencil_12_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_12_write_ctrl_vars[1] = op_hcompute_conv_stencil_12_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_12_write_ctrl_vars[0] = op_hcompute_conv_stencil_12_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_12_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_12_write[0] = op_hcompute_conv_stencil_12_conv_stencil_op_hcompute_conv_stencil_12_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[4] = op_hcompute_conv_stencil_13_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[3] = op_hcompute_conv_stencil_13_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[2] = op_hcompute_conv_stencil_13_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[1] = op_hcompute_conv_stencil_13_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[0] = op_hcompute_conv_stencil_13_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_13_write_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_13_write_ctrl_vars[4] = op_hcompute_conv_stencil_13_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_13_write_ctrl_vars[3] = op_hcompute_conv_stencil_13_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_13_write_ctrl_vars[2] = op_hcompute_conv_stencil_13_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_13_write_ctrl_vars[1] = op_hcompute_conv_stencil_13_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_13_write_ctrl_vars[0] = op_hcompute_conv_stencil_13_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_13_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_13_write[0] = op_hcompute_conv_stencil_13_conv_stencil_op_hcompute_conv_stencil_13_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[4] = op_hcompute_conv_stencil_14_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[3] = op_hcompute_conv_stencil_14_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[2] = op_hcompute_conv_stencil_14_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[1] = op_hcompute_conv_stencil_14_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[0] = op_hcompute_conv_stencil_14_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_14_write_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_14_write_ctrl_vars[4] = op_hcompute_conv_stencil_14_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_14_write_ctrl_vars[3] = op_hcompute_conv_stencil_14_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_14_write_ctrl_vars[2] = op_hcompute_conv_stencil_14_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_14_write_ctrl_vars[1] = op_hcompute_conv_stencil_14_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_14_write_ctrl_vars[0] = op_hcompute_conv_stencil_14_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_14_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_14_write[0] = op_hcompute_conv_stencil_14_conv_stencil_op_hcompute_conv_stencil_14_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[4] = op_hcompute_conv_stencil_15_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[3] = op_hcompute_conv_stencil_15_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[2] = op_hcompute_conv_stencil_15_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[1] = op_hcompute_conv_stencil_15_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[0] = op_hcompute_conv_stencil_15_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_15_write_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_15_write_ctrl_vars[4] = op_hcompute_conv_stencil_15_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_15_write_ctrl_vars[3] = op_hcompute_conv_stencil_15_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_15_write_ctrl_vars[2] = op_hcompute_conv_stencil_15_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_15_write_ctrl_vars[1] = op_hcompute_conv_stencil_15_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_15_write_ctrl_vars[0] = op_hcompute_conv_stencil_15_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_15_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_15_write[0] = op_hcompute_conv_stencil_15_conv_stencil_op_hcompute_conv_stencil_15_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[2] = op_hcompute_conv_stencil_1_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[1] = op_hcompute_conv_stencil_1_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[0] = op_hcompute_conv_stencil_1_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[2] = op_hcompute_conv_stencil_2_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[1] = op_hcompute_conv_stencil_2_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[0] = op_hcompute_conv_stencil_2_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[2] = op_hcompute_conv_stencil_3_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[1] = op_hcompute_conv_stencil_3_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[0] = op_hcompute_conv_stencil_3_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[2] = op_hcompute_conv_stencil_4_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[1] = op_hcompute_conv_stencil_4_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[0] = op_hcompute_conv_stencil_4_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[2] = op_hcompute_conv_stencil_5_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[1] = op_hcompute_conv_stencil_5_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[0] = op_hcompute_conv_stencil_5_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_6_write_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_conv_stencil_6_write_ctrl_vars[2] = op_hcompute_conv_stencil_6_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_6_write_ctrl_vars[1] = op_hcompute_conv_stencil_6_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_6_write_ctrl_vars[0] = op_hcompute_conv_stencil_6_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_6_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_6_write[0] = op_hcompute_conv_stencil_6_conv_stencil_op_hcompute_conv_stencil_6_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_7_write_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_conv_stencil_7_write_ctrl_vars[2] = op_hcompute_conv_stencil_7_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_7_write_ctrl_vars[1] = op_hcompute_conv_stencil_7_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_7_write_ctrl_vars[0] = op_hcompute_conv_stencil_7_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_7_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_7_write[0] = op_hcompute_conv_stencil_7_conv_stencil_op_hcompute_conv_stencil_7_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[4] = op_hcompute_conv_stencil_8_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[3] = op_hcompute_conv_stencil_8_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[2] = op_hcompute_conv_stencil_8_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[1] = op_hcompute_conv_stencil_8_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[0] = op_hcompute_conv_stencil_8_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_8_write_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_8_write_ctrl_vars[4] = op_hcompute_conv_stencil_8_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_8_write_ctrl_vars[3] = op_hcompute_conv_stencil_8_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_8_write_ctrl_vars[2] = op_hcompute_conv_stencil_8_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_8_write_ctrl_vars[1] = op_hcompute_conv_stencil_8_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_8_write_ctrl_vars[0] = op_hcompute_conv_stencil_8_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_8_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_8_write[0] = op_hcompute_conv_stencil_8_conv_stencil_op_hcompute_conv_stencil_8_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[4] = op_hcompute_conv_stencil_9_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[3] = op_hcompute_conv_stencil_9_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[2] = op_hcompute_conv_stencil_9_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[1] = op_hcompute_conv_stencil_9_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[0] = op_hcompute_conv_stencil_9_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_9_write_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_9_write_ctrl_vars[4] = op_hcompute_conv_stencil_9_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_9_write_ctrl_vars[3] = op_hcompute_conv_stencil_9_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_9_write_ctrl_vars[2] = op_hcompute_conv_stencil_9_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_9_write_ctrl_vars[1] = op_hcompute_conv_stencil_9_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_9_write_ctrl_vars[0] = op_hcompute_conv_stencil_9_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_9_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_9_write[0] = op_hcompute_conv_stencil_9_conv_stencil_op_hcompute_conv_stencil_9_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[2] = op_hcompute_conv_stencil_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[1] = op_hcompute_conv_stencil_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[0] = op_hcompute_conv_stencil_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_write[0] = op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write[0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_1_read_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_hw_output_stencil_1_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_1_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_1_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_1_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_1_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_1_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_2_read_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_hw_output_stencil_2_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_2_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_2_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_2_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_2_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_2_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_3_read_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_hw_output_stencil_3_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_3_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_3_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_3_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_3_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_3_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_4_read_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_hw_output_stencil_4_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_4_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_4_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_4_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_4_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_4_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_5_read_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_hw_output_stencil_5_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_5_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_5_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_5_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_5_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_5_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_6_read_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_hw_output_stencil_6_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_6_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_6_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_6_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_6_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_6_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_7_read_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_hw_output_stencil_7_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_7_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_7_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_7_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_7_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_7_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
conv_stencil_ub conv_stencil (
    .clk(clk),
    .flush(flush),
    .rst_n(rst_n),
    .op_hcompute_conv_stencil_10_read_ren(op_hcompute_conv_stencil_10_read_start_out),
    .op_hcompute_conv_stencil_10_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars),
    .op_hcompute_conv_stencil_10_read(conv_stencil_op_hcompute_conv_stencil_10_read),
    .op_hcompute_conv_stencil_10_write_wen(op_hcompute_conv_stencil_10_write_start_out),
    .op_hcompute_conv_stencil_10_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_10_write_ctrl_vars),
    .op_hcompute_conv_stencil_10_write(conv_stencil_op_hcompute_conv_stencil_10_write),
    .op_hcompute_conv_stencil_11_read_ren(op_hcompute_conv_stencil_11_read_start_out),
    .op_hcompute_conv_stencil_11_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars),
    .op_hcompute_conv_stencil_11_read(conv_stencil_op_hcompute_conv_stencil_11_read),
    .op_hcompute_conv_stencil_11_write_wen(op_hcompute_conv_stencil_11_write_start_out),
    .op_hcompute_conv_stencil_11_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_11_write_ctrl_vars),
    .op_hcompute_conv_stencil_11_write(conv_stencil_op_hcompute_conv_stencil_11_write),
    .op_hcompute_conv_stencil_12_read_ren(op_hcompute_conv_stencil_12_read_start_out),
    .op_hcompute_conv_stencil_12_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars),
    .op_hcompute_conv_stencil_12_read(conv_stencil_op_hcompute_conv_stencil_12_read),
    .op_hcompute_conv_stencil_12_write_wen(op_hcompute_conv_stencil_12_write_start_out),
    .op_hcompute_conv_stencil_12_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_12_write_ctrl_vars),
    .op_hcompute_conv_stencil_12_write(conv_stencil_op_hcompute_conv_stencil_12_write),
    .op_hcompute_conv_stencil_13_read_ren(op_hcompute_conv_stencil_13_read_start_out),
    .op_hcompute_conv_stencil_13_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars),
    .op_hcompute_conv_stencil_13_read(conv_stencil_op_hcompute_conv_stencil_13_read),
    .op_hcompute_conv_stencil_13_write_wen(op_hcompute_conv_stencil_13_write_start_out),
    .op_hcompute_conv_stencil_13_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_13_write_ctrl_vars),
    .op_hcompute_conv_stencil_13_write(conv_stencil_op_hcompute_conv_stencil_13_write),
    .op_hcompute_conv_stencil_14_read_ren(op_hcompute_conv_stencil_14_read_start_out),
    .op_hcompute_conv_stencil_14_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars),
    .op_hcompute_conv_stencil_14_read(conv_stencil_op_hcompute_conv_stencil_14_read),
    .op_hcompute_conv_stencil_14_write_wen(op_hcompute_conv_stencil_14_write_start_out),
    .op_hcompute_conv_stencil_14_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_14_write_ctrl_vars),
    .op_hcompute_conv_stencil_14_write(conv_stencil_op_hcompute_conv_stencil_14_write),
    .op_hcompute_conv_stencil_15_read_ren(op_hcompute_conv_stencil_15_read_start_out),
    .op_hcompute_conv_stencil_15_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars),
    .op_hcompute_conv_stencil_15_read(conv_stencil_op_hcompute_conv_stencil_15_read),
    .op_hcompute_conv_stencil_15_write_wen(op_hcompute_conv_stencil_15_write_start_out),
    .op_hcompute_conv_stencil_15_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_15_write_ctrl_vars),
    .op_hcompute_conv_stencil_15_write(conv_stencil_op_hcompute_conv_stencil_15_write),
    .op_hcompute_conv_stencil_1_write_wen(op_hcompute_conv_stencil_1_write_start_out),
    .op_hcompute_conv_stencil_1_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars),
    .op_hcompute_conv_stencil_1_write(conv_stencil_op_hcompute_conv_stencil_1_write),
    .op_hcompute_conv_stencil_2_write_wen(op_hcompute_conv_stencil_2_write_start_out),
    .op_hcompute_conv_stencil_2_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars),
    .op_hcompute_conv_stencil_2_write(conv_stencil_op_hcompute_conv_stencil_2_write),
    .op_hcompute_conv_stencil_3_write_wen(op_hcompute_conv_stencil_3_write_start_out),
    .op_hcompute_conv_stencil_3_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars),
    .op_hcompute_conv_stencil_3_write(conv_stencil_op_hcompute_conv_stencil_3_write),
    .op_hcompute_conv_stencil_4_write_wen(op_hcompute_conv_stencil_4_write_start_out),
    .op_hcompute_conv_stencil_4_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars),
    .op_hcompute_conv_stencil_4_write(conv_stencil_op_hcompute_conv_stencil_4_write),
    .op_hcompute_conv_stencil_5_write_wen(op_hcompute_conv_stencil_5_write_start_out),
    .op_hcompute_conv_stencil_5_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars),
    .op_hcompute_conv_stencil_5_write(conv_stencil_op_hcompute_conv_stencil_5_write),
    .op_hcompute_conv_stencil_6_write_wen(op_hcompute_conv_stencil_6_write_start_out),
    .op_hcompute_conv_stencil_6_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_6_write_ctrl_vars),
    .op_hcompute_conv_stencil_6_write(conv_stencil_op_hcompute_conv_stencil_6_write),
    .op_hcompute_conv_stencil_7_write_wen(op_hcompute_conv_stencil_7_write_start_out),
    .op_hcompute_conv_stencil_7_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_7_write_ctrl_vars),
    .op_hcompute_conv_stencil_7_write(conv_stencil_op_hcompute_conv_stencil_7_write),
    .op_hcompute_conv_stencil_8_read_ren(op_hcompute_conv_stencil_8_read_start_out),
    .op_hcompute_conv_stencil_8_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars),
    .op_hcompute_conv_stencil_8_read(conv_stencil_op_hcompute_conv_stencil_8_read),
    .op_hcompute_conv_stencil_8_write_wen(op_hcompute_conv_stencil_8_write_start_out),
    .op_hcompute_conv_stencil_8_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_8_write_ctrl_vars),
    .op_hcompute_conv_stencil_8_write(conv_stencil_op_hcompute_conv_stencil_8_write),
    .op_hcompute_conv_stencil_9_read_ren(op_hcompute_conv_stencil_9_read_start_out),
    .op_hcompute_conv_stencil_9_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars),
    .op_hcompute_conv_stencil_9_read(conv_stencil_op_hcompute_conv_stencil_9_read),
    .op_hcompute_conv_stencil_9_write_wen(op_hcompute_conv_stencil_9_write_start_out),
    .op_hcompute_conv_stencil_9_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_9_write_ctrl_vars),
    .op_hcompute_conv_stencil_9_write(conv_stencil_op_hcompute_conv_stencil_9_write),
    .op_hcompute_conv_stencil_write_wen(op_hcompute_conv_stencil_write_start_out),
    .op_hcompute_conv_stencil_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars),
    .op_hcompute_conv_stencil_write(conv_stencil_op_hcompute_conv_stencil_write),
    .op_hcompute_hw_output_stencil_1_read_ren(op_hcompute_hw_output_stencil_1_read_start_out),
    .op_hcompute_hw_output_stencil_1_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_1_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_1_read(conv_stencil_op_hcompute_hw_output_stencil_1_read),
    .op_hcompute_hw_output_stencil_2_read_ren(op_hcompute_hw_output_stencil_2_read_start_out),
    .op_hcompute_hw_output_stencil_2_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_2_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_2_read(conv_stencil_op_hcompute_hw_output_stencil_2_read),
    .op_hcompute_hw_output_stencil_3_read_ren(op_hcompute_hw_output_stencil_3_read_start_out),
    .op_hcompute_hw_output_stencil_3_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_3_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_3_read(conv_stencil_op_hcompute_hw_output_stencil_3_read),
    .op_hcompute_hw_output_stencil_4_read_ren(op_hcompute_hw_output_stencil_4_read_start_out),
    .op_hcompute_hw_output_stencil_4_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_4_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_4_read(conv_stencil_op_hcompute_hw_output_stencil_4_read),
    .op_hcompute_hw_output_stencil_5_read_ren(op_hcompute_hw_output_stencil_5_read_start_out),
    .op_hcompute_hw_output_stencil_5_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_5_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_5_read(conv_stencil_op_hcompute_hw_output_stencil_5_read),
    .op_hcompute_hw_output_stencil_6_read_ren(op_hcompute_hw_output_stencil_6_read_start_out),
    .op_hcompute_hw_output_stencil_6_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_6_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_6_read(conv_stencil_op_hcompute_hw_output_stencil_6_read),
    .op_hcompute_hw_output_stencil_7_read_ren(op_hcompute_hw_output_stencil_7_read_start_out),
    .op_hcompute_hw_output_stencil_7_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_7_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_7_read(conv_stencil_op_hcompute_hw_output_stencil_7_read),
    .op_hcompute_hw_output_stencil_read_ren(op_hcompute_hw_output_stencil_read_start_out),
    .op_hcompute_hw_output_stencil_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_read(conv_stencil_op_hcompute_hw_output_stencil_read)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1001 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_11_port_controller_valid),
    .out(delay_reg__U1001_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1002 (
    .clk(clk),
    .in(delay_reg__U1001_out),
    .out(delay_reg__U1002_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1019 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_11_port_controller_valid),
    .out(delay_reg__U1019_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1020 (
    .clk(clk),
    .in(delay_reg__U1019_out),
    .out(delay_reg__U1020_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1021 (
    .clk(clk),
    .in(delay_reg__U1020_out),
    .out(delay_reg__U1021_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1022 (
    .clk(clk),
    .in(delay_reg__U1021_out),
    .out(delay_reg__U1022_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1023 (
    .clk(clk),
    .in(delay_reg__U1022_out),
    .out(delay_reg__U1023_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1024 (
    .clk(clk),
    .in(delay_reg__U1023_out),
    .out(delay_reg__U1024_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1025 (
    .clk(clk),
    .in(delay_reg__U1024_out),
    .out(delay_reg__U1025_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1026 (
    .clk(clk),
    .in(delay_reg__U1025_out),
    .out(delay_reg__U1026_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1027 (
    .clk(clk),
    .in(delay_reg__U1026_out),
    .out(delay_reg__U1027_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1028 (
    .clk(clk),
    .in(delay_reg__U1027_out),
    .out(delay_reg__U1028_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1029 (
    .clk(clk),
    .in(delay_reg__U1028_out),
    .out(delay_reg__U1029_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1030 (
    .clk(clk),
    .in(delay_reg__U1029_out),
    .out(delay_reg__U1030_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1031 (
    .clk(clk),
    .in(delay_reg__U1030_out),
    .out(delay_reg__U1031_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1032 (
    .clk(clk),
    .in(delay_reg__U1031_out),
    .out(delay_reg__U1032_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1033 (
    .clk(clk),
    .in(delay_reg__U1032_out),
    .out(delay_reg__U1033_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1034 (
    .clk(clk),
    .in(delay_reg__U1033_out),
    .out(delay_reg__U1034_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1035 (
    .clk(clk),
    .in(delay_reg__U1034_out),
    .out(delay_reg__U1035_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1189 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_12_port_controller_valid),
    .out(delay_reg__U1189_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1190 (
    .clk(clk),
    .in(delay_reg__U1189_out),
    .out(delay_reg__U1190_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1207 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_12_port_controller_valid),
    .out(delay_reg__U1207_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1208 (
    .clk(clk),
    .in(delay_reg__U1207_out),
    .out(delay_reg__U1208_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1209 (
    .clk(clk),
    .in(delay_reg__U1208_out),
    .out(delay_reg__U1209_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1210 (
    .clk(clk),
    .in(delay_reg__U1209_out),
    .out(delay_reg__U1210_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1211 (
    .clk(clk),
    .in(delay_reg__U1210_out),
    .out(delay_reg__U1211_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1212 (
    .clk(clk),
    .in(delay_reg__U1211_out),
    .out(delay_reg__U1212_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1213 (
    .clk(clk),
    .in(delay_reg__U1212_out),
    .out(delay_reg__U1213_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1214 (
    .clk(clk),
    .in(delay_reg__U1213_out),
    .out(delay_reg__U1214_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1215 (
    .clk(clk),
    .in(delay_reg__U1214_out),
    .out(delay_reg__U1215_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1216 (
    .clk(clk),
    .in(delay_reg__U1215_out),
    .out(delay_reg__U1216_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1217 (
    .clk(clk),
    .in(delay_reg__U1216_out),
    .out(delay_reg__U1217_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1218 (
    .clk(clk),
    .in(delay_reg__U1217_out),
    .out(delay_reg__U1218_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1219 (
    .clk(clk),
    .in(delay_reg__U1218_out),
    .out(delay_reg__U1219_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1220 (
    .clk(clk),
    .in(delay_reg__U1219_out),
    .out(delay_reg__U1220_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1221 (
    .clk(clk),
    .in(delay_reg__U1220_out),
    .out(delay_reg__U1221_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1222 (
    .clk(clk),
    .in(delay_reg__U1221_out),
    .out(delay_reg__U1222_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1223 (
    .clk(clk),
    .in(delay_reg__U1222_out),
    .out(delay_reg__U1223_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1377 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_13_port_controller_valid),
    .out(delay_reg__U1377_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1378 (
    .clk(clk),
    .in(delay_reg__U1377_out),
    .out(delay_reg__U1378_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1395 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_13_port_controller_valid),
    .out(delay_reg__U1395_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1396 (
    .clk(clk),
    .in(delay_reg__U1395_out),
    .out(delay_reg__U1396_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1397 (
    .clk(clk),
    .in(delay_reg__U1396_out),
    .out(delay_reg__U1397_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1398 (
    .clk(clk),
    .in(delay_reg__U1397_out),
    .out(delay_reg__U1398_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1399 (
    .clk(clk),
    .in(delay_reg__U1398_out),
    .out(delay_reg__U1399_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1400 (
    .clk(clk),
    .in(delay_reg__U1399_out),
    .out(delay_reg__U1400_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1401 (
    .clk(clk),
    .in(delay_reg__U1400_out),
    .out(delay_reg__U1401_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1402 (
    .clk(clk),
    .in(delay_reg__U1401_out),
    .out(delay_reg__U1402_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1403 (
    .clk(clk),
    .in(delay_reg__U1402_out),
    .out(delay_reg__U1403_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1404 (
    .clk(clk),
    .in(delay_reg__U1403_out),
    .out(delay_reg__U1404_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1405 (
    .clk(clk),
    .in(delay_reg__U1404_out),
    .out(delay_reg__U1405_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1406 (
    .clk(clk),
    .in(delay_reg__U1405_out),
    .out(delay_reg__U1406_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1407 (
    .clk(clk),
    .in(delay_reg__U1406_out),
    .out(delay_reg__U1407_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1408 (
    .clk(clk),
    .in(delay_reg__U1407_out),
    .out(delay_reg__U1408_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1409 (
    .clk(clk),
    .in(delay_reg__U1408_out),
    .out(delay_reg__U1409_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1410 (
    .clk(clk),
    .in(delay_reg__U1409_out),
    .out(delay_reg__U1410_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1411 (
    .clk(clk),
    .in(delay_reg__U1410_out),
    .out(delay_reg__U1411_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1565 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_14_port_controller_valid),
    .out(delay_reg__U1565_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1566 (
    .clk(clk),
    .in(delay_reg__U1565_out),
    .out(delay_reg__U1566_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1583 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_14_port_controller_valid),
    .out(delay_reg__U1583_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1584 (
    .clk(clk),
    .in(delay_reg__U1583_out),
    .out(delay_reg__U1584_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1585 (
    .clk(clk),
    .in(delay_reg__U1584_out),
    .out(delay_reg__U1585_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1586 (
    .clk(clk),
    .in(delay_reg__U1585_out),
    .out(delay_reg__U1586_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1587 (
    .clk(clk),
    .in(delay_reg__U1586_out),
    .out(delay_reg__U1587_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1588 (
    .clk(clk),
    .in(delay_reg__U1587_out),
    .out(delay_reg__U1588_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1589 (
    .clk(clk),
    .in(delay_reg__U1588_out),
    .out(delay_reg__U1589_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1590 (
    .clk(clk),
    .in(delay_reg__U1589_out),
    .out(delay_reg__U1590_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1591 (
    .clk(clk),
    .in(delay_reg__U1590_out),
    .out(delay_reg__U1591_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1592 (
    .clk(clk),
    .in(delay_reg__U1591_out),
    .out(delay_reg__U1592_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1593 (
    .clk(clk),
    .in(delay_reg__U1592_out),
    .out(delay_reg__U1593_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1594 (
    .clk(clk),
    .in(delay_reg__U1593_out),
    .out(delay_reg__U1594_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1595 (
    .clk(clk),
    .in(delay_reg__U1594_out),
    .out(delay_reg__U1595_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1596 (
    .clk(clk),
    .in(delay_reg__U1595_out),
    .out(delay_reg__U1596_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1597 (
    .clk(clk),
    .in(delay_reg__U1596_out),
    .out(delay_reg__U1597_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1598 (
    .clk(clk),
    .in(delay_reg__U1597_out),
    .out(delay_reg__U1598_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1599 (
    .clk(clk),
    .in(delay_reg__U1598_out),
    .out(delay_reg__U1599_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1753 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_15_port_controller_valid),
    .out(delay_reg__U1753_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1754 (
    .clk(clk),
    .in(delay_reg__U1753_out),
    .out(delay_reg__U1754_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1771 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_15_port_controller_valid),
    .out(delay_reg__U1771_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1772 (
    .clk(clk),
    .in(delay_reg__U1771_out),
    .out(delay_reg__U1772_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1773 (
    .clk(clk),
    .in(delay_reg__U1772_out),
    .out(delay_reg__U1773_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1774 (
    .clk(clk),
    .in(delay_reg__U1773_out),
    .out(delay_reg__U1774_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1775 (
    .clk(clk),
    .in(delay_reg__U1774_out),
    .out(delay_reg__U1775_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1776 (
    .clk(clk),
    .in(delay_reg__U1775_out),
    .out(delay_reg__U1776_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1777 (
    .clk(clk),
    .in(delay_reg__U1776_out),
    .out(delay_reg__U1777_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1778 (
    .clk(clk),
    .in(delay_reg__U1777_out),
    .out(delay_reg__U1778_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1779 (
    .clk(clk),
    .in(delay_reg__U1778_out),
    .out(delay_reg__U1779_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1780 (
    .clk(clk),
    .in(delay_reg__U1779_out),
    .out(delay_reg__U1780_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1781 (
    .clk(clk),
    .in(delay_reg__U1780_out),
    .out(delay_reg__U1781_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1782 (
    .clk(clk),
    .in(delay_reg__U1781_out),
    .out(delay_reg__U1782_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1783 (
    .clk(clk),
    .in(delay_reg__U1782_out),
    .out(delay_reg__U1783_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1784 (
    .clk(clk),
    .in(delay_reg__U1783_out),
    .out(delay_reg__U1784_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1785 (
    .clk(clk),
    .in(delay_reg__U1784_out),
    .out(delay_reg__U1785_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1786 (
    .clk(clk),
    .in(delay_reg__U1785_out),
    .out(delay_reg__U1786_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1787 (
    .clk(clk),
    .in(delay_reg__U1786_out),
    .out(delay_reg__U1787_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1928 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_port_controller_valid),
    .out(delay_reg__U1928_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1929 (
    .clk(clk),
    .in(delay_reg__U1928_out),
    .out(delay_reg__U1929_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1942 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_port_controller_valid),
    .out(delay_reg__U1942_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1943 (
    .clk(clk),
    .in(delay_reg__U1942_out),
    .out(delay_reg__U1943_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1975 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_1_port_controller_valid),
    .out(delay_reg__U1975_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1976 (
    .clk(clk),
    .in(delay_reg__U1975_out),
    .out(delay_reg__U1976_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1989 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_1_port_controller_valid),
    .out(delay_reg__U1989_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1990 (
    .clk(clk),
    .in(delay_reg__U1989_out),
    .out(delay_reg__U1990_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2022 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_2_port_controller_valid),
    .out(delay_reg__U2022_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2023 (
    .clk(clk),
    .in(delay_reg__U2022_out),
    .out(delay_reg__U2023_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2036 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_2_port_controller_valid),
    .out(delay_reg__U2036_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2037 (
    .clk(clk),
    .in(delay_reg__U2036_out),
    .out(delay_reg__U2037_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2069 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_3_port_controller_valid),
    .out(delay_reg__U2069_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2070 (
    .clk(clk),
    .in(delay_reg__U2069_out),
    .out(delay_reg__U2070_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2083 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_3_port_controller_valid),
    .out(delay_reg__U2083_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2084 (
    .clk(clk),
    .in(delay_reg__U2083_out),
    .out(delay_reg__U2084_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2116 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_4_port_controller_valid),
    .out(delay_reg__U2116_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2117 (
    .clk(clk),
    .in(delay_reg__U2116_out),
    .out(delay_reg__U2117_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2130 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_4_port_controller_valid),
    .out(delay_reg__U2130_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2131 (
    .clk(clk),
    .in(delay_reg__U2130_out),
    .out(delay_reg__U2131_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2163 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_5_port_controller_valid),
    .out(delay_reg__U2163_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2164 (
    .clk(clk),
    .in(delay_reg__U2163_out),
    .out(delay_reg__U2164_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2177 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_5_port_controller_valid),
    .out(delay_reg__U2177_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2178 (
    .clk(clk),
    .in(delay_reg__U2177_out),
    .out(delay_reg__U2178_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2210 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_6_port_controller_valid),
    .out(delay_reg__U2210_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2211 (
    .clk(clk),
    .in(delay_reg__U2210_out),
    .out(delay_reg__U2211_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2224 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_6_port_controller_valid),
    .out(delay_reg__U2224_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2225 (
    .clk(clk),
    .in(delay_reg__U2224_out),
    .out(delay_reg__U2225_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2257 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_7_port_controller_valid),
    .out(delay_reg__U2257_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2258 (
    .clk(clk),
    .in(delay_reg__U2257_out),
    .out(delay_reg__U2258_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2271 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_7_port_controller_valid),
    .out(delay_reg__U2271_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2272 (
    .clk(clk),
    .in(delay_reg__U2271_out),
    .out(delay_reg__U2272_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U437 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_8_port_controller_valid),
    .out(delay_reg__U437_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U438 (
    .clk(clk),
    .in(delay_reg__U437_out),
    .out(delay_reg__U438_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U455 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_8_port_controller_valid),
    .out(delay_reg__U455_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U456 (
    .clk(clk),
    .in(delay_reg__U455_out),
    .out(delay_reg__U456_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U457 (
    .clk(clk),
    .in(delay_reg__U456_out),
    .out(delay_reg__U457_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U458 (
    .clk(clk),
    .in(delay_reg__U457_out),
    .out(delay_reg__U458_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U459 (
    .clk(clk),
    .in(delay_reg__U458_out),
    .out(delay_reg__U459_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U460 (
    .clk(clk),
    .in(delay_reg__U459_out),
    .out(delay_reg__U460_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U461 (
    .clk(clk),
    .in(delay_reg__U460_out),
    .out(delay_reg__U461_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U462 (
    .clk(clk),
    .in(delay_reg__U461_out),
    .out(delay_reg__U462_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U463 (
    .clk(clk),
    .in(delay_reg__U462_out),
    .out(delay_reg__U463_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U464 (
    .clk(clk),
    .in(delay_reg__U463_out),
    .out(delay_reg__U464_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U465 (
    .clk(clk),
    .in(delay_reg__U464_out),
    .out(delay_reg__U465_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U466 (
    .clk(clk),
    .in(delay_reg__U465_out),
    .out(delay_reg__U466_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U467 (
    .clk(clk),
    .in(delay_reg__U466_out),
    .out(delay_reg__U467_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U468 (
    .clk(clk),
    .in(delay_reg__U467_out),
    .out(delay_reg__U468_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U469 (
    .clk(clk),
    .in(delay_reg__U468_out),
    .out(delay_reg__U469_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U470 (
    .clk(clk),
    .in(delay_reg__U469_out),
    .out(delay_reg__U470_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U471 (
    .clk(clk),
    .in(delay_reg__U470_out),
    .out(delay_reg__U471_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U625 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_9_port_controller_valid),
    .out(delay_reg__U625_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U626 (
    .clk(clk),
    .in(delay_reg__U625_out),
    .out(delay_reg__U626_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U643 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_9_port_controller_valid),
    .out(delay_reg__U643_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U644 (
    .clk(clk),
    .in(delay_reg__U643_out),
    .out(delay_reg__U644_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U645 (
    .clk(clk),
    .in(delay_reg__U644_out),
    .out(delay_reg__U645_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U646 (
    .clk(clk),
    .in(delay_reg__U645_out),
    .out(delay_reg__U646_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U647 (
    .clk(clk),
    .in(delay_reg__U646_out),
    .out(delay_reg__U647_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U648 (
    .clk(clk),
    .in(delay_reg__U647_out),
    .out(delay_reg__U648_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U649 (
    .clk(clk),
    .in(delay_reg__U648_out),
    .out(delay_reg__U649_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U650 (
    .clk(clk),
    .in(delay_reg__U649_out),
    .out(delay_reg__U650_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U651 (
    .clk(clk),
    .in(delay_reg__U650_out),
    .out(delay_reg__U651_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U652 (
    .clk(clk),
    .in(delay_reg__U651_out),
    .out(delay_reg__U652_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U653 (
    .clk(clk),
    .in(delay_reg__U652_out),
    .out(delay_reg__U653_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U654 (
    .clk(clk),
    .in(delay_reg__U653_out),
    .out(delay_reg__U654_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U655 (
    .clk(clk),
    .in(delay_reg__U654_out),
    .out(delay_reg__U655_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U656 (
    .clk(clk),
    .in(delay_reg__U655_out),
    .out(delay_reg__U656_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U657 (
    .clk(clk),
    .in(delay_reg__U656_out),
    .out(delay_reg__U657_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U658 (
    .clk(clk),
    .in(delay_reg__U657_out),
    .out(delay_reg__U658_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U659 (
    .clk(clk),
    .in(delay_reg__U658_out),
    .out(delay_reg__U659_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U813 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_10_port_controller_valid),
    .out(delay_reg__U813_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U814 (
    .clk(clk),
    .in(delay_reg__U813_out),
    .out(delay_reg__U814_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U831 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_10_port_controller_valid),
    .out(delay_reg__U831_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U832 (
    .clk(clk),
    .in(delay_reg__U831_out),
    .out(delay_reg__U832_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U833 (
    .clk(clk),
    .in(delay_reg__U832_out),
    .out(delay_reg__U833_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U834 (
    .clk(clk),
    .in(delay_reg__U833_out),
    .out(delay_reg__U834_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U835 (
    .clk(clk),
    .in(delay_reg__U834_out),
    .out(delay_reg__U835_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U836 (
    .clk(clk),
    .in(delay_reg__U835_out),
    .out(delay_reg__U836_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U837 (
    .clk(clk),
    .in(delay_reg__U836_out),
    .out(delay_reg__U837_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U838 (
    .clk(clk),
    .in(delay_reg__U837_out),
    .out(delay_reg__U838_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U839 (
    .clk(clk),
    .in(delay_reg__U838_out),
    .out(delay_reg__U839_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U840 (
    .clk(clk),
    .in(delay_reg__U839_out),
    .out(delay_reg__U840_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U841 (
    .clk(clk),
    .in(delay_reg__U840_out),
    .out(delay_reg__U841_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U842 (
    .clk(clk),
    .in(delay_reg__U841_out),
    .out(delay_reg__U842_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U843 (
    .clk(clk),
    .in(delay_reg__U842_out),
    .out(delay_reg__U843_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U844 (
    .clk(clk),
    .in(delay_reg__U843_out),
    .out(delay_reg__U844_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U845 (
    .clk(clk),
    .in(delay_reg__U844_out),
    .out(delay_reg__U845_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U846 (
    .clk(clk),
    .in(delay_reg__U845_out),
    .out(delay_reg__U846_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U847 (
    .clk(clk),
    .in(delay_reg__U846_out),
    .out(delay_reg__U847_out)
);
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars [4:0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[4] = op_hcompute_conv_stencil_10_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[3] = op_hcompute_conv_stencil_10_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[2] = op_hcompute_conv_stencil_10_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[1] = op_hcompute_conv_stencil_10_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[0] = op_hcompute_conv_stencil_10_port_controller_d[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars [4:0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[4] = op_hcompute_conv_stencil_11_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[3] = op_hcompute_conv_stencil_11_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[2] = op_hcompute_conv_stencil_11_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[1] = op_hcompute_conv_stencil_11_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[0] = op_hcompute_conv_stencil_11_port_controller_d[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars [4:0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[4] = op_hcompute_conv_stencil_12_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[3] = op_hcompute_conv_stencil_12_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[2] = op_hcompute_conv_stencil_12_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[1] = op_hcompute_conv_stencil_12_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[0] = op_hcompute_conv_stencil_12_port_controller_d[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars [4:0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[4] = op_hcompute_conv_stencil_13_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[3] = op_hcompute_conv_stencil_13_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[2] = op_hcompute_conv_stencil_13_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[1] = op_hcompute_conv_stencil_13_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[0] = op_hcompute_conv_stencil_13_port_controller_d[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars [4:0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[4] = op_hcompute_conv_stencil_14_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[3] = op_hcompute_conv_stencil_14_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[2] = op_hcompute_conv_stencil_14_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[1] = op_hcompute_conv_stencil_14_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[0] = op_hcompute_conv_stencil_14_port_controller_d[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars [4:0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[4] = op_hcompute_conv_stencil_15_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[3] = op_hcompute_conv_stencil_15_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[2] = op_hcompute_conv_stencil_15_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[1] = op_hcompute_conv_stencil_15_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[0] = op_hcompute_conv_stencil_15_port_controller_d[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars [4:0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[4] = op_hcompute_conv_stencil_8_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[3] = op_hcompute_conv_stencil_8_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[2] = op_hcompute_conv_stencil_8_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[1] = op_hcompute_conv_stencil_8_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[0] = op_hcompute_conv_stencil_8_port_controller_d[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars [4:0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[4] = op_hcompute_conv_stencil_9_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[3] = op_hcompute_conv_stencil_9_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[2] = op_hcompute_conv_stencil_9_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[1] = op_hcompute_conv_stencil_9_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[0] = op_hcompute_conv_stencil_9_port_controller_d[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write_ctrl_vars [2:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_out[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write [0:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write[0] = op_hcompute_hw_input_global_wrapper_stencil_1_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write_ctrl_vars [2:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_out[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write [0:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write[0] = op_hcompute_hw_input_global_wrapper_stencil_2_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write_ctrl_vars [2:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_out[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write [0:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write[0] = op_hcompute_hw_input_global_wrapper_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write_ctrl_vars [2:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_out[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write [0:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write[0] = op_hcompute_hw_input_global_wrapper_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write_ctrl_vars [2:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_out[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write [0:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write[0] = op_hcompute_hw_input_global_wrapper_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write_ctrl_vars [2:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_out[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write [0:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write[0] = op_hcompute_hw_input_global_wrapper_stencil_6_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write_ctrl_vars [2:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_out[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write [0:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write[0] = op_hcompute_hw_input_global_wrapper_stencil_7_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars [2:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0];
hw_input_global_wrapper_stencil_ub hw_input_global_wrapper_stencil (
    .clk(clk),
    .flush(flush),
    .rst_n(rst_n),
    .op_hcompute_conv_stencil_10_read_ren(op_hcompute_conv_stencil_10_read_start_out),
    .op_hcompute_conv_stencil_10_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars),
    .op_hcompute_conv_stencil_10_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read),
    .op_hcompute_conv_stencil_11_read_ren(op_hcompute_conv_stencil_11_read_start_out),
    .op_hcompute_conv_stencil_11_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars),
    .op_hcompute_conv_stencil_11_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read),
    .op_hcompute_conv_stencil_12_read_ren(op_hcompute_conv_stencil_12_read_start_out),
    .op_hcompute_conv_stencil_12_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars),
    .op_hcompute_conv_stencil_12_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read),
    .op_hcompute_conv_stencil_13_read_ren(op_hcompute_conv_stencil_13_read_start_out),
    .op_hcompute_conv_stencil_13_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars),
    .op_hcompute_conv_stencil_13_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read),
    .op_hcompute_conv_stencil_14_read_ren(op_hcompute_conv_stencil_14_read_start_out),
    .op_hcompute_conv_stencil_14_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars),
    .op_hcompute_conv_stencil_14_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read),
    .op_hcompute_conv_stencil_15_read_ren(op_hcompute_conv_stencil_15_read_start_out),
    .op_hcompute_conv_stencil_15_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars),
    .op_hcompute_conv_stencil_15_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read),
    .op_hcompute_conv_stencil_8_read_ren(op_hcompute_conv_stencil_8_read_start_out),
    .op_hcompute_conv_stencil_8_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars),
    .op_hcompute_conv_stencil_8_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read),
    .op_hcompute_conv_stencil_9_read_ren(op_hcompute_conv_stencil_9_read_start_out),
    .op_hcompute_conv_stencil_9_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars),
    .op_hcompute_conv_stencil_9_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read),
    .op_hcompute_hw_input_global_wrapper_stencil_1_write_wen(op_hcompute_hw_input_global_wrapper_stencil_1_write_start_out),
    .op_hcompute_hw_input_global_wrapper_stencil_1_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_1_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write),
    .op_hcompute_hw_input_global_wrapper_stencil_2_write_wen(op_hcompute_hw_input_global_wrapper_stencil_2_write_start_out),
    .op_hcompute_hw_input_global_wrapper_stencil_2_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_2_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write),
    .op_hcompute_hw_input_global_wrapper_stencil_3_write_wen(op_hcompute_hw_input_global_wrapper_stencil_3_write_start_out),
    .op_hcompute_hw_input_global_wrapper_stencil_3_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_3_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write),
    .op_hcompute_hw_input_global_wrapper_stencil_4_write_wen(op_hcompute_hw_input_global_wrapper_stencil_4_write_start_out),
    .op_hcompute_hw_input_global_wrapper_stencil_4_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_4_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write),
    .op_hcompute_hw_input_global_wrapper_stencil_5_write_wen(op_hcompute_hw_input_global_wrapper_stencil_5_write_start_out),
    .op_hcompute_hw_input_global_wrapper_stencil_5_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_5_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write),
    .op_hcompute_hw_input_global_wrapper_stencil_6_write_wen(op_hcompute_hw_input_global_wrapper_stencil_6_write_start_out),
    .op_hcompute_hw_input_global_wrapper_stencil_6_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_6_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write),
    .op_hcompute_hw_input_global_wrapper_stencil_7_write_wen(op_hcompute_hw_input_global_wrapper_stencil_7_write_start_out),
    .op_hcompute_hw_input_global_wrapper_stencil_7_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_7_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write),
    .op_hcompute_hw_input_global_wrapper_stencil_write_wen(op_hcompute_hw_input_global_wrapper_stencil_write_start_out),
    .op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars [4:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[4] = op_hcompute_conv_stencil_10_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[3] = op_hcompute_conv_stencil_10_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[2] = op_hcompute_conv_stencil_10_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[1] = op_hcompute_conv_stencil_10_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[0] = op_hcompute_conv_stencil_10_port_controller_d[0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars [4:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[4] = op_hcompute_conv_stencil_11_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[3] = op_hcompute_conv_stencil_11_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[2] = op_hcompute_conv_stencil_11_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[1] = op_hcompute_conv_stencil_11_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[0] = op_hcompute_conv_stencil_11_port_controller_d[0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars [4:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[4] = op_hcompute_conv_stencil_12_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[3] = op_hcompute_conv_stencil_12_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[2] = op_hcompute_conv_stencil_12_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[1] = op_hcompute_conv_stencil_12_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[0] = op_hcompute_conv_stencil_12_port_controller_d[0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars [4:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[4] = op_hcompute_conv_stencil_13_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[3] = op_hcompute_conv_stencil_13_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[2] = op_hcompute_conv_stencil_13_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[1] = op_hcompute_conv_stencil_13_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[0] = op_hcompute_conv_stencil_13_port_controller_d[0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars [4:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[4] = op_hcompute_conv_stencil_14_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[3] = op_hcompute_conv_stencil_14_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[2] = op_hcompute_conv_stencil_14_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[1] = op_hcompute_conv_stencil_14_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[0] = op_hcompute_conv_stencil_14_port_controller_d[0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars [4:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[4] = op_hcompute_conv_stencil_15_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[3] = op_hcompute_conv_stencil_15_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[2] = op_hcompute_conv_stencil_15_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[1] = op_hcompute_conv_stencil_15_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[0] = op_hcompute_conv_stencil_15_port_controller_d[0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars [4:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[4] = op_hcompute_conv_stencil_8_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[3] = op_hcompute_conv_stencil_8_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[2] = op_hcompute_conv_stencil_8_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[1] = op_hcompute_conv_stencil_8_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[0] = op_hcompute_conv_stencil_8_port_controller_d[0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars [4:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[4] = op_hcompute_conv_stencil_9_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[3] = op_hcompute_conv_stencil_9_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[2] = op_hcompute_conv_stencil_9_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[1] = op_hcompute_conv_stencil_9_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[0] = op_hcompute_conv_stencil_9_port_controller_d[0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars [4:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[4] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0];
hw_kernel_global_wrapper_stencil_ub hw_kernel_global_wrapper_stencil (
    .clk(clk),
    .flush(flush),
    .rst_n(rst_n),
    .op_hcompute_conv_stencil_10_read_ren(op_hcompute_conv_stencil_10_read_start_out),
    .op_hcompute_conv_stencil_10_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars),
    .op_hcompute_conv_stencil_10_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read),
    .op_hcompute_conv_stencil_11_read_ren(op_hcompute_conv_stencil_11_read_start_out),
    .op_hcompute_conv_stencil_11_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars),
    .op_hcompute_conv_stencil_11_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read),
    .op_hcompute_conv_stencil_12_read_ren(op_hcompute_conv_stencil_12_read_start_out),
    .op_hcompute_conv_stencil_12_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars),
    .op_hcompute_conv_stencil_12_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read),
    .op_hcompute_conv_stencil_13_read_ren(op_hcompute_conv_stencil_13_read_start_out),
    .op_hcompute_conv_stencil_13_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars),
    .op_hcompute_conv_stencil_13_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read),
    .op_hcompute_conv_stencil_14_read_ren(op_hcompute_conv_stencil_14_read_start_out),
    .op_hcompute_conv_stencil_14_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars),
    .op_hcompute_conv_stencil_14_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read),
    .op_hcompute_conv_stencil_15_read_ren(op_hcompute_conv_stencil_15_read_start_out),
    .op_hcompute_conv_stencil_15_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars),
    .op_hcompute_conv_stencil_15_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read),
    .op_hcompute_conv_stencil_8_read_ren(op_hcompute_conv_stencil_8_read_start_out),
    .op_hcompute_conv_stencil_8_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars),
    .op_hcompute_conv_stencil_8_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read),
    .op_hcompute_conv_stencil_9_read_ren(op_hcompute_conv_stencil_9_read_start_out),
    .op_hcompute_conv_stencil_9_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars),
    .op_hcompute_conv_stencil_9_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_wen(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
cu_op_hcompute_conv_stencil op_hcompute_conv_stencil (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_write(op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write)
);
cu_op_hcompute_conv_stencil_1 op_hcompute_conv_stencil_1 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_1_write(op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write)
);
wire [15:0] op_hcompute_conv_stencil_10_conv_stencil_op_hcompute_conv_stencil_10_read [0:0];
assign op_hcompute_conv_stencil_10_conv_stencil_op_hcompute_conv_stencil_10_read[0] = conv_stencil_op_hcompute_conv_stencil_10_read[0];
wire [15:0] op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read [7:0];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[7];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[6];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[5];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[4];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[3];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[2];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[1];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[0];
wire [15:0] op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read [7:0];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[7];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[6];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[5];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[4];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[3];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[2];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[1];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[0];
cu_op_hcompute_conv_stencil_10 op_hcompute_conv_stencil_10 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_10_read(op_hcompute_conv_stencil_10_conv_stencil_op_hcompute_conv_stencil_10_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read(op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read(op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read),
    .conv_stencil_op_hcompute_conv_stencil_10_write(op_hcompute_conv_stencil_10_conv_stencil_op_hcompute_conv_stencil_10_write)
);
op_hcompute_conv_stencil_10_exe_start_pt__U812 op_hcompute_conv_stencil_10_exe_start (
    .in(delay_reg__U814_out),
    .out(op_hcompute_conv_stencil_10_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_10_exe_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_10_exe_start_control_vars_in[4] = arr__U823_out[4];
assign op_hcompute_conv_stencil_10_exe_start_control_vars_in[3] = arr__U823_out[3];
assign op_hcompute_conv_stencil_10_exe_start_control_vars_in[2] = arr__U823_out[2];
assign op_hcompute_conv_stencil_10_exe_start_control_vars_in[1] = arr__U823_out[1];
assign op_hcompute_conv_stencil_10_exe_start_control_vars_in[0] = arr__U823_out[0];
op_hcompute_conv_stencil_10_exe_start_control_vars_pt__U815 op_hcompute_conv_stencil_10_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_10_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_10_exe_start_control_vars_out)
);
affine_controller__U780 op_hcompute_conv_stencil_10_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_10_port_controller_valid),
    .d(op_hcompute_conv_stencil_10_port_controller_d)
);
op_hcompute_conv_stencil_10_read_start_pt__U810 op_hcompute_conv_stencil_10_read_start (
    .in(op_hcompute_conv_stencil_10_port_controller_valid),
    .out(op_hcompute_conv_stencil_10_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_10_read_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_10_read_start_control_vars_in[4] = op_hcompute_conv_stencil_10_port_controller_d[4];
assign op_hcompute_conv_stencil_10_read_start_control_vars_in[3] = op_hcompute_conv_stencil_10_port_controller_d[3];
assign op_hcompute_conv_stencil_10_read_start_control_vars_in[2] = op_hcompute_conv_stencil_10_port_controller_d[2];
assign op_hcompute_conv_stencil_10_read_start_control_vars_in[1] = op_hcompute_conv_stencil_10_port_controller_d[1];
assign op_hcompute_conv_stencil_10_read_start_control_vars_in[0] = op_hcompute_conv_stencil_10_port_controller_d[0];
op_hcompute_conv_stencil_10_read_start_control_vars_pt__U811 op_hcompute_conv_stencil_10_read_start_control_vars (
    .in(op_hcompute_conv_stencil_10_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_10_read_start_control_vars_out)
);
op_hcompute_conv_stencil_10_write_start_pt__U830 op_hcompute_conv_stencil_10_write_start (
    .in(delay_reg__U847_out),
    .out(op_hcompute_conv_stencil_10_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_10_write_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_10_write_start_control_vars_in[4] = arr__U961_out[4];
assign op_hcompute_conv_stencil_10_write_start_control_vars_in[3] = arr__U961_out[3];
assign op_hcompute_conv_stencil_10_write_start_control_vars_in[2] = arr__U961_out[2];
assign op_hcompute_conv_stencil_10_write_start_control_vars_in[1] = arr__U961_out[1];
assign op_hcompute_conv_stencil_10_write_start_control_vars_in[0] = arr__U961_out[0];
op_hcompute_conv_stencil_10_write_start_control_vars_pt__U848 op_hcompute_conv_stencil_10_write_start_control_vars (
    .in(op_hcompute_conv_stencil_10_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_10_write_start_control_vars_out)
);
wire [15:0] op_hcompute_conv_stencil_11_conv_stencil_op_hcompute_conv_stencil_11_read [0:0];
assign op_hcompute_conv_stencil_11_conv_stencil_op_hcompute_conv_stencil_11_read[0] = conv_stencil_op_hcompute_conv_stencil_11_read[0];
wire [15:0] op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read [7:0];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[7];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[6];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[5];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[4];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[3];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[2];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[1];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[0];
wire [15:0] op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read [7:0];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[7];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[6];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[5];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[4];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[3];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[2];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[1];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[0];
cu_op_hcompute_conv_stencil_11 op_hcompute_conv_stencil_11 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_11_read(op_hcompute_conv_stencil_11_conv_stencil_op_hcompute_conv_stencil_11_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read(op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read(op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read),
    .conv_stencil_op_hcompute_conv_stencil_11_write(op_hcompute_conv_stencil_11_conv_stencil_op_hcompute_conv_stencil_11_write)
);
op_hcompute_conv_stencil_11_exe_start_pt__U1000 op_hcompute_conv_stencil_11_exe_start (
    .in(delay_reg__U1002_out),
    .out(op_hcompute_conv_stencil_11_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_11_exe_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_11_exe_start_control_vars_in[4] = arr__U1011_out[4];
assign op_hcompute_conv_stencil_11_exe_start_control_vars_in[3] = arr__U1011_out[3];
assign op_hcompute_conv_stencil_11_exe_start_control_vars_in[2] = arr__U1011_out[2];
assign op_hcompute_conv_stencil_11_exe_start_control_vars_in[1] = arr__U1011_out[1];
assign op_hcompute_conv_stencil_11_exe_start_control_vars_in[0] = arr__U1011_out[0];
op_hcompute_conv_stencil_11_exe_start_control_vars_pt__U1003 op_hcompute_conv_stencil_11_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_11_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_11_exe_start_control_vars_out)
);
affine_controller__U968 op_hcompute_conv_stencil_11_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_11_port_controller_valid),
    .d(op_hcompute_conv_stencil_11_port_controller_d)
);
op_hcompute_conv_stencil_11_read_start_pt__U998 op_hcompute_conv_stencil_11_read_start (
    .in(op_hcompute_conv_stencil_11_port_controller_valid),
    .out(op_hcompute_conv_stencil_11_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_11_read_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_11_read_start_control_vars_in[4] = op_hcompute_conv_stencil_11_port_controller_d[4];
assign op_hcompute_conv_stencil_11_read_start_control_vars_in[3] = op_hcompute_conv_stencil_11_port_controller_d[3];
assign op_hcompute_conv_stencil_11_read_start_control_vars_in[2] = op_hcompute_conv_stencil_11_port_controller_d[2];
assign op_hcompute_conv_stencil_11_read_start_control_vars_in[1] = op_hcompute_conv_stencil_11_port_controller_d[1];
assign op_hcompute_conv_stencil_11_read_start_control_vars_in[0] = op_hcompute_conv_stencil_11_port_controller_d[0];
op_hcompute_conv_stencil_11_read_start_control_vars_pt__U999 op_hcompute_conv_stencil_11_read_start_control_vars (
    .in(op_hcompute_conv_stencil_11_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_11_read_start_control_vars_out)
);
op_hcompute_conv_stencil_11_write_start_pt__U1018 op_hcompute_conv_stencil_11_write_start (
    .in(delay_reg__U1035_out),
    .out(op_hcompute_conv_stencil_11_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_11_write_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_11_write_start_control_vars_in[4] = arr__U1149_out[4];
assign op_hcompute_conv_stencil_11_write_start_control_vars_in[3] = arr__U1149_out[3];
assign op_hcompute_conv_stencil_11_write_start_control_vars_in[2] = arr__U1149_out[2];
assign op_hcompute_conv_stencil_11_write_start_control_vars_in[1] = arr__U1149_out[1];
assign op_hcompute_conv_stencil_11_write_start_control_vars_in[0] = arr__U1149_out[0];
op_hcompute_conv_stencil_11_write_start_control_vars_pt__U1036 op_hcompute_conv_stencil_11_write_start_control_vars (
    .in(op_hcompute_conv_stencil_11_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_11_write_start_control_vars_out)
);
wire [15:0] op_hcompute_conv_stencil_12_conv_stencil_op_hcompute_conv_stencil_12_read [0:0];
assign op_hcompute_conv_stencil_12_conv_stencil_op_hcompute_conv_stencil_12_read[0] = conv_stencil_op_hcompute_conv_stencil_12_read[0];
wire [15:0] op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read [7:0];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[7];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[6];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[5];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[4];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[3];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[2];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[1];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[0];
wire [15:0] op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read [7:0];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[7];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[6];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[5];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[4];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[3];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[2];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[1];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[0];
cu_op_hcompute_conv_stencil_12 op_hcompute_conv_stencil_12 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_12_read(op_hcompute_conv_stencil_12_conv_stencil_op_hcompute_conv_stencil_12_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read(op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read(op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read),
    .conv_stencil_op_hcompute_conv_stencil_12_write(op_hcompute_conv_stencil_12_conv_stencil_op_hcompute_conv_stencil_12_write)
);
op_hcompute_conv_stencil_12_exe_start_pt__U1188 op_hcompute_conv_stencil_12_exe_start (
    .in(delay_reg__U1190_out),
    .out(op_hcompute_conv_stencil_12_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_12_exe_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_12_exe_start_control_vars_in[4] = arr__U1199_out[4];
assign op_hcompute_conv_stencil_12_exe_start_control_vars_in[3] = arr__U1199_out[3];
assign op_hcompute_conv_stencil_12_exe_start_control_vars_in[2] = arr__U1199_out[2];
assign op_hcompute_conv_stencil_12_exe_start_control_vars_in[1] = arr__U1199_out[1];
assign op_hcompute_conv_stencil_12_exe_start_control_vars_in[0] = arr__U1199_out[0];
op_hcompute_conv_stencil_12_exe_start_control_vars_pt__U1191 op_hcompute_conv_stencil_12_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_12_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_12_exe_start_control_vars_out)
);
affine_controller__U1156 op_hcompute_conv_stencil_12_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_12_port_controller_valid),
    .d(op_hcompute_conv_stencil_12_port_controller_d)
);
op_hcompute_conv_stencil_12_read_start_pt__U1186 op_hcompute_conv_stencil_12_read_start (
    .in(op_hcompute_conv_stencil_12_port_controller_valid),
    .out(op_hcompute_conv_stencil_12_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_12_read_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_12_read_start_control_vars_in[4] = op_hcompute_conv_stencil_12_port_controller_d[4];
assign op_hcompute_conv_stencil_12_read_start_control_vars_in[3] = op_hcompute_conv_stencil_12_port_controller_d[3];
assign op_hcompute_conv_stencil_12_read_start_control_vars_in[2] = op_hcompute_conv_stencil_12_port_controller_d[2];
assign op_hcompute_conv_stencil_12_read_start_control_vars_in[1] = op_hcompute_conv_stencil_12_port_controller_d[1];
assign op_hcompute_conv_stencil_12_read_start_control_vars_in[0] = op_hcompute_conv_stencil_12_port_controller_d[0];
op_hcompute_conv_stencil_12_read_start_control_vars_pt__U1187 op_hcompute_conv_stencil_12_read_start_control_vars (
    .in(op_hcompute_conv_stencil_12_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_12_read_start_control_vars_out)
);
op_hcompute_conv_stencil_12_write_start_pt__U1206 op_hcompute_conv_stencil_12_write_start (
    .in(delay_reg__U1223_out),
    .out(op_hcompute_conv_stencil_12_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_12_write_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_12_write_start_control_vars_in[4] = arr__U1337_out[4];
assign op_hcompute_conv_stencil_12_write_start_control_vars_in[3] = arr__U1337_out[3];
assign op_hcompute_conv_stencil_12_write_start_control_vars_in[2] = arr__U1337_out[2];
assign op_hcompute_conv_stencil_12_write_start_control_vars_in[1] = arr__U1337_out[1];
assign op_hcompute_conv_stencil_12_write_start_control_vars_in[0] = arr__U1337_out[0];
op_hcompute_conv_stencil_12_write_start_control_vars_pt__U1224 op_hcompute_conv_stencil_12_write_start_control_vars (
    .in(op_hcompute_conv_stencil_12_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_12_write_start_control_vars_out)
);
wire [15:0] op_hcompute_conv_stencil_13_conv_stencil_op_hcompute_conv_stencil_13_read [0:0];
assign op_hcompute_conv_stencil_13_conv_stencil_op_hcompute_conv_stencil_13_read[0] = conv_stencil_op_hcompute_conv_stencil_13_read[0];
wire [15:0] op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read [7:0];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[7];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[6];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[5];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[4];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[3];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[2];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[1];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[0];
wire [15:0] op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read [7:0];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[7];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[6];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[5];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[4];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[3];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[2];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[1];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[0];
cu_op_hcompute_conv_stencil_13 op_hcompute_conv_stencil_13 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_13_read(op_hcompute_conv_stencil_13_conv_stencil_op_hcompute_conv_stencil_13_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read(op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read(op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read),
    .conv_stencil_op_hcompute_conv_stencil_13_write(op_hcompute_conv_stencil_13_conv_stencil_op_hcompute_conv_stencil_13_write)
);
op_hcompute_conv_stencil_13_exe_start_pt__U1376 op_hcompute_conv_stencil_13_exe_start (
    .in(delay_reg__U1378_out),
    .out(op_hcompute_conv_stencil_13_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_13_exe_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_13_exe_start_control_vars_in[4] = arr__U1387_out[4];
assign op_hcompute_conv_stencil_13_exe_start_control_vars_in[3] = arr__U1387_out[3];
assign op_hcompute_conv_stencil_13_exe_start_control_vars_in[2] = arr__U1387_out[2];
assign op_hcompute_conv_stencil_13_exe_start_control_vars_in[1] = arr__U1387_out[1];
assign op_hcompute_conv_stencil_13_exe_start_control_vars_in[0] = arr__U1387_out[0];
op_hcompute_conv_stencil_13_exe_start_control_vars_pt__U1379 op_hcompute_conv_stencil_13_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_13_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_13_exe_start_control_vars_out)
);
affine_controller__U1344 op_hcompute_conv_stencil_13_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_13_port_controller_valid),
    .d(op_hcompute_conv_stencil_13_port_controller_d)
);
op_hcompute_conv_stencil_13_read_start_pt__U1374 op_hcompute_conv_stencil_13_read_start (
    .in(op_hcompute_conv_stencil_13_port_controller_valid),
    .out(op_hcompute_conv_stencil_13_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_13_read_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_13_read_start_control_vars_in[4] = op_hcompute_conv_stencil_13_port_controller_d[4];
assign op_hcompute_conv_stencil_13_read_start_control_vars_in[3] = op_hcompute_conv_stencil_13_port_controller_d[3];
assign op_hcompute_conv_stencil_13_read_start_control_vars_in[2] = op_hcompute_conv_stencil_13_port_controller_d[2];
assign op_hcompute_conv_stencil_13_read_start_control_vars_in[1] = op_hcompute_conv_stencil_13_port_controller_d[1];
assign op_hcompute_conv_stencil_13_read_start_control_vars_in[0] = op_hcompute_conv_stencil_13_port_controller_d[0];
op_hcompute_conv_stencil_13_read_start_control_vars_pt__U1375 op_hcompute_conv_stencil_13_read_start_control_vars (
    .in(op_hcompute_conv_stencil_13_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_13_read_start_control_vars_out)
);
op_hcompute_conv_stencil_13_write_start_pt__U1394 op_hcompute_conv_stencil_13_write_start (
    .in(delay_reg__U1411_out),
    .out(op_hcompute_conv_stencil_13_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_13_write_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_13_write_start_control_vars_in[4] = arr__U1525_out[4];
assign op_hcompute_conv_stencil_13_write_start_control_vars_in[3] = arr__U1525_out[3];
assign op_hcompute_conv_stencil_13_write_start_control_vars_in[2] = arr__U1525_out[2];
assign op_hcompute_conv_stencil_13_write_start_control_vars_in[1] = arr__U1525_out[1];
assign op_hcompute_conv_stencil_13_write_start_control_vars_in[0] = arr__U1525_out[0];
op_hcompute_conv_stencil_13_write_start_control_vars_pt__U1412 op_hcompute_conv_stencil_13_write_start_control_vars (
    .in(op_hcompute_conv_stencil_13_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_13_write_start_control_vars_out)
);
wire [15:0] op_hcompute_conv_stencil_14_conv_stencil_op_hcompute_conv_stencil_14_read [0:0];
assign op_hcompute_conv_stencil_14_conv_stencil_op_hcompute_conv_stencil_14_read[0] = conv_stencil_op_hcompute_conv_stencil_14_read[0];
wire [15:0] op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read [7:0];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[7];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[6];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[5];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[4];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[3];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[2];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[1];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[0];
wire [15:0] op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read [7:0];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[7];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[6];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[5];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[4];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[3];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[2];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[1];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[0];
cu_op_hcompute_conv_stencil_14 op_hcompute_conv_stencil_14 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_14_read(op_hcompute_conv_stencil_14_conv_stencil_op_hcompute_conv_stencil_14_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read(op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read(op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read),
    .conv_stencil_op_hcompute_conv_stencil_14_write(op_hcompute_conv_stencil_14_conv_stencil_op_hcompute_conv_stencil_14_write)
);
op_hcompute_conv_stencil_14_exe_start_pt__U1564 op_hcompute_conv_stencil_14_exe_start (
    .in(delay_reg__U1566_out),
    .out(op_hcompute_conv_stencil_14_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_14_exe_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_14_exe_start_control_vars_in[4] = arr__U1575_out[4];
assign op_hcompute_conv_stencil_14_exe_start_control_vars_in[3] = arr__U1575_out[3];
assign op_hcompute_conv_stencil_14_exe_start_control_vars_in[2] = arr__U1575_out[2];
assign op_hcompute_conv_stencil_14_exe_start_control_vars_in[1] = arr__U1575_out[1];
assign op_hcompute_conv_stencil_14_exe_start_control_vars_in[0] = arr__U1575_out[0];
op_hcompute_conv_stencil_14_exe_start_control_vars_pt__U1567 op_hcompute_conv_stencil_14_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_14_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_14_exe_start_control_vars_out)
);
affine_controller__U1532 op_hcompute_conv_stencil_14_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_14_port_controller_valid),
    .d(op_hcompute_conv_stencil_14_port_controller_d)
);
op_hcompute_conv_stencil_14_read_start_pt__U1562 op_hcompute_conv_stencil_14_read_start (
    .in(op_hcompute_conv_stencil_14_port_controller_valid),
    .out(op_hcompute_conv_stencil_14_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_14_read_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_14_read_start_control_vars_in[4] = op_hcompute_conv_stencil_14_port_controller_d[4];
assign op_hcompute_conv_stencil_14_read_start_control_vars_in[3] = op_hcompute_conv_stencil_14_port_controller_d[3];
assign op_hcompute_conv_stencil_14_read_start_control_vars_in[2] = op_hcompute_conv_stencil_14_port_controller_d[2];
assign op_hcompute_conv_stencil_14_read_start_control_vars_in[1] = op_hcompute_conv_stencil_14_port_controller_d[1];
assign op_hcompute_conv_stencil_14_read_start_control_vars_in[0] = op_hcompute_conv_stencil_14_port_controller_d[0];
op_hcompute_conv_stencil_14_read_start_control_vars_pt__U1563 op_hcompute_conv_stencil_14_read_start_control_vars (
    .in(op_hcompute_conv_stencil_14_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_14_read_start_control_vars_out)
);
op_hcompute_conv_stencil_14_write_start_pt__U1582 op_hcompute_conv_stencil_14_write_start (
    .in(delay_reg__U1599_out),
    .out(op_hcompute_conv_stencil_14_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_14_write_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_14_write_start_control_vars_in[4] = arr__U1713_out[4];
assign op_hcompute_conv_stencil_14_write_start_control_vars_in[3] = arr__U1713_out[3];
assign op_hcompute_conv_stencil_14_write_start_control_vars_in[2] = arr__U1713_out[2];
assign op_hcompute_conv_stencil_14_write_start_control_vars_in[1] = arr__U1713_out[1];
assign op_hcompute_conv_stencil_14_write_start_control_vars_in[0] = arr__U1713_out[0];
op_hcompute_conv_stencil_14_write_start_control_vars_pt__U1600 op_hcompute_conv_stencil_14_write_start_control_vars (
    .in(op_hcompute_conv_stencil_14_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_14_write_start_control_vars_out)
);
wire [15:0] op_hcompute_conv_stencil_15_conv_stencil_op_hcompute_conv_stencil_15_read [0:0];
assign op_hcompute_conv_stencil_15_conv_stencil_op_hcompute_conv_stencil_15_read[0] = conv_stencil_op_hcompute_conv_stencil_15_read[0];
wire [15:0] op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read [7:0];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[7];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[6];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[5];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[4];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[3];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[2];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[1];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[0];
wire [15:0] op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read [7:0];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[7];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[6];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[5];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[4];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[3];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[2];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[1];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[0];
cu_op_hcompute_conv_stencil_15 op_hcompute_conv_stencil_15 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_15_read(op_hcompute_conv_stencil_15_conv_stencil_op_hcompute_conv_stencil_15_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read(op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read(op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read),
    .conv_stencil_op_hcompute_conv_stencil_15_write(op_hcompute_conv_stencil_15_conv_stencil_op_hcompute_conv_stencil_15_write)
);
op_hcompute_conv_stencil_15_exe_start_pt__U1752 op_hcompute_conv_stencil_15_exe_start (
    .in(delay_reg__U1754_out),
    .out(op_hcompute_conv_stencil_15_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_15_exe_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_15_exe_start_control_vars_in[4] = arr__U1763_out[4];
assign op_hcompute_conv_stencil_15_exe_start_control_vars_in[3] = arr__U1763_out[3];
assign op_hcompute_conv_stencil_15_exe_start_control_vars_in[2] = arr__U1763_out[2];
assign op_hcompute_conv_stencil_15_exe_start_control_vars_in[1] = arr__U1763_out[1];
assign op_hcompute_conv_stencil_15_exe_start_control_vars_in[0] = arr__U1763_out[0];
op_hcompute_conv_stencil_15_exe_start_control_vars_pt__U1755 op_hcompute_conv_stencil_15_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_15_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_15_exe_start_control_vars_out)
);
affine_controller__U1720 op_hcompute_conv_stencil_15_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_15_port_controller_valid),
    .d(op_hcompute_conv_stencil_15_port_controller_d)
);
op_hcompute_conv_stencil_15_read_start_pt__U1750 op_hcompute_conv_stencil_15_read_start (
    .in(op_hcompute_conv_stencil_15_port_controller_valid),
    .out(op_hcompute_conv_stencil_15_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_15_read_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_15_read_start_control_vars_in[4] = op_hcompute_conv_stencil_15_port_controller_d[4];
assign op_hcompute_conv_stencil_15_read_start_control_vars_in[3] = op_hcompute_conv_stencil_15_port_controller_d[3];
assign op_hcompute_conv_stencil_15_read_start_control_vars_in[2] = op_hcompute_conv_stencil_15_port_controller_d[2];
assign op_hcompute_conv_stencil_15_read_start_control_vars_in[1] = op_hcompute_conv_stencil_15_port_controller_d[1];
assign op_hcompute_conv_stencil_15_read_start_control_vars_in[0] = op_hcompute_conv_stencil_15_port_controller_d[0];
op_hcompute_conv_stencil_15_read_start_control_vars_pt__U1751 op_hcompute_conv_stencil_15_read_start_control_vars (
    .in(op_hcompute_conv_stencil_15_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_15_read_start_control_vars_out)
);
op_hcompute_conv_stencil_15_write_start_pt__U1770 op_hcompute_conv_stencil_15_write_start (
    .in(delay_reg__U1787_out),
    .out(op_hcompute_conv_stencil_15_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_15_write_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_15_write_start_control_vars_in[4] = arr__U1901_out[4];
assign op_hcompute_conv_stencil_15_write_start_control_vars_in[3] = arr__U1901_out[3];
assign op_hcompute_conv_stencil_15_write_start_control_vars_in[2] = arr__U1901_out[2];
assign op_hcompute_conv_stencil_15_write_start_control_vars_in[1] = arr__U1901_out[1];
assign op_hcompute_conv_stencil_15_write_start_control_vars_in[0] = arr__U1901_out[0];
op_hcompute_conv_stencil_15_write_start_control_vars_pt__U1788 op_hcompute_conv_stencil_15_write_start_control_vars (
    .in(op_hcompute_conv_stencil_15_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_15_write_start_control_vars_out)
);
op_hcompute_conv_stencil_1_exe_start_pt__U262 op_hcompute_conv_stencil_1_exe_start (
    .in(op_hcompute_conv_stencil_1_port_controller_valid),
    .out(op_hcompute_conv_stencil_1_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U263 op_hcompute_conv_stencil_1_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_1_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_exe_start_control_vars_out)
);
affine_controller__U243 op_hcompute_conv_stencil_1_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_1_port_controller_valid),
    .d(op_hcompute_conv_stencil_1_port_controller_d)
);
op_hcompute_conv_stencil_1_read_start_pt__U260 op_hcompute_conv_stencil_1_read_start (
    .in(op_hcompute_conv_stencil_1_port_controller_valid),
    .out(op_hcompute_conv_stencil_1_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_read_start_control_vars_pt__U261 op_hcompute_conv_stencil_1_read_start_control_vars (
    .in(op_hcompute_conv_stencil_1_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_read_start_control_vars_out)
);
op_hcompute_conv_stencil_1_write_start_pt__U264 op_hcompute_conv_stencil_1_write_start (
    .in(op_hcompute_conv_stencil_1_port_controller_valid),
    .out(op_hcompute_conv_stencil_1_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_write_start_control_vars_pt__U265 op_hcompute_conv_stencil_1_write_start_control_vars (
    .in(op_hcompute_conv_stencil_1_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_write_start_control_vars_out)
);
cu_op_hcompute_conv_stencil_2 op_hcompute_conv_stencil_2 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_2_write(op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write)
);
op_hcompute_conv_stencil_2_exe_start_pt__U285 op_hcompute_conv_stencil_2_exe_start (
    .in(op_hcompute_conv_stencil_2_port_controller_valid),
    .out(op_hcompute_conv_stencil_2_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U286 op_hcompute_conv_stencil_2_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_2_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_exe_start_control_vars_out)
);
affine_controller__U266 op_hcompute_conv_stencil_2_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_2_port_controller_valid),
    .d(op_hcompute_conv_stencil_2_port_controller_d)
);
op_hcompute_conv_stencil_2_read_start_pt__U283 op_hcompute_conv_stencil_2_read_start (
    .in(op_hcompute_conv_stencil_2_port_controller_valid),
    .out(op_hcompute_conv_stencil_2_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_read_start_control_vars_pt__U284 op_hcompute_conv_stencil_2_read_start_control_vars (
    .in(op_hcompute_conv_stencil_2_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_read_start_control_vars_out)
);
op_hcompute_conv_stencil_2_write_start_pt__U287 op_hcompute_conv_stencil_2_write_start (
    .in(op_hcompute_conv_stencil_2_port_controller_valid),
    .out(op_hcompute_conv_stencil_2_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_write_start_control_vars_pt__U288 op_hcompute_conv_stencil_2_write_start_control_vars (
    .in(op_hcompute_conv_stencil_2_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_write_start_control_vars_out)
);
cu_op_hcompute_conv_stencil_3 op_hcompute_conv_stencil_3 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_3_write(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write)
);
op_hcompute_conv_stencil_3_exe_start_pt__U308 op_hcompute_conv_stencil_3_exe_start (
    .in(op_hcompute_conv_stencil_3_port_controller_valid),
    .out(op_hcompute_conv_stencil_3_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U309 op_hcompute_conv_stencil_3_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_3_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_exe_start_control_vars_out)
);
affine_controller__U289 op_hcompute_conv_stencil_3_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_3_port_controller_valid),
    .d(op_hcompute_conv_stencil_3_port_controller_d)
);
op_hcompute_conv_stencil_3_read_start_pt__U306 op_hcompute_conv_stencil_3_read_start (
    .in(op_hcompute_conv_stencil_3_port_controller_valid),
    .out(op_hcompute_conv_stencil_3_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
op_hcompute_conv_stencil_3_read_start_control_vars_pt__U307 op_hcompute_conv_stencil_3_read_start_control_vars (
    .in(op_hcompute_conv_stencil_3_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_read_start_control_vars_out)
);
op_hcompute_conv_stencil_3_write_start_pt__U310 op_hcompute_conv_stencil_3_write_start (
    .in(op_hcompute_conv_stencil_3_port_controller_valid),
    .out(op_hcompute_conv_stencil_3_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
op_hcompute_conv_stencil_3_write_start_control_vars_pt__U311 op_hcompute_conv_stencil_3_write_start_control_vars (
    .in(op_hcompute_conv_stencil_3_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_write_start_control_vars_out)
);
cu_op_hcompute_conv_stencil_4 op_hcompute_conv_stencil_4 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_4_write(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write)
);
op_hcompute_conv_stencil_4_exe_start_pt__U331 op_hcompute_conv_stencil_4_exe_start (
    .in(op_hcompute_conv_stencil_4_port_controller_valid),
    .out(op_hcompute_conv_stencil_4_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U332 op_hcompute_conv_stencil_4_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_4_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_exe_start_control_vars_out)
);
affine_controller__U312 op_hcompute_conv_stencil_4_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_4_port_controller_valid),
    .d(op_hcompute_conv_stencil_4_port_controller_d)
);
op_hcompute_conv_stencil_4_read_start_pt__U329 op_hcompute_conv_stencil_4_read_start (
    .in(op_hcompute_conv_stencil_4_port_controller_valid),
    .out(op_hcompute_conv_stencil_4_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
op_hcompute_conv_stencil_4_read_start_control_vars_pt__U330 op_hcompute_conv_stencil_4_read_start_control_vars (
    .in(op_hcompute_conv_stencil_4_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_read_start_control_vars_out)
);
op_hcompute_conv_stencil_4_write_start_pt__U333 op_hcompute_conv_stencil_4_write_start (
    .in(op_hcompute_conv_stencil_4_port_controller_valid),
    .out(op_hcompute_conv_stencil_4_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
op_hcompute_conv_stencil_4_write_start_control_vars_pt__U334 op_hcompute_conv_stencil_4_write_start_control_vars (
    .in(op_hcompute_conv_stencil_4_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_write_start_control_vars_out)
);
cu_op_hcompute_conv_stencil_5 op_hcompute_conv_stencil_5 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_5_write(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write)
);
op_hcompute_conv_stencil_5_exe_start_pt__U354 op_hcompute_conv_stencil_5_exe_start (
    .in(op_hcompute_conv_stencil_5_port_controller_valid),
    .out(op_hcompute_conv_stencil_5_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U355 op_hcompute_conv_stencil_5_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_5_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_exe_start_control_vars_out)
);
affine_controller__U335 op_hcompute_conv_stencil_5_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_5_port_controller_valid),
    .d(op_hcompute_conv_stencil_5_port_controller_d)
);
op_hcompute_conv_stencil_5_read_start_pt__U352 op_hcompute_conv_stencil_5_read_start (
    .in(op_hcompute_conv_stencil_5_port_controller_valid),
    .out(op_hcompute_conv_stencil_5_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
op_hcompute_conv_stencil_5_read_start_control_vars_pt__U353 op_hcompute_conv_stencil_5_read_start_control_vars (
    .in(op_hcompute_conv_stencil_5_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_read_start_control_vars_out)
);
op_hcompute_conv_stencil_5_write_start_pt__U356 op_hcompute_conv_stencil_5_write_start (
    .in(op_hcompute_conv_stencil_5_port_controller_valid),
    .out(op_hcompute_conv_stencil_5_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
op_hcompute_conv_stencil_5_write_start_control_vars_pt__U357 op_hcompute_conv_stencil_5_write_start_control_vars (
    .in(op_hcompute_conv_stencil_5_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_write_start_control_vars_out)
);
cu_op_hcompute_conv_stencil_6 op_hcompute_conv_stencil_6 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_6_write(op_hcompute_conv_stencil_6_conv_stencil_op_hcompute_conv_stencil_6_write)
);
op_hcompute_conv_stencil_6_exe_start_pt__U377 op_hcompute_conv_stencil_6_exe_start (
    .in(op_hcompute_conv_stencil_6_port_controller_valid),
    .out(op_hcompute_conv_stencil_6_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_6_exe_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_6_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_6_port_controller_d[2];
assign op_hcompute_conv_stencil_6_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_6_port_controller_d[1];
assign op_hcompute_conv_stencil_6_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_6_port_controller_d[0];
op_hcompute_conv_stencil_6_exe_start_control_vars_pt__U378 op_hcompute_conv_stencil_6_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_6_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_6_exe_start_control_vars_out)
);
affine_controller__U358 op_hcompute_conv_stencil_6_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_6_port_controller_valid),
    .d(op_hcompute_conv_stencil_6_port_controller_d)
);
op_hcompute_conv_stencil_6_read_start_pt__U375 op_hcompute_conv_stencil_6_read_start (
    .in(op_hcompute_conv_stencil_6_port_controller_valid),
    .out(op_hcompute_conv_stencil_6_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_6_read_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_6_read_start_control_vars_in[2] = op_hcompute_conv_stencil_6_port_controller_d[2];
assign op_hcompute_conv_stencil_6_read_start_control_vars_in[1] = op_hcompute_conv_stencil_6_port_controller_d[1];
assign op_hcompute_conv_stencil_6_read_start_control_vars_in[0] = op_hcompute_conv_stencil_6_port_controller_d[0];
op_hcompute_conv_stencil_6_read_start_control_vars_pt__U376 op_hcompute_conv_stencil_6_read_start_control_vars (
    .in(op_hcompute_conv_stencil_6_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_6_read_start_control_vars_out)
);
op_hcompute_conv_stencil_6_write_start_pt__U379 op_hcompute_conv_stencil_6_write_start (
    .in(op_hcompute_conv_stencil_6_port_controller_valid),
    .out(op_hcompute_conv_stencil_6_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_6_write_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_6_write_start_control_vars_in[2] = op_hcompute_conv_stencil_6_port_controller_d[2];
assign op_hcompute_conv_stencil_6_write_start_control_vars_in[1] = op_hcompute_conv_stencil_6_port_controller_d[1];
assign op_hcompute_conv_stencil_6_write_start_control_vars_in[0] = op_hcompute_conv_stencil_6_port_controller_d[0];
op_hcompute_conv_stencil_6_write_start_control_vars_pt__U380 op_hcompute_conv_stencil_6_write_start_control_vars (
    .in(op_hcompute_conv_stencil_6_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_6_write_start_control_vars_out)
);
cu_op_hcompute_conv_stencil_7 op_hcompute_conv_stencil_7 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_7_write(op_hcompute_conv_stencil_7_conv_stencil_op_hcompute_conv_stencil_7_write)
);
op_hcompute_conv_stencil_7_exe_start_pt__U400 op_hcompute_conv_stencil_7_exe_start (
    .in(op_hcompute_conv_stencil_7_port_controller_valid),
    .out(op_hcompute_conv_stencil_7_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_7_exe_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_7_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_7_port_controller_d[2];
assign op_hcompute_conv_stencil_7_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_7_port_controller_d[1];
assign op_hcompute_conv_stencil_7_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_7_port_controller_d[0];
op_hcompute_conv_stencil_7_exe_start_control_vars_pt__U401 op_hcompute_conv_stencil_7_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_7_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_7_exe_start_control_vars_out)
);
affine_controller__U381 op_hcompute_conv_stencil_7_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_7_port_controller_valid),
    .d(op_hcompute_conv_stencil_7_port_controller_d)
);
op_hcompute_conv_stencil_7_read_start_pt__U398 op_hcompute_conv_stencil_7_read_start (
    .in(op_hcompute_conv_stencil_7_port_controller_valid),
    .out(op_hcompute_conv_stencil_7_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_7_read_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_7_read_start_control_vars_in[2] = op_hcompute_conv_stencil_7_port_controller_d[2];
assign op_hcompute_conv_stencil_7_read_start_control_vars_in[1] = op_hcompute_conv_stencil_7_port_controller_d[1];
assign op_hcompute_conv_stencil_7_read_start_control_vars_in[0] = op_hcompute_conv_stencil_7_port_controller_d[0];
op_hcompute_conv_stencil_7_read_start_control_vars_pt__U399 op_hcompute_conv_stencil_7_read_start_control_vars (
    .in(op_hcompute_conv_stencil_7_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_7_read_start_control_vars_out)
);
op_hcompute_conv_stencil_7_write_start_pt__U402 op_hcompute_conv_stencil_7_write_start (
    .in(op_hcompute_conv_stencil_7_port_controller_valid),
    .out(op_hcompute_conv_stencil_7_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_7_write_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_7_write_start_control_vars_in[2] = op_hcompute_conv_stencil_7_port_controller_d[2];
assign op_hcompute_conv_stencil_7_write_start_control_vars_in[1] = op_hcompute_conv_stencil_7_port_controller_d[1];
assign op_hcompute_conv_stencil_7_write_start_control_vars_in[0] = op_hcompute_conv_stencil_7_port_controller_d[0];
op_hcompute_conv_stencil_7_write_start_control_vars_pt__U403 op_hcompute_conv_stencil_7_write_start_control_vars (
    .in(op_hcompute_conv_stencil_7_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_7_write_start_control_vars_out)
);
wire [15:0] op_hcompute_conv_stencil_8_conv_stencil_op_hcompute_conv_stencil_8_read [0:0];
assign op_hcompute_conv_stencil_8_conv_stencil_op_hcompute_conv_stencil_8_read[0] = conv_stencil_op_hcompute_conv_stencil_8_read[0];
wire [15:0] op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read [7:0];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[7];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[6];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[5];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[4];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[3];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[2];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[1];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[0];
wire [15:0] op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read [7:0];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[7];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[6];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[5];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[4];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[3];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[2];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[1];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[0];
cu_op_hcompute_conv_stencil_8 op_hcompute_conv_stencil_8 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_8_read(op_hcompute_conv_stencil_8_conv_stencil_op_hcompute_conv_stencil_8_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read(op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read(op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read),
    .conv_stencil_op_hcompute_conv_stencil_8_write(op_hcompute_conv_stencil_8_conv_stencil_op_hcompute_conv_stencil_8_write)
);
op_hcompute_conv_stencil_8_exe_start_pt__U436 op_hcompute_conv_stencil_8_exe_start (
    .in(delay_reg__U438_out),
    .out(op_hcompute_conv_stencil_8_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_8_exe_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_8_exe_start_control_vars_in[4] = arr__U447_out[4];
assign op_hcompute_conv_stencil_8_exe_start_control_vars_in[3] = arr__U447_out[3];
assign op_hcompute_conv_stencil_8_exe_start_control_vars_in[2] = arr__U447_out[2];
assign op_hcompute_conv_stencil_8_exe_start_control_vars_in[1] = arr__U447_out[1];
assign op_hcompute_conv_stencil_8_exe_start_control_vars_in[0] = arr__U447_out[0];
op_hcompute_conv_stencil_8_exe_start_control_vars_pt__U439 op_hcompute_conv_stencil_8_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_8_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_8_exe_start_control_vars_out)
);
affine_controller__U404 op_hcompute_conv_stencil_8_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_8_port_controller_valid),
    .d(op_hcompute_conv_stencil_8_port_controller_d)
);
op_hcompute_conv_stencil_8_read_start_pt__U434 op_hcompute_conv_stencil_8_read_start (
    .in(op_hcompute_conv_stencil_8_port_controller_valid),
    .out(op_hcompute_conv_stencil_8_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_8_read_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_8_read_start_control_vars_in[4] = op_hcompute_conv_stencil_8_port_controller_d[4];
assign op_hcompute_conv_stencil_8_read_start_control_vars_in[3] = op_hcompute_conv_stencil_8_port_controller_d[3];
assign op_hcompute_conv_stencil_8_read_start_control_vars_in[2] = op_hcompute_conv_stencil_8_port_controller_d[2];
assign op_hcompute_conv_stencil_8_read_start_control_vars_in[1] = op_hcompute_conv_stencil_8_port_controller_d[1];
assign op_hcompute_conv_stencil_8_read_start_control_vars_in[0] = op_hcompute_conv_stencil_8_port_controller_d[0];
op_hcompute_conv_stencil_8_read_start_control_vars_pt__U435 op_hcompute_conv_stencil_8_read_start_control_vars (
    .in(op_hcompute_conv_stencil_8_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_8_read_start_control_vars_out)
);
op_hcompute_conv_stencil_8_write_start_pt__U454 op_hcompute_conv_stencil_8_write_start (
    .in(delay_reg__U471_out),
    .out(op_hcompute_conv_stencil_8_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_8_write_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_8_write_start_control_vars_in[4] = arr__U585_out[4];
assign op_hcompute_conv_stencil_8_write_start_control_vars_in[3] = arr__U585_out[3];
assign op_hcompute_conv_stencil_8_write_start_control_vars_in[2] = arr__U585_out[2];
assign op_hcompute_conv_stencil_8_write_start_control_vars_in[1] = arr__U585_out[1];
assign op_hcompute_conv_stencil_8_write_start_control_vars_in[0] = arr__U585_out[0];
op_hcompute_conv_stencil_8_write_start_control_vars_pt__U472 op_hcompute_conv_stencil_8_write_start_control_vars (
    .in(op_hcompute_conv_stencil_8_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_8_write_start_control_vars_out)
);
wire [15:0] op_hcompute_conv_stencil_9_conv_stencil_op_hcompute_conv_stencil_9_read [0:0];
assign op_hcompute_conv_stencil_9_conv_stencil_op_hcompute_conv_stencil_9_read[0] = conv_stencil_op_hcompute_conv_stencil_9_read[0];
wire [15:0] op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read [7:0];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[7];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[6];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[5];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[4];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[3];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[2];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[1];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[0];
wire [15:0] op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read [7:0];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[7];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[6];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[5];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[4];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[3];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[2];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[1];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[0];
cu_op_hcompute_conv_stencil_9 op_hcompute_conv_stencil_9 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_9_read(op_hcompute_conv_stencil_9_conv_stencil_op_hcompute_conv_stencil_9_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read(op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read(op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read),
    .conv_stencil_op_hcompute_conv_stencil_9_write(op_hcompute_conv_stencil_9_conv_stencil_op_hcompute_conv_stencil_9_write)
);
op_hcompute_conv_stencil_9_exe_start_pt__U624 op_hcompute_conv_stencil_9_exe_start (
    .in(delay_reg__U626_out),
    .out(op_hcompute_conv_stencil_9_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_9_exe_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_9_exe_start_control_vars_in[4] = arr__U635_out[4];
assign op_hcompute_conv_stencil_9_exe_start_control_vars_in[3] = arr__U635_out[3];
assign op_hcompute_conv_stencil_9_exe_start_control_vars_in[2] = arr__U635_out[2];
assign op_hcompute_conv_stencil_9_exe_start_control_vars_in[1] = arr__U635_out[1];
assign op_hcompute_conv_stencil_9_exe_start_control_vars_in[0] = arr__U635_out[0];
op_hcompute_conv_stencil_9_exe_start_control_vars_pt__U627 op_hcompute_conv_stencil_9_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_9_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_9_exe_start_control_vars_out)
);
affine_controller__U592 op_hcompute_conv_stencil_9_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_9_port_controller_valid),
    .d(op_hcompute_conv_stencil_9_port_controller_d)
);
op_hcompute_conv_stencil_9_read_start_pt__U622 op_hcompute_conv_stencil_9_read_start (
    .in(op_hcompute_conv_stencil_9_port_controller_valid),
    .out(op_hcompute_conv_stencil_9_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_9_read_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_9_read_start_control_vars_in[4] = op_hcompute_conv_stencil_9_port_controller_d[4];
assign op_hcompute_conv_stencil_9_read_start_control_vars_in[3] = op_hcompute_conv_stencil_9_port_controller_d[3];
assign op_hcompute_conv_stencil_9_read_start_control_vars_in[2] = op_hcompute_conv_stencil_9_port_controller_d[2];
assign op_hcompute_conv_stencil_9_read_start_control_vars_in[1] = op_hcompute_conv_stencil_9_port_controller_d[1];
assign op_hcompute_conv_stencil_9_read_start_control_vars_in[0] = op_hcompute_conv_stencil_9_port_controller_d[0];
op_hcompute_conv_stencil_9_read_start_control_vars_pt__U623 op_hcompute_conv_stencil_9_read_start_control_vars (
    .in(op_hcompute_conv_stencil_9_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_9_read_start_control_vars_out)
);
op_hcompute_conv_stencil_9_write_start_pt__U642 op_hcompute_conv_stencil_9_write_start (
    .in(delay_reg__U659_out),
    .out(op_hcompute_conv_stencil_9_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_9_write_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_9_write_start_control_vars_in[4] = arr__U773_out[4];
assign op_hcompute_conv_stencil_9_write_start_control_vars_in[3] = arr__U773_out[3];
assign op_hcompute_conv_stencil_9_write_start_control_vars_in[2] = arr__U773_out[2];
assign op_hcompute_conv_stencil_9_write_start_control_vars_in[1] = arr__U773_out[1];
assign op_hcompute_conv_stencil_9_write_start_control_vars_in[0] = arr__U773_out[0];
op_hcompute_conv_stencil_9_write_start_control_vars_pt__U660 op_hcompute_conv_stencil_9_write_start_control_vars (
    .in(op_hcompute_conv_stencil_9_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_9_write_start_control_vars_out)
);
op_hcompute_conv_stencil_exe_start_pt__U239 op_hcompute_conv_stencil_exe_start (
    .in(op_hcompute_conv_stencil_port_controller_valid),
    .out(op_hcompute_conv_stencil_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_exe_start_control_vars_pt__U240 op_hcompute_conv_stencil_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_exe_start_control_vars_out)
);
affine_controller__U220 op_hcompute_conv_stencil_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_port_controller_valid),
    .d(op_hcompute_conv_stencil_port_controller_d)
);
op_hcompute_conv_stencil_read_start_pt__U237 op_hcompute_conv_stencil_read_start (
    .in(op_hcompute_conv_stencil_port_controller_valid),
    .out(op_hcompute_conv_stencil_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_read_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_read_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_read_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_read_start_control_vars_pt__U238 op_hcompute_conv_stencil_read_start_control_vars (
    .in(op_hcompute_conv_stencil_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_read_start_control_vars_out)
);
op_hcompute_conv_stencil_write_start_pt__U241 op_hcompute_conv_stencil_write_start (
    .in(op_hcompute_conv_stencil_port_controller_valid),
    .out(op_hcompute_conv_stencil_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_write_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_write_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_write_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_write_start_control_vars_pt__U242 op_hcompute_conv_stencil_write_start_control_vars (
    .in(op_hcompute_conv_stencil_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read [0:0];
assign op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read[0] = hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil op_hcompute_hw_input_global_wrapper_stencil (
    .clk(clk),
    .hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read(op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write(op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read [0:0];
assign op_hcompute_hw_input_global_wrapper_stencil_1_hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read[0] = hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil_1 op_hcompute_hw_input_global_wrapper_stencil_1 (
    .clk(clk),
    .hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read(op_hcompute_hw_input_global_wrapper_stencil_1_hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write(op_hcompute_hw_input_global_wrapper_stencil_1_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write)
);
op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_pt__U42 op_hcompute_hw_input_global_wrapper_stencil_1_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_pt__U43 op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_out)
);
affine_controller__U23 op_hcompute_hw_input_global_wrapper_stencil_1_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d)
);
op_hcompute_hw_input_global_wrapper_stencil_1_read_start_pt__U40 op_hcompute_hw_input_global_wrapper_stencil_1_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_valid),
    .out(hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read_en)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_pt__U41 op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_out)
);
op_hcompute_hw_input_global_wrapper_stencil_1_write_start_pt__U44 op_hcompute_hw_input_global_wrapper_stencil_1_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_1_write_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_pt__U45 op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read [0:0];
assign op_hcompute_hw_input_global_wrapper_stencil_2_hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read[0] = hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil_2 op_hcompute_hw_input_global_wrapper_stencil_2 (
    .clk(clk),
    .hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read(op_hcompute_hw_input_global_wrapper_stencil_2_hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write(op_hcompute_hw_input_global_wrapper_stencil_2_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write)
);
op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_pt__U65 op_hcompute_hw_input_global_wrapper_stencil_2_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_pt__U66 op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_out)
);
affine_controller__U46 op_hcompute_hw_input_global_wrapper_stencil_2_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d)
);
op_hcompute_hw_input_global_wrapper_stencil_2_read_start_pt__U63 op_hcompute_hw_input_global_wrapper_stencil_2_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_valid),
    .out(hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read_en)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_pt__U64 op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_out)
);
op_hcompute_hw_input_global_wrapper_stencil_2_write_start_pt__U67 op_hcompute_hw_input_global_wrapper_stencil_2_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_2_write_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_pt__U68 op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read [0:0];
assign op_hcompute_hw_input_global_wrapper_stencil_3_hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read[0] = hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil_3 op_hcompute_hw_input_global_wrapper_stencil_3 (
    .clk(clk),
    .hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read(op_hcompute_hw_input_global_wrapper_stencil_3_hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write(op_hcompute_hw_input_global_wrapper_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write)
);
op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_pt__U88 op_hcompute_hw_input_global_wrapper_stencil_3_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_pt__U89 op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_out)
);
affine_controller__U69 op_hcompute_hw_input_global_wrapper_stencil_3_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d)
);
op_hcompute_hw_input_global_wrapper_stencil_3_read_start_pt__U86 op_hcompute_hw_input_global_wrapper_stencil_3_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_valid),
    .out(hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read_en)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_pt__U87 op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_out)
);
op_hcompute_hw_input_global_wrapper_stencil_3_write_start_pt__U90 op_hcompute_hw_input_global_wrapper_stencil_3_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_3_write_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_pt__U91 op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read [0:0];
assign op_hcompute_hw_input_global_wrapper_stencil_4_hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read[0] = hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil_4 op_hcompute_hw_input_global_wrapper_stencil_4 (
    .clk(clk),
    .hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read(op_hcompute_hw_input_global_wrapper_stencil_4_hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write(op_hcompute_hw_input_global_wrapper_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write)
);
op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_pt__U111 op_hcompute_hw_input_global_wrapper_stencil_4_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_pt__U112 op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_out)
);
affine_controller__U92 op_hcompute_hw_input_global_wrapper_stencil_4_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d)
);
op_hcompute_hw_input_global_wrapper_stencil_4_read_start_pt__U109 op_hcompute_hw_input_global_wrapper_stencil_4_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_valid),
    .out(hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read_en)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_pt__U110 op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_out)
);
op_hcompute_hw_input_global_wrapper_stencil_4_write_start_pt__U113 op_hcompute_hw_input_global_wrapper_stencil_4_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_4_write_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_pt__U114 op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read [0:0];
assign op_hcompute_hw_input_global_wrapper_stencil_5_hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read[0] = hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil_5 op_hcompute_hw_input_global_wrapper_stencil_5 (
    .clk(clk),
    .hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read(op_hcompute_hw_input_global_wrapper_stencil_5_hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write(op_hcompute_hw_input_global_wrapper_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write)
);
op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_pt__U134 op_hcompute_hw_input_global_wrapper_stencil_5_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_pt__U135 op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_out)
);
affine_controller__U115 op_hcompute_hw_input_global_wrapper_stencil_5_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d)
);
op_hcompute_hw_input_global_wrapper_stencil_5_read_start_pt__U132 op_hcompute_hw_input_global_wrapper_stencil_5_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_valid),
    .out(hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read_en)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_pt__U133 op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_out)
);
op_hcompute_hw_input_global_wrapper_stencil_5_write_start_pt__U136 op_hcompute_hw_input_global_wrapper_stencil_5_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_5_write_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_pt__U137 op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read [0:0];
assign op_hcompute_hw_input_global_wrapper_stencil_6_hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read[0] = hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil_6 op_hcompute_hw_input_global_wrapper_stencil_6 (
    .clk(clk),
    .hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read(op_hcompute_hw_input_global_wrapper_stencil_6_hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write(op_hcompute_hw_input_global_wrapper_stencil_6_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write)
);
op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_pt__U157 op_hcompute_hw_input_global_wrapper_stencil_6_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_pt__U158 op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_out)
);
affine_controller__U138 op_hcompute_hw_input_global_wrapper_stencil_6_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d)
);
op_hcompute_hw_input_global_wrapper_stencil_6_read_start_pt__U155 op_hcompute_hw_input_global_wrapper_stencil_6_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_valid),
    .out(hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read_en)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_pt__U156 op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_out)
);
op_hcompute_hw_input_global_wrapper_stencil_6_write_start_pt__U159 op_hcompute_hw_input_global_wrapper_stencil_6_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_6_write_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_pt__U160 op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read [0:0];
assign op_hcompute_hw_input_global_wrapper_stencil_7_hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read[0] = hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil_7 op_hcompute_hw_input_global_wrapper_stencil_7 (
    .clk(clk),
    .hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read(op_hcompute_hw_input_global_wrapper_stencil_7_hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write(op_hcompute_hw_input_global_wrapper_stencil_7_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write)
);
op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_pt__U180 op_hcompute_hw_input_global_wrapper_stencil_7_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_pt__U181 op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_out)
);
affine_controller__U161 op_hcompute_hw_input_global_wrapper_stencil_7_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d)
);
op_hcompute_hw_input_global_wrapper_stencil_7_read_start_pt__U178 op_hcompute_hw_input_global_wrapper_stencil_7_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_valid),
    .out(hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read_en)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_pt__U179 op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_out)
);
op_hcompute_hw_input_global_wrapper_stencil_7_write_start_pt__U182 op_hcompute_hw_input_global_wrapper_stencil_7_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_7_write_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_pt__U183 op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_out)
);
op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U19 op_hcompute_hw_input_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U20 op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out)
);
affine_controller__U0 op_hcompute_hw_input_global_wrapper_stencil_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_port_controller_d)
);
op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U17 op_hcompute_hw_input_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .out(hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read_en)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U18 op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out)
);
op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U21 op_hcompute_hw_input_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in [2:0];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U22 op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0];
assign op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_kernel_global_wrapper_stencil op_hcompute_hw_kernel_global_wrapper_stencil (
    .clk(clk),
    .hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U216 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out)
);
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in [4:0];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U217 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out)
);
affine_controller__U184 op_hcompute_hw_kernel_global_wrapper_stencil_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d)
);
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U214 op_hcompute_hw_kernel_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .out(hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en)
);
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in [4:0];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U215 op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out)
);
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U218 op_hcompute_hw_kernel_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out)
);
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in [4:0];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U219 op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
assign op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
cu_op_hcompute_hw_output_stencil op_hcompute_hw_output_stencil (
    .clk(clk),
    .conv_stencil_op_hcompute_hw_output_stencil_read(op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read),
    .hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write(op_hcompute_hw_output_stencil_hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write)
);
wire [15:0] op_hcompute_hw_output_stencil_1_conv_stencil_op_hcompute_hw_output_stencil_1_read [0:0];
assign op_hcompute_hw_output_stencil_1_conv_stencil_op_hcompute_hw_output_stencil_1_read[0] = conv_stencil_op_hcompute_hw_output_stencil_1_read[0];
cu_op_hcompute_hw_output_stencil_1 op_hcompute_hw_output_stencil_1 (
    .clk(clk),
    .conv_stencil_op_hcompute_hw_output_stencil_1_read(op_hcompute_hw_output_stencil_1_conv_stencil_op_hcompute_hw_output_stencil_1_read),
    .hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write(op_hcompute_hw_output_stencil_1_hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write)
);
op_hcompute_hw_output_stencil_1_exe_start_pt__U1974 op_hcompute_hw_output_stencil_1_exe_start (
    .in(delay_reg__U1976_out),
    .out(op_hcompute_hw_output_stencil_1_exe_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_1_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_1_exe_start_control_vars_in[2] = arr__U1983_out[2];
assign op_hcompute_hw_output_stencil_1_exe_start_control_vars_in[1] = arr__U1983_out[1];
assign op_hcompute_hw_output_stencil_1_exe_start_control_vars_in[0] = arr__U1983_out[0];
op_hcompute_hw_output_stencil_1_exe_start_control_vars_pt__U1977 op_hcompute_hw_output_stencil_1_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_1_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_1_exe_start_control_vars_out)
);
affine_controller__U1955 op_hcompute_hw_output_stencil_1_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_output_stencil_1_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_1_port_controller_d)
);
op_hcompute_hw_output_stencil_1_read_start_pt__U1972 op_hcompute_hw_output_stencil_1_read_start (
    .in(op_hcompute_hw_output_stencil_1_port_controller_valid),
    .out(op_hcompute_hw_output_stencil_1_read_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_1_read_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_1_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_1_port_controller_d[2];
assign op_hcompute_hw_output_stencil_1_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_1_port_controller_d[1];
assign op_hcompute_hw_output_stencil_1_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_1_port_controller_d[0];
op_hcompute_hw_output_stencil_1_read_start_control_vars_pt__U1973 op_hcompute_hw_output_stencil_1_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_1_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_1_read_start_control_vars_out)
);
op_hcompute_hw_output_stencil_1_write_start_pt__U1988 op_hcompute_hw_output_stencil_1_write_start (
    .in(delay_reg__U1990_out),
    .out(hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write_valid)
);
wire [15:0] op_hcompute_hw_output_stencil_1_write_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_1_write_start_control_vars_in[2] = arr__U1997_out[2];
assign op_hcompute_hw_output_stencil_1_write_start_control_vars_in[1] = arr__U1997_out[1];
assign op_hcompute_hw_output_stencil_1_write_start_control_vars_in[0] = arr__U1997_out[0];
op_hcompute_hw_output_stencil_1_write_start_control_vars_pt__U1991 op_hcompute_hw_output_stencil_1_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_1_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_1_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_output_stencil_2_conv_stencil_op_hcompute_hw_output_stencil_2_read [0:0];
assign op_hcompute_hw_output_stencil_2_conv_stencil_op_hcompute_hw_output_stencil_2_read[0] = conv_stencil_op_hcompute_hw_output_stencil_2_read[0];
cu_op_hcompute_hw_output_stencil_2 op_hcompute_hw_output_stencil_2 (
    .clk(clk),
    .conv_stencil_op_hcompute_hw_output_stencil_2_read(op_hcompute_hw_output_stencil_2_conv_stencil_op_hcompute_hw_output_stencil_2_read),
    .hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write(op_hcompute_hw_output_stencil_2_hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write)
);
op_hcompute_hw_output_stencil_2_exe_start_pt__U2021 op_hcompute_hw_output_stencil_2_exe_start (
    .in(delay_reg__U2023_out),
    .out(op_hcompute_hw_output_stencil_2_exe_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_2_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_2_exe_start_control_vars_in[2] = arr__U2030_out[2];
assign op_hcompute_hw_output_stencil_2_exe_start_control_vars_in[1] = arr__U2030_out[1];
assign op_hcompute_hw_output_stencil_2_exe_start_control_vars_in[0] = arr__U2030_out[0];
op_hcompute_hw_output_stencil_2_exe_start_control_vars_pt__U2024 op_hcompute_hw_output_stencil_2_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_2_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_2_exe_start_control_vars_out)
);
affine_controller__U2002 op_hcompute_hw_output_stencil_2_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_output_stencil_2_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_2_port_controller_d)
);
op_hcompute_hw_output_stencil_2_read_start_pt__U2019 op_hcompute_hw_output_stencil_2_read_start (
    .in(op_hcompute_hw_output_stencil_2_port_controller_valid),
    .out(op_hcompute_hw_output_stencil_2_read_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_2_read_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_2_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_2_port_controller_d[2];
assign op_hcompute_hw_output_stencil_2_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_2_port_controller_d[1];
assign op_hcompute_hw_output_stencil_2_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_2_port_controller_d[0];
op_hcompute_hw_output_stencil_2_read_start_control_vars_pt__U2020 op_hcompute_hw_output_stencil_2_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_2_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_2_read_start_control_vars_out)
);
op_hcompute_hw_output_stencil_2_write_start_pt__U2035 op_hcompute_hw_output_stencil_2_write_start (
    .in(delay_reg__U2037_out),
    .out(hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write_valid)
);
wire [15:0] op_hcompute_hw_output_stencil_2_write_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_2_write_start_control_vars_in[2] = arr__U2044_out[2];
assign op_hcompute_hw_output_stencil_2_write_start_control_vars_in[1] = arr__U2044_out[1];
assign op_hcompute_hw_output_stencil_2_write_start_control_vars_in[0] = arr__U2044_out[0];
op_hcompute_hw_output_stencil_2_write_start_control_vars_pt__U2038 op_hcompute_hw_output_stencil_2_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_2_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_2_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_output_stencil_3_conv_stencil_op_hcompute_hw_output_stencil_3_read [0:0];
assign op_hcompute_hw_output_stencil_3_conv_stencil_op_hcompute_hw_output_stencil_3_read[0] = conv_stencil_op_hcompute_hw_output_stencil_3_read[0];
cu_op_hcompute_hw_output_stencil_3 op_hcompute_hw_output_stencil_3 (
    .clk(clk),
    .conv_stencil_op_hcompute_hw_output_stencil_3_read(op_hcompute_hw_output_stencil_3_conv_stencil_op_hcompute_hw_output_stencil_3_read),
    .hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write(op_hcompute_hw_output_stencil_3_hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write)
);
op_hcompute_hw_output_stencil_3_exe_start_pt__U2068 op_hcompute_hw_output_stencil_3_exe_start (
    .in(delay_reg__U2070_out),
    .out(op_hcompute_hw_output_stencil_3_exe_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_3_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_3_exe_start_control_vars_in[2] = arr__U2077_out[2];
assign op_hcompute_hw_output_stencil_3_exe_start_control_vars_in[1] = arr__U2077_out[1];
assign op_hcompute_hw_output_stencil_3_exe_start_control_vars_in[0] = arr__U2077_out[0];
op_hcompute_hw_output_stencil_3_exe_start_control_vars_pt__U2071 op_hcompute_hw_output_stencil_3_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_3_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_3_exe_start_control_vars_out)
);
affine_controller__U2049 op_hcompute_hw_output_stencil_3_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_output_stencil_3_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_3_port_controller_d)
);
op_hcompute_hw_output_stencil_3_read_start_pt__U2066 op_hcompute_hw_output_stencil_3_read_start (
    .in(op_hcompute_hw_output_stencil_3_port_controller_valid),
    .out(op_hcompute_hw_output_stencil_3_read_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_3_read_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_3_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_3_port_controller_d[2];
assign op_hcompute_hw_output_stencil_3_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_3_port_controller_d[1];
assign op_hcompute_hw_output_stencil_3_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_3_port_controller_d[0];
op_hcompute_hw_output_stencil_3_read_start_control_vars_pt__U2067 op_hcompute_hw_output_stencil_3_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_3_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_3_read_start_control_vars_out)
);
op_hcompute_hw_output_stencil_3_write_start_pt__U2082 op_hcompute_hw_output_stencil_3_write_start (
    .in(delay_reg__U2084_out),
    .out(hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write_valid)
);
wire [15:0] op_hcompute_hw_output_stencil_3_write_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_3_write_start_control_vars_in[2] = arr__U2091_out[2];
assign op_hcompute_hw_output_stencil_3_write_start_control_vars_in[1] = arr__U2091_out[1];
assign op_hcompute_hw_output_stencil_3_write_start_control_vars_in[0] = arr__U2091_out[0];
op_hcompute_hw_output_stencil_3_write_start_control_vars_pt__U2085 op_hcompute_hw_output_stencil_3_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_3_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_3_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_output_stencil_4_conv_stencil_op_hcompute_hw_output_stencil_4_read [0:0];
assign op_hcompute_hw_output_stencil_4_conv_stencil_op_hcompute_hw_output_stencil_4_read[0] = conv_stencil_op_hcompute_hw_output_stencil_4_read[0];
cu_op_hcompute_hw_output_stencil_4 op_hcompute_hw_output_stencil_4 (
    .clk(clk),
    .conv_stencil_op_hcompute_hw_output_stencil_4_read(op_hcompute_hw_output_stencil_4_conv_stencil_op_hcompute_hw_output_stencil_4_read),
    .hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write(op_hcompute_hw_output_stencil_4_hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write)
);
op_hcompute_hw_output_stencil_4_exe_start_pt__U2115 op_hcompute_hw_output_stencil_4_exe_start (
    .in(delay_reg__U2117_out),
    .out(op_hcompute_hw_output_stencil_4_exe_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_4_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_4_exe_start_control_vars_in[2] = arr__U2124_out[2];
assign op_hcompute_hw_output_stencil_4_exe_start_control_vars_in[1] = arr__U2124_out[1];
assign op_hcompute_hw_output_stencil_4_exe_start_control_vars_in[0] = arr__U2124_out[0];
op_hcompute_hw_output_stencil_4_exe_start_control_vars_pt__U2118 op_hcompute_hw_output_stencil_4_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_4_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_4_exe_start_control_vars_out)
);
affine_controller__U2096 op_hcompute_hw_output_stencil_4_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_output_stencil_4_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_4_port_controller_d)
);
op_hcompute_hw_output_stencil_4_read_start_pt__U2113 op_hcompute_hw_output_stencil_4_read_start (
    .in(op_hcompute_hw_output_stencil_4_port_controller_valid),
    .out(op_hcompute_hw_output_stencil_4_read_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_4_read_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_4_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_4_port_controller_d[2];
assign op_hcompute_hw_output_stencil_4_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_4_port_controller_d[1];
assign op_hcompute_hw_output_stencil_4_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_4_port_controller_d[0];
op_hcompute_hw_output_stencil_4_read_start_control_vars_pt__U2114 op_hcompute_hw_output_stencil_4_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_4_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_4_read_start_control_vars_out)
);
op_hcompute_hw_output_stencil_4_write_start_pt__U2129 op_hcompute_hw_output_stencil_4_write_start (
    .in(delay_reg__U2131_out),
    .out(hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write_valid)
);
wire [15:0] op_hcompute_hw_output_stencil_4_write_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_4_write_start_control_vars_in[2] = arr__U2138_out[2];
assign op_hcompute_hw_output_stencil_4_write_start_control_vars_in[1] = arr__U2138_out[1];
assign op_hcompute_hw_output_stencil_4_write_start_control_vars_in[0] = arr__U2138_out[0];
op_hcompute_hw_output_stencil_4_write_start_control_vars_pt__U2132 op_hcompute_hw_output_stencil_4_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_4_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_4_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_output_stencil_5_conv_stencil_op_hcompute_hw_output_stencil_5_read [0:0];
assign op_hcompute_hw_output_stencil_5_conv_stencil_op_hcompute_hw_output_stencil_5_read[0] = conv_stencil_op_hcompute_hw_output_stencil_5_read[0];
cu_op_hcompute_hw_output_stencil_5 op_hcompute_hw_output_stencil_5 (
    .clk(clk),
    .conv_stencil_op_hcompute_hw_output_stencil_5_read(op_hcompute_hw_output_stencil_5_conv_stencil_op_hcompute_hw_output_stencil_5_read),
    .hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write(op_hcompute_hw_output_stencil_5_hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write)
);
op_hcompute_hw_output_stencil_5_exe_start_pt__U2162 op_hcompute_hw_output_stencil_5_exe_start (
    .in(delay_reg__U2164_out),
    .out(op_hcompute_hw_output_stencil_5_exe_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_5_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_5_exe_start_control_vars_in[2] = arr__U2171_out[2];
assign op_hcompute_hw_output_stencil_5_exe_start_control_vars_in[1] = arr__U2171_out[1];
assign op_hcompute_hw_output_stencil_5_exe_start_control_vars_in[0] = arr__U2171_out[0];
op_hcompute_hw_output_stencil_5_exe_start_control_vars_pt__U2165 op_hcompute_hw_output_stencil_5_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_5_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_5_exe_start_control_vars_out)
);
affine_controller__U2143 op_hcompute_hw_output_stencil_5_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_output_stencil_5_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_5_port_controller_d)
);
op_hcompute_hw_output_stencil_5_read_start_pt__U2160 op_hcompute_hw_output_stencil_5_read_start (
    .in(op_hcompute_hw_output_stencil_5_port_controller_valid),
    .out(op_hcompute_hw_output_stencil_5_read_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_5_read_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_5_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_5_port_controller_d[2];
assign op_hcompute_hw_output_stencil_5_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_5_port_controller_d[1];
assign op_hcompute_hw_output_stencil_5_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_5_port_controller_d[0];
op_hcompute_hw_output_stencil_5_read_start_control_vars_pt__U2161 op_hcompute_hw_output_stencil_5_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_5_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_5_read_start_control_vars_out)
);
op_hcompute_hw_output_stencil_5_write_start_pt__U2176 op_hcompute_hw_output_stencil_5_write_start (
    .in(delay_reg__U2178_out),
    .out(hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write_valid)
);
wire [15:0] op_hcompute_hw_output_stencil_5_write_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_5_write_start_control_vars_in[2] = arr__U2185_out[2];
assign op_hcompute_hw_output_stencil_5_write_start_control_vars_in[1] = arr__U2185_out[1];
assign op_hcompute_hw_output_stencil_5_write_start_control_vars_in[0] = arr__U2185_out[0];
op_hcompute_hw_output_stencil_5_write_start_control_vars_pt__U2179 op_hcompute_hw_output_stencil_5_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_5_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_5_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_output_stencil_6_conv_stencil_op_hcompute_hw_output_stencil_6_read [0:0];
assign op_hcompute_hw_output_stencil_6_conv_stencil_op_hcompute_hw_output_stencil_6_read[0] = conv_stencil_op_hcompute_hw_output_stencil_6_read[0];
cu_op_hcompute_hw_output_stencil_6 op_hcompute_hw_output_stencil_6 (
    .clk(clk),
    .conv_stencil_op_hcompute_hw_output_stencil_6_read(op_hcompute_hw_output_stencil_6_conv_stencil_op_hcompute_hw_output_stencil_6_read),
    .hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write(op_hcompute_hw_output_stencil_6_hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write)
);
op_hcompute_hw_output_stencil_6_exe_start_pt__U2209 op_hcompute_hw_output_stencil_6_exe_start (
    .in(delay_reg__U2211_out),
    .out(op_hcompute_hw_output_stencil_6_exe_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_6_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_6_exe_start_control_vars_in[2] = arr__U2218_out[2];
assign op_hcompute_hw_output_stencil_6_exe_start_control_vars_in[1] = arr__U2218_out[1];
assign op_hcompute_hw_output_stencil_6_exe_start_control_vars_in[0] = arr__U2218_out[0];
op_hcompute_hw_output_stencil_6_exe_start_control_vars_pt__U2212 op_hcompute_hw_output_stencil_6_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_6_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_6_exe_start_control_vars_out)
);
affine_controller__U2190 op_hcompute_hw_output_stencil_6_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_output_stencil_6_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_6_port_controller_d)
);
op_hcompute_hw_output_stencil_6_read_start_pt__U2207 op_hcompute_hw_output_stencil_6_read_start (
    .in(op_hcompute_hw_output_stencil_6_port_controller_valid),
    .out(op_hcompute_hw_output_stencil_6_read_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_6_read_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_6_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_6_port_controller_d[2];
assign op_hcompute_hw_output_stencil_6_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_6_port_controller_d[1];
assign op_hcompute_hw_output_stencil_6_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_6_port_controller_d[0];
op_hcompute_hw_output_stencil_6_read_start_control_vars_pt__U2208 op_hcompute_hw_output_stencil_6_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_6_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_6_read_start_control_vars_out)
);
op_hcompute_hw_output_stencil_6_write_start_pt__U2223 op_hcompute_hw_output_stencil_6_write_start (
    .in(delay_reg__U2225_out),
    .out(hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write_valid)
);
wire [15:0] op_hcompute_hw_output_stencil_6_write_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_6_write_start_control_vars_in[2] = arr__U2232_out[2];
assign op_hcompute_hw_output_stencil_6_write_start_control_vars_in[1] = arr__U2232_out[1];
assign op_hcompute_hw_output_stencil_6_write_start_control_vars_in[0] = arr__U2232_out[0];
op_hcompute_hw_output_stencil_6_write_start_control_vars_pt__U2226 op_hcompute_hw_output_stencil_6_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_6_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_6_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_output_stencil_7_conv_stencil_op_hcompute_hw_output_stencil_7_read [0:0];
assign op_hcompute_hw_output_stencil_7_conv_stencil_op_hcompute_hw_output_stencil_7_read[0] = conv_stencil_op_hcompute_hw_output_stencil_7_read[0];
cu_op_hcompute_hw_output_stencil_7 op_hcompute_hw_output_stencil_7 (
    .clk(clk),
    .conv_stencil_op_hcompute_hw_output_stencil_7_read(op_hcompute_hw_output_stencil_7_conv_stencil_op_hcompute_hw_output_stencil_7_read),
    .hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write(op_hcompute_hw_output_stencil_7_hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write)
);
op_hcompute_hw_output_stencil_7_exe_start_pt__U2256 op_hcompute_hw_output_stencil_7_exe_start (
    .in(delay_reg__U2258_out),
    .out(op_hcompute_hw_output_stencil_7_exe_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_7_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_7_exe_start_control_vars_in[2] = arr__U2265_out[2];
assign op_hcompute_hw_output_stencil_7_exe_start_control_vars_in[1] = arr__U2265_out[1];
assign op_hcompute_hw_output_stencil_7_exe_start_control_vars_in[0] = arr__U2265_out[0];
op_hcompute_hw_output_stencil_7_exe_start_control_vars_pt__U2259 op_hcompute_hw_output_stencil_7_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_7_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_7_exe_start_control_vars_out)
);
affine_controller__U2237 op_hcompute_hw_output_stencil_7_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_output_stencil_7_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_7_port_controller_d)
);
op_hcompute_hw_output_stencil_7_read_start_pt__U2254 op_hcompute_hw_output_stencil_7_read_start (
    .in(op_hcompute_hw_output_stencil_7_port_controller_valid),
    .out(op_hcompute_hw_output_stencil_7_read_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_7_read_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_7_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_7_port_controller_d[2];
assign op_hcompute_hw_output_stencil_7_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_7_port_controller_d[1];
assign op_hcompute_hw_output_stencil_7_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_7_port_controller_d[0];
op_hcompute_hw_output_stencil_7_read_start_control_vars_pt__U2255 op_hcompute_hw_output_stencil_7_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_7_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_7_read_start_control_vars_out)
);
op_hcompute_hw_output_stencil_7_write_start_pt__U2270 op_hcompute_hw_output_stencil_7_write_start (
    .in(delay_reg__U2272_out),
    .out(hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write_valid)
);
wire [15:0] op_hcompute_hw_output_stencil_7_write_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_7_write_start_control_vars_in[2] = arr__U2279_out[2];
assign op_hcompute_hw_output_stencil_7_write_start_control_vars_in[1] = arr__U2279_out[1];
assign op_hcompute_hw_output_stencil_7_write_start_control_vars_in[0] = arr__U2279_out[0];
op_hcompute_hw_output_stencil_7_write_start_control_vars_pt__U2273 op_hcompute_hw_output_stencil_7_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_7_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_7_write_start_control_vars_out)
);
op_hcompute_hw_output_stencil_exe_start_pt__U1927 op_hcompute_hw_output_stencil_exe_start (
    .in(delay_reg__U1929_out),
    .out(op_hcompute_hw_output_stencil_exe_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[2] = arr__U1936_out[2];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[1] = arr__U1936_out[1];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[0] = arr__U1936_out[0];
op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U1930 op_hcompute_hw_output_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_exe_start_control_vars_out)
);
affine_controller__U1908 op_hcompute_hw_output_stencil_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_output_stencil_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_port_controller_d)
);
op_hcompute_hw_output_stencil_read_start_pt__U1925 op_hcompute_hw_output_stencil_read_start (
    .in(op_hcompute_hw_output_stencil_port_controller_valid),
    .out(op_hcompute_hw_output_stencil_read_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
op_hcompute_hw_output_stencil_read_start_control_vars_pt__U1926 op_hcompute_hw_output_stencil_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_read_start_control_vars_out)
);
op_hcompute_hw_output_stencil_write_start_pt__U1941 op_hcompute_hw_output_stencil_write_start (
    .in(delay_reg__U1943_out),
    .out(hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write_valid)
);
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_in [2:0];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[2] = arr__U1950_out[2];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[1] = arr__U1950_out[1];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[0] = arr__U1950_out[0];
op_hcompute_hw_output_stencil_write_start_control_vars_pt__U1944 op_hcompute_hw_output_stencil_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_write_start_control_vars_out)
);
assign hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write[0] = op_hcompute_hw_output_stencil_2_hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write[0];
assign hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write[0] = op_hcompute_hw_output_stencil_3_hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write[0];
assign hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write[0] = op_hcompute_hw_output_stencil_4_hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write[0];
assign hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write[0] = op_hcompute_hw_output_stencil_5_hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write[0];
assign hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write[0] = op_hcompute_hw_output_stencil_6_hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write[0];
assign hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write[0] = op_hcompute_hw_output_stencil_7_hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write[0];
assign hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write[0] = op_hcompute_hw_output_stencil_hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write[0];
assign hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write[0] = op_hcompute_hw_output_stencil_1_hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write[0];
endmodule

