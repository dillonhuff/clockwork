// Module `hw_kernel_global_wrapper_stencil_ub` defined externally
// Module `hw_input_global_wrapper_stencil_ub` defined externally
// Module `conv_stencil_ub` defined externally
module op_hcompute_hw_output_stencil_write_start_pt__U1941 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_write_start_control_vars_pt__U1944 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_read_start_pt__U1925 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_read_start_control_vars_pt__U1926 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_exe_start_pt__U1927 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U1930 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_7_write_start_pt__U2270 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_7_write_start_control_vars_pt__U2273 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_7_read_start_pt__U2254 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_7_read_start_control_vars_pt__U2255 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_7_exe_start_pt__U2256 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_7_exe_start_control_vars_pt__U2259 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_6_write_start_pt__U2223 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_6_write_start_control_vars_pt__U2226 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_6_read_start_pt__U2207 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_6_read_start_control_vars_pt__U2208 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_6_exe_start_pt__U2209 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_6_exe_start_control_vars_pt__U2212 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_5_write_start_pt__U2176 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_5_write_start_control_vars_pt__U2179 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_5_read_start_pt__U2160 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_5_read_start_control_vars_pt__U2161 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_5_exe_start_pt__U2162 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_5_exe_start_control_vars_pt__U2165 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_4_write_start_pt__U2129 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_4_write_start_control_vars_pt__U2132 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_4_read_start_pt__U2113 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_4_read_start_control_vars_pt__U2114 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_4_exe_start_pt__U2115 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_4_exe_start_control_vars_pt__U2118 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_3_write_start_pt__U2082 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_3_write_start_control_vars_pt__U2085 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_3_read_start_pt__U2066 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_3_read_start_control_vars_pt__U2067 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_3_exe_start_pt__U2068 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_3_exe_start_control_vars_pt__U2071 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_2_write_start_pt__U2035 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_2_write_start_control_vars_pt__U2038 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_2_read_start_pt__U2019 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_2_read_start_control_vars_pt__U2020 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_2_exe_start_pt__U2021 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_2_exe_start_control_vars_pt__U2024 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_1_write_start_pt__U1988 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_1_write_start_control_vars_pt__U1991 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_1_read_start_pt__U1972 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_1_read_start_control_vars_pt__U1973 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_1_exe_start_pt__U1974 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_1_exe_start_control_vars_pt__U1977 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U218 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U219 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U214 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U215 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U216 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U217 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U21 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U22 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U17 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U18 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U19 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U20 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_7_write_start_pt__U182 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_pt__U183 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_7_read_start_pt__U178 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_pt__U179 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_pt__U180 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_pt__U181 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_6_write_start_pt__U159 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_pt__U160 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_6_read_start_pt__U155 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_pt__U156 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_pt__U157 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_pt__U158 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_5_write_start_pt__U136 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_pt__U137 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_5_read_start_pt__U132 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_pt__U133 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_pt__U134 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_pt__U135 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_4_write_start_pt__U113 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_pt__U114 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_4_read_start_pt__U109 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_pt__U110 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_pt__U111 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_pt__U112 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_3_write_start_pt__U90 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_pt__U91 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_3_read_start_pt__U86 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_pt__U87 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_pt__U88 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_pt__U89 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_2_write_start_pt__U67 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_pt__U68 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_2_read_start_pt__U63 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_pt__U64 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_pt__U65 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_pt__U66 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_1_write_start_pt__U44 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_pt__U45 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_1_read_start_pt__U40 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_pt__U41 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_pt__U42 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_pt__U43 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_write_start_pt__U241 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_write_start_control_vars_pt__U242 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_read_start_pt__U237 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_read_start_control_vars_pt__U238 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_exe_start_pt__U239 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_exe_start_control_vars_pt__U240 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_9_write_start_pt__U642 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_9_write_start_control_vars_pt__U660 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_9_read_start_pt__U622 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_9_read_start_control_vars_pt__U623 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_9_exe_start_pt__U624 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_9_exe_start_control_vars_pt__U627 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_8_write_start_pt__U454 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_8_write_start_control_vars_pt__U472 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_8_read_start_pt__U434 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_8_read_start_control_vars_pt__U435 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_8_exe_start_pt__U436 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_8_exe_start_control_vars_pt__U439 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_7_write_start_pt__U402 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_7_write_start_control_vars_pt__U403 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_7_read_start_pt__U398 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_7_read_start_control_vars_pt__U399 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_7_exe_start_pt__U400 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_7_exe_start_control_vars_pt__U401 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_6_write_start_pt__U379 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_6_write_start_control_vars_pt__U380 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_6_read_start_pt__U375 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_6_read_start_control_vars_pt__U376 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_6_exe_start_pt__U377 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_6_exe_start_control_vars_pt__U378 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_write_start_pt__U356 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_write_start_control_vars_pt__U357 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_read_start_pt__U352 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_read_start_control_vars_pt__U353 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_exe_start_pt__U354 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U355 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_write_start_pt__U333 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_write_start_control_vars_pt__U334 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_read_start_pt__U329 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_read_start_control_vars_pt__U330 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_exe_start_pt__U331 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U332 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_write_start_pt__U310 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_write_start_control_vars_pt__U311 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_read_start_pt__U306 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_read_start_control_vars_pt__U307 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_exe_start_pt__U308 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U309 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_write_start_pt__U287 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_write_start_control_vars_pt__U288 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_read_start_pt__U283 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_read_start_control_vars_pt__U284 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_exe_start_pt__U285 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U286 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_write_start_pt__U264 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_write_start_control_vars_pt__U265 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_read_start_pt__U260 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_read_start_control_vars_pt__U261 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_exe_start_pt__U262 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U263 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_15_write_start_pt__U1770 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_15_write_start_control_vars_pt__U1788 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_15_read_start_pt__U1750 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_15_read_start_control_vars_pt__U1751 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_15_exe_start_pt__U1752 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_15_exe_start_control_vars_pt__U1755 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_14_write_start_pt__U1582 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_14_write_start_control_vars_pt__U1600 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_14_read_start_pt__U1562 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_14_read_start_control_vars_pt__U1563 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_14_exe_start_pt__U1564 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_14_exe_start_control_vars_pt__U1567 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_13_write_start_pt__U1394 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_13_write_start_control_vars_pt__U1412 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_13_read_start_pt__U1374 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_13_read_start_control_vars_pt__U1375 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_13_exe_start_pt__U1376 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_13_exe_start_control_vars_pt__U1379 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_12_write_start_pt__U1206 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_12_write_start_control_vars_pt__U1224 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_12_read_start_pt__U1186 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_12_read_start_control_vars_pt__U1187 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_12_exe_start_pt__U1188 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_12_exe_start_control_vars_pt__U1191 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_11_write_start_pt__U1018 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_11_write_start_control_vars_pt__U1036 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_11_read_start_pt__U998 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_11_read_start_control_vars_pt__U999 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_11_exe_start_pt__U1000 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_11_exe_start_control_vars_pt__U1003 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_10_write_start_pt__U830 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_10_write_start_control_vars_pt__U848 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_10_read_start_pt__U810 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_10_read_start_control_vars_pt__U811 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_10_exe_start_pt__U812 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_10_exe_start_control_vars_pt__U815 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module coreir_reg #(
    parameter width = 1,
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input [width-1:0] in,
    output [width-1:0] out
);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out
);
wire reg0_clk;
wire [15:0] reg0_in;
assign reg0_clk = clk;
assign reg0_in = in;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(reg0_clk),
    .in(reg0_in),
    .out(out)
);
endmodule

module mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out,
    input en
);
wire reg0_clk;
wire [15:0] reg0_in;
assign reg0_clk = clk;
assign reg0_in = en ? in : out;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(reg0_clk),
    .in(reg0_in),
    .out(out)
);
endmodule

module corebit_reg #(
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input in,
    output out
);
reg outReg = init;
always @(posedge clk) begin
  outReg <= in;
end
assign out = outReg;
endmodule

module array_delay_U962 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U963_in;
wire _U963_clk;
wire [15:0] _U963_out;
wire [15:0] _U964_in;
wire _U964_clk;
wire [15:0] _U964_out;
wire [15:0] _U965_in;
wire _U965_clk;
wire [15:0] _U965_out;
wire [15:0] _U966_in;
wire _U966_clk;
wire [15:0] _U966_out;
wire [15:0] _U967_in;
wire _U967_clk;
wire [15:0] _U967_out;
assign _U963_in = in[0];
assign _U963_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U963 (
    .in(_U963_in),
    .clk(_U963_clk),
    .out(_U963_out)
);
assign _U964_in = in[1];
assign _U964_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U964 (
    .in(_U964_in),
    .clk(_U964_clk),
    .out(_U964_out)
);
assign _U965_in = in[2];
assign _U965_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U965 (
    .in(_U965_in),
    .clk(_U965_clk),
    .out(_U965_out)
);
assign _U966_in = in[3];
assign _U966_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U966 (
    .in(_U966_in),
    .clk(_U966_clk),
    .out(_U966_out)
);
assign _U967_in = in[4];
assign _U967_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U967 (
    .in(_U967_in),
    .clk(_U967_clk),
    .out(_U967_out)
);
assign out[4] = _U967_out;
assign out[3] = _U966_out;
assign out[2] = _U965_out;
assign out[1] = _U964_out;
assign out[0] = _U963_out;
endmodule

module array_delay_U955 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U956_in;
wire _U956_clk;
wire [15:0] _U956_out;
wire [15:0] _U957_in;
wire _U957_clk;
wire [15:0] _U957_out;
wire [15:0] _U958_in;
wire _U958_clk;
wire [15:0] _U958_out;
wire [15:0] _U959_in;
wire _U959_clk;
wire [15:0] _U959_out;
wire [15:0] _U960_in;
wire _U960_clk;
wire [15:0] _U960_out;
assign _U956_in = in[0];
assign _U956_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U956 (
    .in(_U956_in),
    .clk(_U956_clk),
    .out(_U956_out)
);
assign _U957_in = in[1];
assign _U957_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U957 (
    .in(_U957_in),
    .clk(_U957_clk),
    .out(_U957_out)
);
assign _U958_in = in[2];
assign _U958_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U958 (
    .in(_U958_in),
    .clk(_U958_clk),
    .out(_U958_out)
);
assign _U959_in = in[3];
assign _U959_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U959 (
    .in(_U959_in),
    .clk(_U959_clk),
    .out(_U959_out)
);
assign _U960_in = in[4];
assign _U960_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U960 (
    .in(_U960_in),
    .clk(_U960_clk),
    .out(_U960_out)
);
assign out[4] = _U960_out;
assign out[3] = _U959_out;
assign out[2] = _U958_out;
assign out[1] = _U957_out;
assign out[0] = _U956_out;
endmodule

module array_delay_U948 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U949_in;
wire _U949_clk;
wire [15:0] _U949_out;
wire [15:0] _U950_in;
wire _U950_clk;
wire [15:0] _U950_out;
wire [15:0] _U951_in;
wire _U951_clk;
wire [15:0] _U951_out;
wire [15:0] _U952_in;
wire _U952_clk;
wire [15:0] _U952_out;
wire [15:0] _U953_in;
wire _U953_clk;
wire [15:0] _U953_out;
assign _U949_in = in[0];
assign _U949_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U949 (
    .in(_U949_in),
    .clk(_U949_clk),
    .out(_U949_out)
);
assign _U950_in = in[1];
assign _U950_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U950 (
    .in(_U950_in),
    .clk(_U950_clk),
    .out(_U950_out)
);
assign _U951_in = in[2];
assign _U951_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U951 (
    .in(_U951_in),
    .clk(_U951_clk),
    .out(_U951_out)
);
assign _U952_in = in[3];
assign _U952_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U952 (
    .in(_U952_in),
    .clk(_U952_clk),
    .out(_U952_out)
);
assign _U953_in = in[4];
assign _U953_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U953 (
    .in(_U953_in),
    .clk(_U953_clk),
    .out(_U953_out)
);
assign out[4] = _U953_out;
assign out[3] = _U952_out;
assign out[2] = _U951_out;
assign out[1] = _U950_out;
assign out[0] = _U949_out;
endmodule

module array_delay_U941 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U942_in;
wire _U942_clk;
wire [15:0] _U942_out;
wire [15:0] _U943_in;
wire _U943_clk;
wire [15:0] _U943_out;
wire [15:0] _U944_in;
wire _U944_clk;
wire [15:0] _U944_out;
wire [15:0] _U945_in;
wire _U945_clk;
wire [15:0] _U945_out;
wire [15:0] _U946_in;
wire _U946_clk;
wire [15:0] _U946_out;
assign _U942_in = in[0];
assign _U942_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U942 (
    .in(_U942_in),
    .clk(_U942_clk),
    .out(_U942_out)
);
assign _U943_in = in[1];
assign _U943_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U943 (
    .in(_U943_in),
    .clk(_U943_clk),
    .out(_U943_out)
);
assign _U944_in = in[2];
assign _U944_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U944 (
    .in(_U944_in),
    .clk(_U944_clk),
    .out(_U944_out)
);
assign _U945_in = in[3];
assign _U945_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U945 (
    .in(_U945_in),
    .clk(_U945_clk),
    .out(_U945_out)
);
assign _U946_in = in[4];
assign _U946_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U946 (
    .in(_U946_in),
    .clk(_U946_clk),
    .out(_U946_out)
);
assign out[4] = _U946_out;
assign out[3] = _U945_out;
assign out[2] = _U944_out;
assign out[1] = _U943_out;
assign out[0] = _U942_out;
endmodule

module array_delay_U934 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U935_in;
wire _U935_clk;
wire [15:0] _U935_out;
wire [15:0] _U936_in;
wire _U936_clk;
wire [15:0] _U936_out;
wire [15:0] _U937_in;
wire _U937_clk;
wire [15:0] _U937_out;
wire [15:0] _U938_in;
wire _U938_clk;
wire [15:0] _U938_out;
wire [15:0] _U939_in;
wire _U939_clk;
wire [15:0] _U939_out;
assign _U935_in = in[0];
assign _U935_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U935 (
    .in(_U935_in),
    .clk(_U935_clk),
    .out(_U935_out)
);
assign _U936_in = in[1];
assign _U936_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U936 (
    .in(_U936_in),
    .clk(_U936_clk),
    .out(_U936_out)
);
assign _U937_in = in[2];
assign _U937_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U937 (
    .in(_U937_in),
    .clk(_U937_clk),
    .out(_U937_out)
);
assign _U938_in = in[3];
assign _U938_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U938 (
    .in(_U938_in),
    .clk(_U938_clk),
    .out(_U938_out)
);
assign _U939_in = in[4];
assign _U939_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U939 (
    .in(_U939_in),
    .clk(_U939_clk),
    .out(_U939_out)
);
assign out[4] = _U939_out;
assign out[3] = _U938_out;
assign out[2] = _U937_out;
assign out[1] = _U936_out;
assign out[0] = _U935_out;
endmodule

module array_delay_U927 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U928_in;
wire _U928_clk;
wire [15:0] _U928_out;
wire [15:0] _U929_in;
wire _U929_clk;
wire [15:0] _U929_out;
wire [15:0] _U930_in;
wire _U930_clk;
wire [15:0] _U930_out;
wire [15:0] _U931_in;
wire _U931_clk;
wire [15:0] _U931_out;
wire [15:0] _U932_in;
wire _U932_clk;
wire [15:0] _U932_out;
assign _U928_in = in[0];
assign _U928_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U928 (
    .in(_U928_in),
    .clk(_U928_clk),
    .out(_U928_out)
);
assign _U929_in = in[1];
assign _U929_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U929 (
    .in(_U929_in),
    .clk(_U929_clk),
    .out(_U929_out)
);
assign _U930_in = in[2];
assign _U930_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U930 (
    .in(_U930_in),
    .clk(_U930_clk),
    .out(_U930_out)
);
assign _U931_in = in[3];
assign _U931_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U931 (
    .in(_U931_in),
    .clk(_U931_clk),
    .out(_U931_out)
);
assign _U932_in = in[4];
assign _U932_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U932 (
    .in(_U932_in),
    .clk(_U932_clk),
    .out(_U932_out)
);
assign out[4] = _U932_out;
assign out[3] = _U931_out;
assign out[2] = _U930_out;
assign out[1] = _U929_out;
assign out[0] = _U928_out;
endmodule

module array_delay_U920 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U921_in;
wire _U921_clk;
wire [15:0] _U921_out;
wire [15:0] _U922_in;
wire _U922_clk;
wire [15:0] _U922_out;
wire [15:0] _U923_in;
wire _U923_clk;
wire [15:0] _U923_out;
wire [15:0] _U924_in;
wire _U924_clk;
wire [15:0] _U924_out;
wire [15:0] _U925_in;
wire _U925_clk;
wire [15:0] _U925_out;
assign _U921_in = in[0];
assign _U921_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U921 (
    .in(_U921_in),
    .clk(_U921_clk),
    .out(_U921_out)
);
assign _U922_in = in[1];
assign _U922_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U922 (
    .in(_U922_in),
    .clk(_U922_clk),
    .out(_U922_out)
);
assign _U923_in = in[2];
assign _U923_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U923 (
    .in(_U923_in),
    .clk(_U923_clk),
    .out(_U923_out)
);
assign _U924_in = in[3];
assign _U924_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U924 (
    .in(_U924_in),
    .clk(_U924_clk),
    .out(_U924_out)
);
assign _U925_in = in[4];
assign _U925_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U925 (
    .in(_U925_in),
    .clk(_U925_clk),
    .out(_U925_out)
);
assign out[4] = _U925_out;
assign out[3] = _U924_out;
assign out[2] = _U923_out;
assign out[1] = _U922_out;
assign out[0] = _U921_out;
endmodule

module array_delay_U913 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U914_in;
wire _U914_clk;
wire [15:0] _U914_out;
wire [15:0] _U915_in;
wire _U915_clk;
wire [15:0] _U915_out;
wire [15:0] _U916_in;
wire _U916_clk;
wire [15:0] _U916_out;
wire [15:0] _U917_in;
wire _U917_clk;
wire [15:0] _U917_out;
wire [15:0] _U918_in;
wire _U918_clk;
wire [15:0] _U918_out;
assign _U914_in = in[0];
assign _U914_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U914 (
    .in(_U914_in),
    .clk(_U914_clk),
    .out(_U914_out)
);
assign _U915_in = in[1];
assign _U915_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U915 (
    .in(_U915_in),
    .clk(_U915_clk),
    .out(_U915_out)
);
assign _U916_in = in[2];
assign _U916_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U916 (
    .in(_U916_in),
    .clk(_U916_clk),
    .out(_U916_out)
);
assign _U917_in = in[3];
assign _U917_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U917 (
    .in(_U917_in),
    .clk(_U917_clk),
    .out(_U917_out)
);
assign _U918_in = in[4];
assign _U918_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U918 (
    .in(_U918_in),
    .clk(_U918_clk),
    .out(_U918_out)
);
assign out[4] = _U918_out;
assign out[3] = _U917_out;
assign out[2] = _U916_out;
assign out[1] = _U915_out;
assign out[0] = _U914_out;
endmodule

module array_delay_U906 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U907_in;
wire _U907_clk;
wire [15:0] _U907_out;
wire [15:0] _U908_in;
wire _U908_clk;
wire [15:0] _U908_out;
wire [15:0] _U909_in;
wire _U909_clk;
wire [15:0] _U909_out;
wire [15:0] _U910_in;
wire _U910_clk;
wire [15:0] _U910_out;
wire [15:0] _U911_in;
wire _U911_clk;
wire [15:0] _U911_out;
assign _U907_in = in[0];
assign _U907_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U907 (
    .in(_U907_in),
    .clk(_U907_clk),
    .out(_U907_out)
);
assign _U908_in = in[1];
assign _U908_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U908 (
    .in(_U908_in),
    .clk(_U908_clk),
    .out(_U908_out)
);
assign _U909_in = in[2];
assign _U909_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U909 (
    .in(_U909_in),
    .clk(_U909_clk),
    .out(_U909_out)
);
assign _U910_in = in[3];
assign _U910_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U910 (
    .in(_U910_in),
    .clk(_U910_clk),
    .out(_U910_out)
);
assign _U911_in = in[4];
assign _U911_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U911 (
    .in(_U911_in),
    .clk(_U911_clk),
    .out(_U911_out)
);
assign out[4] = _U911_out;
assign out[3] = _U910_out;
assign out[2] = _U909_out;
assign out[1] = _U908_out;
assign out[0] = _U907_out;
endmodule

module array_delay_U899 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U900_in;
wire _U900_clk;
wire [15:0] _U900_out;
wire [15:0] _U901_in;
wire _U901_clk;
wire [15:0] _U901_out;
wire [15:0] _U902_in;
wire _U902_clk;
wire [15:0] _U902_out;
wire [15:0] _U903_in;
wire _U903_clk;
wire [15:0] _U903_out;
wire [15:0] _U904_in;
wire _U904_clk;
wire [15:0] _U904_out;
assign _U900_in = in[0];
assign _U900_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U900 (
    .in(_U900_in),
    .clk(_U900_clk),
    .out(_U900_out)
);
assign _U901_in = in[1];
assign _U901_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U901 (
    .in(_U901_in),
    .clk(_U901_clk),
    .out(_U901_out)
);
assign _U902_in = in[2];
assign _U902_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U902 (
    .in(_U902_in),
    .clk(_U902_clk),
    .out(_U902_out)
);
assign _U903_in = in[3];
assign _U903_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U903 (
    .in(_U903_in),
    .clk(_U903_clk),
    .out(_U903_out)
);
assign _U904_in = in[4];
assign _U904_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U904 (
    .in(_U904_in),
    .clk(_U904_clk),
    .out(_U904_out)
);
assign out[4] = _U904_out;
assign out[3] = _U903_out;
assign out[2] = _U902_out;
assign out[1] = _U901_out;
assign out[0] = _U900_out;
endmodule

module array_delay_U892 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U893_in;
wire _U893_clk;
wire [15:0] _U893_out;
wire [15:0] _U894_in;
wire _U894_clk;
wire [15:0] _U894_out;
wire [15:0] _U895_in;
wire _U895_clk;
wire [15:0] _U895_out;
wire [15:0] _U896_in;
wire _U896_clk;
wire [15:0] _U896_out;
wire [15:0] _U897_in;
wire _U897_clk;
wire [15:0] _U897_out;
assign _U893_in = in[0];
assign _U893_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U893 (
    .in(_U893_in),
    .clk(_U893_clk),
    .out(_U893_out)
);
assign _U894_in = in[1];
assign _U894_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U894 (
    .in(_U894_in),
    .clk(_U894_clk),
    .out(_U894_out)
);
assign _U895_in = in[2];
assign _U895_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U895 (
    .in(_U895_in),
    .clk(_U895_clk),
    .out(_U895_out)
);
assign _U896_in = in[3];
assign _U896_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U896 (
    .in(_U896_in),
    .clk(_U896_clk),
    .out(_U896_out)
);
assign _U897_in = in[4];
assign _U897_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U897 (
    .in(_U897_in),
    .clk(_U897_clk),
    .out(_U897_out)
);
assign out[4] = _U897_out;
assign out[3] = _U896_out;
assign out[2] = _U895_out;
assign out[1] = _U894_out;
assign out[0] = _U893_out;
endmodule

module array_delay_U885 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U886_in;
wire _U886_clk;
wire [15:0] _U886_out;
wire [15:0] _U887_in;
wire _U887_clk;
wire [15:0] _U887_out;
wire [15:0] _U888_in;
wire _U888_clk;
wire [15:0] _U888_out;
wire [15:0] _U889_in;
wire _U889_clk;
wire [15:0] _U889_out;
wire [15:0] _U890_in;
wire _U890_clk;
wire [15:0] _U890_out;
assign _U886_in = in[0];
assign _U886_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U886 (
    .in(_U886_in),
    .clk(_U886_clk),
    .out(_U886_out)
);
assign _U887_in = in[1];
assign _U887_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U887 (
    .in(_U887_in),
    .clk(_U887_clk),
    .out(_U887_out)
);
assign _U888_in = in[2];
assign _U888_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U888 (
    .in(_U888_in),
    .clk(_U888_clk),
    .out(_U888_out)
);
assign _U889_in = in[3];
assign _U889_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U889 (
    .in(_U889_in),
    .clk(_U889_clk),
    .out(_U889_out)
);
assign _U890_in = in[4];
assign _U890_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U890 (
    .in(_U890_in),
    .clk(_U890_clk),
    .out(_U890_out)
);
assign out[4] = _U890_out;
assign out[3] = _U889_out;
assign out[2] = _U888_out;
assign out[1] = _U887_out;
assign out[0] = _U886_out;
endmodule

module array_delay_U878 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U879_in;
wire _U879_clk;
wire [15:0] _U879_out;
wire [15:0] _U880_in;
wire _U880_clk;
wire [15:0] _U880_out;
wire [15:0] _U881_in;
wire _U881_clk;
wire [15:0] _U881_out;
wire [15:0] _U882_in;
wire _U882_clk;
wire [15:0] _U882_out;
wire [15:0] _U883_in;
wire _U883_clk;
wire [15:0] _U883_out;
assign _U879_in = in[0];
assign _U879_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U879 (
    .in(_U879_in),
    .clk(_U879_clk),
    .out(_U879_out)
);
assign _U880_in = in[1];
assign _U880_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U880 (
    .in(_U880_in),
    .clk(_U880_clk),
    .out(_U880_out)
);
assign _U881_in = in[2];
assign _U881_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U881 (
    .in(_U881_in),
    .clk(_U881_clk),
    .out(_U881_out)
);
assign _U882_in = in[3];
assign _U882_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U882 (
    .in(_U882_in),
    .clk(_U882_clk),
    .out(_U882_out)
);
assign _U883_in = in[4];
assign _U883_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U883 (
    .in(_U883_in),
    .clk(_U883_clk),
    .out(_U883_out)
);
assign out[4] = _U883_out;
assign out[3] = _U882_out;
assign out[2] = _U881_out;
assign out[1] = _U880_out;
assign out[0] = _U879_out;
endmodule

module array_delay_U871 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U872_in;
wire _U872_clk;
wire [15:0] _U872_out;
wire [15:0] _U873_in;
wire _U873_clk;
wire [15:0] _U873_out;
wire [15:0] _U874_in;
wire _U874_clk;
wire [15:0] _U874_out;
wire [15:0] _U875_in;
wire _U875_clk;
wire [15:0] _U875_out;
wire [15:0] _U876_in;
wire _U876_clk;
wire [15:0] _U876_out;
assign _U872_in = in[0];
assign _U872_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U872 (
    .in(_U872_in),
    .clk(_U872_clk),
    .out(_U872_out)
);
assign _U873_in = in[1];
assign _U873_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U873 (
    .in(_U873_in),
    .clk(_U873_clk),
    .out(_U873_out)
);
assign _U874_in = in[2];
assign _U874_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U874 (
    .in(_U874_in),
    .clk(_U874_clk),
    .out(_U874_out)
);
assign _U875_in = in[3];
assign _U875_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U875 (
    .in(_U875_in),
    .clk(_U875_clk),
    .out(_U875_out)
);
assign _U876_in = in[4];
assign _U876_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U876 (
    .in(_U876_in),
    .clk(_U876_clk),
    .out(_U876_out)
);
assign out[4] = _U876_out;
assign out[3] = _U875_out;
assign out[2] = _U874_out;
assign out[1] = _U873_out;
assign out[0] = _U872_out;
endmodule

module array_delay_U864 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U865_in;
wire _U865_clk;
wire [15:0] _U865_out;
wire [15:0] _U866_in;
wire _U866_clk;
wire [15:0] _U866_out;
wire [15:0] _U867_in;
wire _U867_clk;
wire [15:0] _U867_out;
wire [15:0] _U868_in;
wire _U868_clk;
wire [15:0] _U868_out;
wire [15:0] _U869_in;
wire _U869_clk;
wire [15:0] _U869_out;
assign _U865_in = in[0];
assign _U865_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U865 (
    .in(_U865_in),
    .clk(_U865_clk),
    .out(_U865_out)
);
assign _U866_in = in[1];
assign _U866_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U866 (
    .in(_U866_in),
    .clk(_U866_clk),
    .out(_U866_out)
);
assign _U867_in = in[2];
assign _U867_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U867 (
    .in(_U867_in),
    .clk(_U867_clk),
    .out(_U867_out)
);
assign _U868_in = in[3];
assign _U868_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U868 (
    .in(_U868_in),
    .clk(_U868_clk),
    .out(_U868_out)
);
assign _U869_in = in[4];
assign _U869_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U869 (
    .in(_U869_in),
    .clk(_U869_clk),
    .out(_U869_out)
);
assign out[4] = _U869_out;
assign out[3] = _U868_out;
assign out[2] = _U867_out;
assign out[1] = _U866_out;
assign out[0] = _U865_out;
endmodule

module array_delay_U857 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U858_in;
wire _U858_clk;
wire [15:0] _U858_out;
wire [15:0] _U859_in;
wire _U859_clk;
wire [15:0] _U859_out;
wire [15:0] _U860_in;
wire _U860_clk;
wire [15:0] _U860_out;
wire [15:0] _U861_in;
wire _U861_clk;
wire [15:0] _U861_out;
wire [15:0] _U862_in;
wire _U862_clk;
wire [15:0] _U862_out;
assign _U858_in = in[0];
assign _U858_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U858 (
    .in(_U858_in),
    .clk(_U858_clk),
    .out(_U858_out)
);
assign _U859_in = in[1];
assign _U859_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U859 (
    .in(_U859_in),
    .clk(_U859_clk),
    .out(_U859_out)
);
assign _U860_in = in[2];
assign _U860_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U860 (
    .in(_U860_in),
    .clk(_U860_clk),
    .out(_U860_out)
);
assign _U861_in = in[3];
assign _U861_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U861 (
    .in(_U861_in),
    .clk(_U861_clk),
    .out(_U861_out)
);
assign _U862_in = in[4];
assign _U862_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U862 (
    .in(_U862_in),
    .clk(_U862_clk),
    .out(_U862_out)
);
assign out[4] = _U862_out;
assign out[3] = _U861_out;
assign out[2] = _U860_out;
assign out[1] = _U859_out;
assign out[0] = _U858_out;
endmodule

module array_delay_U850 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U851_in;
wire _U851_clk;
wire [15:0] _U851_out;
wire [15:0] _U852_in;
wire _U852_clk;
wire [15:0] _U852_out;
wire [15:0] _U853_in;
wire _U853_clk;
wire [15:0] _U853_out;
wire [15:0] _U854_in;
wire _U854_clk;
wire [15:0] _U854_out;
wire [15:0] _U855_in;
wire _U855_clk;
wire [15:0] _U855_out;
assign _U851_in = in[0];
assign _U851_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U851 (
    .in(_U851_in),
    .clk(_U851_clk),
    .out(_U851_out)
);
assign _U852_in = in[1];
assign _U852_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U852 (
    .in(_U852_in),
    .clk(_U852_clk),
    .out(_U852_out)
);
assign _U853_in = in[2];
assign _U853_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U853 (
    .in(_U853_in),
    .clk(_U853_clk),
    .out(_U853_out)
);
assign _U854_in = in[3];
assign _U854_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U854 (
    .in(_U854_in),
    .clk(_U854_clk),
    .out(_U854_out)
);
assign _U855_in = in[4];
assign _U855_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U855 (
    .in(_U855_in),
    .clk(_U855_clk),
    .out(_U855_out)
);
assign out[4] = _U855_out;
assign out[3] = _U854_out;
assign out[2] = _U853_out;
assign out[1] = _U852_out;
assign out[0] = _U851_out;
endmodule

module array_delay_U824 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U825_in;
wire _U825_clk;
wire [15:0] _U825_out;
wire [15:0] _U826_in;
wire _U826_clk;
wire [15:0] _U826_out;
wire [15:0] _U827_in;
wire _U827_clk;
wire [15:0] _U827_out;
wire [15:0] _U828_in;
wire _U828_clk;
wire [15:0] _U828_out;
wire [15:0] _U829_in;
wire _U829_clk;
wire [15:0] _U829_out;
assign _U825_in = in[0];
assign _U825_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U825 (
    .in(_U825_in),
    .clk(_U825_clk),
    .out(_U825_out)
);
assign _U826_in = in[1];
assign _U826_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U826 (
    .in(_U826_in),
    .clk(_U826_clk),
    .out(_U826_out)
);
assign _U827_in = in[2];
assign _U827_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U827 (
    .in(_U827_in),
    .clk(_U827_clk),
    .out(_U827_out)
);
assign _U828_in = in[3];
assign _U828_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U828 (
    .in(_U828_in),
    .clk(_U828_clk),
    .out(_U828_out)
);
assign _U829_in = in[4];
assign _U829_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U829 (
    .in(_U829_in),
    .clk(_U829_clk),
    .out(_U829_out)
);
assign out[4] = _U829_out;
assign out[3] = _U828_out;
assign out[2] = _U827_out;
assign out[1] = _U826_out;
assign out[0] = _U825_out;
endmodule

module array_delay_U817 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U818_in;
wire _U818_clk;
wire [15:0] _U818_out;
wire [15:0] _U819_in;
wire _U819_clk;
wire [15:0] _U819_out;
wire [15:0] _U820_in;
wire _U820_clk;
wire [15:0] _U820_out;
wire [15:0] _U821_in;
wire _U821_clk;
wire [15:0] _U821_out;
wire [15:0] _U822_in;
wire _U822_clk;
wire [15:0] _U822_out;
assign _U818_in = in[0];
assign _U818_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U818 (
    .in(_U818_in),
    .clk(_U818_clk),
    .out(_U818_out)
);
assign _U819_in = in[1];
assign _U819_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U819 (
    .in(_U819_in),
    .clk(_U819_clk),
    .out(_U819_out)
);
assign _U820_in = in[2];
assign _U820_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U820 (
    .in(_U820_in),
    .clk(_U820_clk),
    .out(_U820_out)
);
assign _U821_in = in[3];
assign _U821_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U821 (
    .in(_U821_in),
    .clk(_U821_clk),
    .out(_U821_out)
);
assign _U822_in = in[4];
assign _U822_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U822 (
    .in(_U822_in),
    .clk(_U822_clk),
    .out(_U822_out)
);
assign out[4] = _U822_out;
assign out[3] = _U821_out;
assign out[2] = _U820_out;
assign out[1] = _U819_out;
assign out[0] = _U818_out;
endmodule

module array_delay_U774 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U775_in;
wire _U775_clk;
wire [15:0] _U775_out;
wire [15:0] _U776_in;
wire _U776_clk;
wire [15:0] _U776_out;
wire [15:0] _U777_in;
wire _U777_clk;
wire [15:0] _U777_out;
wire [15:0] _U778_in;
wire _U778_clk;
wire [15:0] _U778_out;
wire [15:0] _U779_in;
wire _U779_clk;
wire [15:0] _U779_out;
assign _U775_in = in[0];
assign _U775_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U775 (
    .in(_U775_in),
    .clk(_U775_clk),
    .out(_U775_out)
);
assign _U776_in = in[1];
assign _U776_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U776 (
    .in(_U776_in),
    .clk(_U776_clk),
    .out(_U776_out)
);
assign _U777_in = in[2];
assign _U777_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U777 (
    .in(_U777_in),
    .clk(_U777_clk),
    .out(_U777_out)
);
assign _U778_in = in[3];
assign _U778_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U778 (
    .in(_U778_in),
    .clk(_U778_clk),
    .out(_U778_out)
);
assign _U779_in = in[4];
assign _U779_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U779 (
    .in(_U779_in),
    .clk(_U779_clk),
    .out(_U779_out)
);
assign out[4] = _U779_out;
assign out[3] = _U778_out;
assign out[2] = _U777_out;
assign out[1] = _U776_out;
assign out[0] = _U775_out;
endmodule

module array_delay_U767 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U768_in;
wire _U768_clk;
wire [15:0] _U768_out;
wire [15:0] _U769_in;
wire _U769_clk;
wire [15:0] _U769_out;
wire [15:0] _U770_in;
wire _U770_clk;
wire [15:0] _U770_out;
wire [15:0] _U771_in;
wire _U771_clk;
wire [15:0] _U771_out;
wire [15:0] _U772_in;
wire _U772_clk;
wire [15:0] _U772_out;
assign _U768_in = in[0];
assign _U768_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U768 (
    .in(_U768_in),
    .clk(_U768_clk),
    .out(_U768_out)
);
assign _U769_in = in[1];
assign _U769_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U769 (
    .in(_U769_in),
    .clk(_U769_clk),
    .out(_U769_out)
);
assign _U770_in = in[2];
assign _U770_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U770 (
    .in(_U770_in),
    .clk(_U770_clk),
    .out(_U770_out)
);
assign _U771_in = in[3];
assign _U771_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U771 (
    .in(_U771_in),
    .clk(_U771_clk),
    .out(_U771_out)
);
assign _U772_in = in[4];
assign _U772_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U772 (
    .in(_U772_in),
    .clk(_U772_clk),
    .out(_U772_out)
);
assign out[4] = _U772_out;
assign out[3] = _U771_out;
assign out[2] = _U770_out;
assign out[1] = _U769_out;
assign out[0] = _U768_out;
endmodule

module array_delay_U760 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U761_in;
wire _U761_clk;
wire [15:0] _U761_out;
wire [15:0] _U762_in;
wire _U762_clk;
wire [15:0] _U762_out;
wire [15:0] _U763_in;
wire _U763_clk;
wire [15:0] _U763_out;
wire [15:0] _U764_in;
wire _U764_clk;
wire [15:0] _U764_out;
wire [15:0] _U765_in;
wire _U765_clk;
wire [15:0] _U765_out;
assign _U761_in = in[0];
assign _U761_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U761 (
    .in(_U761_in),
    .clk(_U761_clk),
    .out(_U761_out)
);
assign _U762_in = in[1];
assign _U762_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U762 (
    .in(_U762_in),
    .clk(_U762_clk),
    .out(_U762_out)
);
assign _U763_in = in[2];
assign _U763_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U763 (
    .in(_U763_in),
    .clk(_U763_clk),
    .out(_U763_out)
);
assign _U764_in = in[3];
assign _U764_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U764 (
    .in(_U764_in),
    .clk(_U764_clk),
    .out(_U764_out)
);
assign _U765_in = in[4];
assign _U765_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U765 (
    .in(_U765_in),
    .clk(_U765_clk),
    .out(_U765_out)
);
assign out[4] = _U765_out;
assign out[3] = _U764_out;
assign out[2] = _U763_out;
assign out[1] = _U762_out;
assign out[0] = _U761_out;
endmodule

module array_delay_U753 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U754_in;
wire _U754_clk;
wire [15:0] _U754_out;
wire [15:0] _U755_in;
wire _U755_clk;
wire [15:0] _U755_out;
wire [15:0] _U756_in;
wire _U756_clk;
wire [15:0] _U756_out;
wire [15:0] _U757_in;
wire _U757_clk;
wire [15:0] _U757_out;
wire [15:0] _U758_in;
wire _U758_clk;
wire [15:0] _U758_out;
assign _U754_in = in[0];
assign _U754_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U754 (
    .in(_U754_in),
    .clk(_U754_clk),
    .out(_U754_out)
);
assign _U755_in = in[1];
assign _U755_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U755 (
    .in(_U755_in),
    .clk(_U755_clk),
    .out(_U755_out)
);
assign _U756_in = in[2];
assign _U756_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U756 (
    .in(_U756_in),
    .clk(_U756_clk),
    .out(_U756_out)
);
assign _U757_in = in[3];
assign _U757_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U757 (
    .in(_U757_in),
    .clk(_U757_clk),
    .out(_U757_out)
);
assign _U758_in = in[4];
assign _U758_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U758 (
    .in(_U758_in),
    .clk(_U758_clk),
    .out(_U758_out)
);
assign out[4] = _U758_out;
assign out[3] = _U757_out;
assign out[2] = _U756_out;
assign out[1] = _U755_out;
assign out[0] = _U754_out;
endmodule

module array_delay_U746 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U747_in;
wire _U747_clk;
wire [15:0] _U747_out;
wire [15:0] _U748_in;
wire _U748_clk;
wire [15:0] _U748_out;
wire [15:0] _U749_in;
wire _U749_clk;
wire [15:0] _U749_out;
wire [15:0] _U750_in;
wire _U750_clk;
wire [15:0] _U750_out;
wire [15:0] _U751_in;
wire _U751_clk;
wire [15:0] _U751_out;
assign _U747_in = in[0];
assign _U747_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U747 (
    .in(_U747_in),
    .clk(_U747_clk),
    .out(_U747_out)
);
assign _U748_in = in[1];
assign _U748_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U748 (
    .in(_U748_in),
    .clk(_U748_clk),
    .out(_U748_out)
);
assign _U749_in = in[2];
assign _U749_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U749 (
    .in(_U749_in),
    .clk(_U749_clk),
    .out(_U749_out)
);
assign _U750_in = in[3];
assign _U750_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U750 (
    .in(_U750_in),
    .clk(_U750_clk),
    .out(_U750_out)
);
assign _U751_in = in[4];
assign _U751_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U751 (
    .in(_U751_in),
    .clk(_U751_clk),
    .out(_U751_out)
);
assign out[4] = _U751_out;
assign out[3] = _U750_out;
assign out[2] = _U749_out;
assign out[1] = _U748_out;
assign out[0] = _U747_out;
endmodule

module array_delay_U739 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U740_in;
wire _U740_clk;
wire [15:0] _U740_out;
wire [15:0] _U741_in;
wire _U741_clk;
wire [15:0] _U741_out;
wire [15:0] _U742_in;
wire _U742_clk;
wire [15:0] _U742_out;
wire [15:0] _U743_in;
wire _U743_clk;
wire [15:0] _U743_out;
wire [15:0] _U744_in;
wire _U744_clk;
wire [15:0] _U744_out;
assign _U740_in = in[0];
assign _U740_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U740 (
    .in(_U740_in),
    .clk(_U740_clk),
    .out(_U740_out)
);
assign _U741_in = in[1];
assign _U741_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U741 (
    .in(_U741_in),
    .clk(_U741_clk),
    .out(_U741_out)
);
assign _U742_in = in[2];
assign _U742_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U742 (
    .in(_U742_in),
    .clk(_U742_clk),
    .out(_U742_out)
);
assign _U743_in = in[3];
assign _U743_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U743 (
    .in(_U743_in),
    .clk(_U743_clk),
    .out(_U743_out)
);
assign _U744_in = in[4];
assign _U744_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U744 (
    .in(_U744_in),
    .clk(_U744_clk),
    .out(_U744_out)
);
assign out[4] = _U744_out;
assign out[3] = _U743_out;
assign out[2] = _U742_out;
assign out[1] = _U741_out;
assign out[0] = _U740_out;
endmodule

module array_delay_U732 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U733_in;
wire _U733_clk;
wire [15:0] _U733_out;
wire [15:0] _U734_in;
wire _U734_clk;
wire [15:0] _U734_out;
wire [15:0] _U735_in;
wire _U735_clk;
wire [15:0] _U735_out;
wire [15:0] _U736_in;
wire _U736_clk;
wire [15:0] _U736_out;
wire [15:0] _U737_in;
wire _U737_clk;
wire [15:0] _U737_out;
assign _U733_in = in[0];
assign _U733_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U733 (
    .in(_U733_in),
    .clk(_U733_clk),
    .out(_U733_out)
);
assign _U734_in = in[1];
assign _U734_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U734 (
    .in(_U734_in),
    .clk(_U734_clk),
    .out(_U734_out)
);
assign _U735_in = in[2];
assign _U735_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U735 (
    .in(_U735_in),
    .clk(_U735_clk),
    .out(_U735_out)
);
assign _U736_in = in[3];
assign _U736_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U736 (
    .in(_U736_in),
    .clk(_U736_clk),
    .out(_U736_out)
);
assign _U737_in = in[4];
assign _U737_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U737 (
    .in(_U737_in),
    .clk(_U737_clk),
    .out(_U737_out)
);
assign out[4] = _U737_out;
assign out[3] = _U736_out;
assign out[2] = _U735_out;
assign out[1] = _U734_out;
assign out[0] = _U733_out;
endmodule

module array_delay_U725 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U726_in;
wire _U726_clk;
wire [15:0] _U726_out;
wire [15:0] _U727_in;
wire _U727_clk;
wire [15:0] _U727_out;
wire [15:0] _U728_in;
wire _U728_clk;
wire [15:0] _U728_out;
wire [15:0] _U729_in;
wire _U729_clk;
wire [15:0] _U729_out;
wire [15:0] _U730_in;
wire _U730_clk;
wire [15:0] _U730_out;
assign _U726_in = in[0];
assign _U726_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U726 (
    .in(_U726_in),
    .clk(_U726_clk),
    .out(_U726_out)
);
assign _U727_in = in[1];
assign _U727_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U727 (
    .in(_U727_in),
    .clk(_U727_clk),
    .out(_U727_out)
);
assign _U728_in = in[2];
assign _U728_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U728 (
    .in(_U728_in),
    .clk(_U728_clk),
    .out(_U728_out)
);
assign _U729_in = in[3];
assign _U729_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U729 (
    .in(_U729_in),
    .clk(_U729_clk),
    .out(_U729_out)
);
assign _U730_in = in[4];
assign _U730_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U730 (
    .in(_U730_in),
    .clk(_U730_clk),
    .out(_U730_out)
);
assign out[4] = _U730_out;
assign out[3] = _U729_out;
assign out[2] = _U728_out;
assign out[1] = _U727_out;
assign out[0] = _U726_out;
endmodule

module array_delay_U718 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U719_in;
wire _U719_clk;
wire [15:0] _U719_out;
wire [15:0] _U720_in;
wire _U720_clk;
wire [15:0] _U720_out;
wire [15:0] _U721_in;
wire _U721_clk;
wire [15:0] _U721_out;
wire [15:0] _U722_in;
wire _U722_clk;
wire [15:0] _U722_out;
wire [15:0] _U723_in;
wire _U723_clk;
wire [15:0] _U723_out;
assign _U719_in = in[0];
assign _U719_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U719 (
    .in(_U719_in),
    .clk(_U719_clk),
    .out(_U719_out)
);
assign _U720_in = in[1];
assign _U720_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U720 (
    .in(_U720_in),
    .clk(_U720_clk),
    .out(_U720_out)
);
assign _U721_in = in[2];
assign _U721_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U721 (
    .in(_U721_in),
    .clk(_U721_clk),
    .out(_U721_out)
);
assign _U722_in = in[3];
assign _U722_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U722 (
    .in(_U722_in),
    .clk(_U722_clk),
    .out(_U722_out)
);
assign _U723_in = in[4];
assign _U723_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U723 (
    .in(_U723_in),
    .clk(_U723_clk),
    .out(_U723_out)
);
assign out[4] = _U723_out;
assign out[3] = _U722_out;
assign out[2] = _U721_out;
assign out[1] = _U720_out;
assign out[0] = _U719_out;
endmodule

module array_delay_U711 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U712_in;
wire _U712_clk;
wire [15:0] _U712_out;
wire [15:0] _U713_in;
wire _U713_clk;
wire [15:0] _U713_out;
wire [15:0] _U714_in;
wire _U714_clk;
wire [15:0] _U714_out;
wire [15:0] _U715_in;
wire _U715_clk;
wire [15:0] _U715_out;
wire [15:0] _U716_in;
wire _U716_clk;
wire [15:0] _U716_out;
assign _U712_in = in[0];
assign _U712_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U712 (
    .in(_U712_in),
    .clk(_U712_clk),
    .out(_U712_out)
);
assign _U713_in = in[1];
assign _U713_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U713 (
    .in(_U713_in),
    .clk(_U713_clk),
    .out(_U713_out)
);
assign _U714_in = in[2];
assign _U714_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U714 (
    .in(_U714_in),
    .clk(_U714_clk),
    .out(_U714_out)
);
assign _U715_in = in[3];
assign _U715_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U715 (
    .in(_U715_in),
    .clk(_U715_clk),
    .out(_U715_out)
);
assign _U716_in = in[4];
assign _U716_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U716 (
    .in(_U716_in),
    .clk(_U716_clk),
    .out(_U716_out)
);
assign out[4] = _U716_out;
assign out[3] = _U715_out;
assign out[2] = _U714_out;
assign out[1] = _U713_out;
assign out[0] = _U712_out;
endmodule

module array_delay_U704 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U705_in;
wire _U705_clk;
wire [15:0] _U705_out;
wire [15:0] _U706_in;
wire _U706_clk;
wire [15:0] _U706_out;
wire [15:0] _U707_in;
wire _U707_clk;
wire [15:0] _U707_out;
wire [15:0] _U708_in;
wire _U708_clk;
wire [15:0] _U708_out;
wire [15:0] _U709_in;
wire _U709_clk;
wire [15:0] _U709_out;
assign _U705_in = in[0];
assign _U705_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U705 (
    .in(_U705_in),
    .clk(_U705_clk),
    .out(_U705_out)
);
assign _U706_in = in[1];
assign _U706_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U706 (
    .in(_U706_in),
    .clk(_U706_clk),
    .out(_U706_out)
);
assign _U707_in = in[2];
assign _U707_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U707 (
    .in(_U707_in),
    .clk(_U707_clk),
    .out(_U707_out)
);
assign _U708_in = in[3];
assign _U708_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U708 (
    .in(_U708_in),
    .clk(_U708_clk),
    .out(_U708_out)
);
assign _U709_in = in[4];
assign _U709_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U709 (
    .in(_U709_in),
    .clk(_U709_clk),
    .out(_U709_out)
);
assign out[4] = _U709_out;
assign out[3] = _U708_out;
assign out[2] = _U707_out;
assign out[1] = _U706_out;
assign out[0] = _U705_out;
endmodule

module array_delay_U697 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U698_in;
wire _U698_clk;
wire [15:0] _U698_out;
wire [15:0] _U699_in;
wire _U699_clk;
wire [15:0] _U699_out;
wire [15:0] _U700_in;
wire _U700_clk;
wire [15:0] _U700_out;
wire [15:0] _U701_in;
wire _U701_clk;
wire [15:0] _U701_out;
wire [15:0] _U702_in;
wire _U702_clk;
wire [15:0] _U702_out;
assign _U698_in = in[0];
assign _U698_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U698 (
    .in(_U698_in),
    .clk(_U698_clk),
    .out(_U698_out)
);
assign _U699_in = in[1];
assign _U699_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U699 (
    .in(_U699_in),
    .clk(_U699_clk),
    .out(_U699_out)
);
assign _U700_in = in[2];
assign _U700_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U700 (
    .in(_U700_in),
    .clk(_U700_clk),
    .out(_U700_out)
);
assign _U701_in = in[3];
assign _U701_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U701 (
    .in(_U701_in),
    .clk(_U701_clk),
    .out(_U701_out)
);
assign _U702_in = in[4];
assign _U702_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U702 (
    .in(_U702_in),
    .clk(_U702_clk),
    .out(_U702_out)
);
assign out[4] = _U702_out;
assign out[3] = _U701_out;
assign out[2] = _U700_out;
assign out[1] = _U699_out;
assign out[0] = _U698_out;
endmodule

module array_delay_U690 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U691_in;
wire _U691_clk;
wire [15:0] _U691_out;
wire [15:0] _U692_in;
wire _U692_clk;
wire [15:0] _U692_out;
wire [15:0] _U693_in;
wire _U693_clk;
wire [15:0] _U693_out;
wire [15:0] _U694_in;
wire _U694_clk;
wire [15:0] _U694_out;
wire [15:0] _U695_in;
wire _U695_clk;
wire [15:0] _U695_out;
assign _U691_in = in[0];
assign _U691_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U691 (
    .in(_U691_in),
    .clk(_U691_clk),
    .out(_U691_out)
);
assign _U692_in = in[1];
assign _U692_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U692 (
    .in(_U692_in),
    .clk(_U692_clk),
    .out(_U692_out)
);
assign _U693_in = in[2];
assign _U693_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U693 (
    .in(_U693_in),
    .clk(_U693_clk),
    .out(_U693_out)
);
assign _U694_in = in[3];
assign _U694_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U694 (
    .in(_U694_in),
    .clk(_U694_clk),
    .out(_U694_out)
);
assign _U695_in = in[4];
assign _U695_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U695 (
    .in(_U695_in),
    .clk(_U695_clk),
    .out(_U695_out)
);
assign out[4] = _U695_out;
assign out[3] = _U694_out;
assign out[2] = _U693_out;
assign out[1] = _U692_out;
assign out[0] = _U691_out;
endmodule

module array_delay_U683 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U684_in;
wire _U684_clk;
wire [15:0] _U684_out;
wire [15:0] _U685_in;
wire _U685_clk;
wire [15:0] _U685_out;
wire [15:0] _U686_in;
wire _U686_clk;
wire [15:0] _U686_out;
wire [15:0] _U687_in;
wire _U687_clk;
wire [15:0] _U687_out;
wire [15:0] _U688_in;
wire _U688_clk;
wire [15:0] _U688_out;
assign _U684_in = in[0];
assign _U684_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U684 (
    .in(_U684_in),
    .clk(_U684_clk),
    .out(_U684_out)
);
assign _U685_in = in[1];
assign _U685_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U685 (
    .in(_U685_in),
    .clk(_U685_clk),
    .out(_U685_out)
);
assign _U686_in = in[2];
assign _U686_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U686 (
    .in(_U686_in),
    .clk(_U686_clk),
    .out(_U686_out)
);
assign _U687_in = in[3];
assign _U687_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U687 (
    .in(_U687_in),
    .clk(_U687_clk),
    .out(_U687_out)
);
assign _U688_in = in[4];
assign _U688_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U688 (
    .in(_U688_in),
    .clk(_U688_clk),
    .out(_U688_out)
);
assign out[4] = _U688_out;
assign out[3] = _U687_out;
assign out[2] = _U686_out;
assign out[1] = _U685_out;
assign out[0] = _U684_out;
endmodule

module array_delay_U676 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U677_in;
wire _U677_clk;
wire [15:0] _U677_out;
wire [15:0] _U678_in;
wire _U678_clk;
wire [15:0] _U678_out;
wire [15:0] _U679_in;
wire _U679_clk;
wire [15:0] _U679_out;
wire [15:0] _U680_in;
wire _U680_clk;
wire [15:0] _U680_out;
wire [15:0] _U681_in;
wire _U681_clk;
wire [15:0] _U681_out;
assign _U677_in = in[0];
assign _U677_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U677 (
    .in(_U677_in),
    .clk(_U677_clk),
    .out(_U677_out)
);
assign _U678_in = in[1];
assign _U678_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U678 (
    .in(_U678_in),
    .clk(_U678_clk),
    .out(_U678_out)
);
assign _U679_in = in[2];
assign _U679_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U679 (
    .in(_U679_in),
    .clk(_U679_clk),
    .out(_U679_out)
);
assign _U680_in = in[3];
assign _U680_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U680 (
    .in(_U680_in),
    .clk(_U680_clk),
    .out(_U680_out)
);
assign _U681_in = in[4];
assign _U681_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U681 (
    .in(_U681_in),
    .clk(_U681_clk),
    .out(_U681_out)
);
assign out[4] = _U681_out;
assign out[3] = _U680_out;
assign out[2] = _U679_out;
assign out[1] = _U678_out;
assign out[0] = _U677_out;
endmodule

module array_delay_U669 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U670_in;
wire _U670_clk;
wire [15:0] _U670_out;
wire [15:0] _U671_in;
wire _U671_clk;
wire [15:0] _U671_out;
wire [15:0] _U672_in;
wire _U672_clk;
wire [15:0] _U672_out;
wire [15:0] _U673_in;
wire _U673_clk;
wire [15:0] _U673_out;
wire [15:0] _U674_in;
wire _U674_clk;
wire [15:0] _U674_out;
assign _U670_in = in[0];
assign _U670_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U670 (
    .in(_U670_in),
    .clk(_U670_clk),
    .out(_U670_out)
);
assign _U671_in = in[1];
assign _U671_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U671 (
    .in(_U671_in),
    .clk(_U671_clk),
    .out(_U671_out)
);
assign _U672_in = in[2];
assign _U672_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U672 (
    .in(_U672_in),
    .clk(_U672_clk),
    .out(_U672_out)
);
assign _U673_in = in[3];
assign _U673_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U673 (
    .in(_U673_in),
    .clk(_U673_clk),
    .out(_U673_out)
);
assign _U674_in = in[4];
assign _U674_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U674 (
    .in(_U674_in),
    .clk(_U674_clk),
    .out(_U674_out)
);
assign out[4] = _U674_out;
assign out[3] = _U673_out;
assign out[2] = _U672_out;
assign out[1] = _U671_out;
assign out[0] = _U670_out;
endmodule

module array_delay_U662 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U663_in;
wire _U663_clk;
wire [15:0] _U663_out;
wire [15:0] _U664_in;
wire _U664_clk;
wire [15:0] _U664_out;
wire [15:0] _U665_in;
wire _U665_clk;
wire [15:0] _U665_out;
wire [15:0] _U666_in;
wire _U666_clk;
wire [15:0] _U666_out;
wire [15:0] _U667_in;
wire _U667_clk;
wire [15:0] _U667_out;
assign _U663_in = in[0];
assign _U663_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U663 (
    .in(_U663_in),
    .clk(_U663_clk),
    .out(_U663_out)
);
assign _U664_in = in[1];
assign _U664_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U664 (
    .in(_U664_in),
    .clk(_U664_clk),
    .out(_U664_out)
);
assign _U665_in = in[2];
assign _U665_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U665 (
    .in(_U665_in),
    .clk(_U665_clk),
    .out(_U665_out)
);
assign _U666_in = in[3];
assign _U666_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U666 (
    .in(_U666_in),
    .clk(_U666_clk),
    .out(_U666_out)
);
assign _U667_in = in[4];
assign _U667_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U667 (
    .in(_U667_in),
    .clk(_U667_clk),
    .out(_U667_out)
);
assign out[4] = _U667_out;
assign out[3] = _U666_out;
assign out[2] = _U665_out;
assign out[1] = _U664_out;
assign out[0] = _U663_out;
endmodule

module array_delay_U636 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U637_in;
wire _U637_clk;
wire [15:0] _U637_out;
wire [15:0] _U638_in;
wire _U638_clk;
wire [15:0] _U638_out;
wire [15:0] _U639_in;
wire _U639_clk;
wire [15:0] _U639_out;
wire [15:0] _U640_in;
wire _U640_clk;
wire [15:0] _U640_out;
wire [15:0] _U641_in;
wire _U641_clk;
wire [15:0] _U641_out;
assign _U637_in = in[0];
assign _U637_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U637 (
    .in(_U637_in),
    .clk(_U637_clk),
    .out(_U637_out)
);
assign _U638_in = in[1];
assign _U638_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U638 (
    .in(_U638_in),
    .clk(_U638_clk),
    .out(_U638_out)
);
assign _U639_in = in[2];
assign _U639_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U639 (
    .in(_U639_in),
    .clk(_U639_clk),
    .out(_U639_out)
);
assign _U640_in = in[3];
assign _U640_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U640 (
    .in(_U640_in),
    .clk(_U640_clk),
    .out(_U640_out)
);
assign _U641_in = in[4];
assign _U641_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U641 (
    .in(_U641_in),
    .clk(_U641_clk),
    .out(_U641_out)
);
assign out[4] = _U641_out;
assign out[3] = _U640_out;
assign out[2] = _U639_out;
assign out[1] = _U638_out;
assign out[0] = _U637_out;
endmodule

module array_delay_U629 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U630_in;
wire _U630_clk;
wire [15:0] _U630_out;
wire [15:0] _U631_in;
wire _U631_clk;
wire [15:0] _U631_out;
wire [15:0] _U632_in;
wire _U632_clk;
wire [15:0] _U632_out;
wire [15:0] _U633_in;
wire _U633_clk;
wire [15:0] _U633_out;
wire [15:0] _U634_in;
wire _U634_clk;
wire [15:0] _U634_out;
assign _U630_in = in[0];
assign _U630_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U630 (
    .in(_U630_in),
    .clk(_U630_clk),
    .out(_U630_out)
);
assign _U631_in = in[1];
assign _U631_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U631 (
    .in(_U631_in),
    .clk(_U631_clk),
    .out(_U631_out)
);
assign _U632_in = in[2];
assign _U632_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U632 (
    .in(_U632_in),
    .clk(_U632_clk),
    .out(_U632_out)
);
assign _U633_in = in[3];
assign _U633_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U633 (
    .in(_U633_in),
    .clk(_U633_clk),
    .out(_U633_out)
);
assign _U634_in = in[4];
assign _U634_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U634 (
    .in(_U634_in),
    .clk(_U634_clk),
    .out(_U634_out)
);
assign out[4] = _U634_out;
assign out[3] = _U633_out;
assign out[2] = _U632_out;
assign out[1] = _U631_out;
assign out[0] = _U630_out;
endmodule

module array_delay_U586 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U587_in;
wire _U587_clk;
wire [15:0] _U587_out;
wire [15:0] _U588_in;
wire _U588_clk;
wire [15:0] _U588_out;
wire [15:0] _U589_in;
wire _U589_clk;
wire [15:0] _U589_out;
wire [15:0] _U590_in;
wire _U590_clk;
wire [15:0] _U590_out;
wire [15:0] _U591_in;
wire _U591_clk;
wire [15:0] _U591_out;
assign _U587_in = in[0];
assign _U587_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U587 (
    .in(_U587_in),
    .clk(_U587_clk),
    .out(_U587_out)
);
assign _U588_in = in[1];
assign _U588_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U588 (
    .in(_U588_in),
    .clk(_U588_clk),
    .out(_U588_out)
);
assign _U589_in = in[2];
assign _U589_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U589 (
    .in(_U589_in),
    .clk(_U589_clk),
    .out(_U589_out)
);
assign _U590_in = in[3];
assign _U590_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U590 (
    .in(_U590_in),
    .clk(_U590_clk),
    .out(_U590_out)
);
assign _U591_in = in[4];
assign _U591_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U591 (
    .in(_U591_in),
    .clk(_U591_clk),
    .out(_U591_out)
);
assign out[4] = _U591_out;
assign out[3] = _U590_out;
assign out[2] = _U589_out;
assign out[1] = _U588_out;
assign out[0] = _U587_out;
endmodule

module array_delay_U579 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U580_in;
wire _U580_clk;
wire [15:0] _U580_out;
wire [15:0] _U581_in;
wire _U581_clk;
wire [15:0] _U581_out;
wire [15:0] _U582_in;
wire _U582_clk;
wire [15:0] _U582_out;
wire [15:0] _U583_in;
wire _U583_clk;
wire [15:0] _U583_out;
wire [15:0] _U584_in;
wire _U584_clk;
wire [15:0] _U584_out;
assign _U580_in = in[0];
assign _U580_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U580 (
    .in(_U580_in),
    .clk(_U580_clk),
    .out(_U580_out)
);
assign _U581_in = in[1];
assign _U581_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U581 (
    .in(_U581_in),
    .clk(_U581_clk),
    .out(_U581_out)
);
assign _U582_in = in[2];
assign _U582_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U582 (
    .in(_U582_in),
    .clk(_U582_clk),
    .out(_U582_out)
);
assign _U583_in = in[3];
assign _U583_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U583 (
    .in(_U583_in),
    .clk(_U583_clk),
    .out(_U583_out)
);
assign _U584_in = in[4];
assign _U584_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U584 (
    .in(_U584_in),
    .clk(_U584_clk),
    .out(_U584_out)
);
assign out[4] = _U584_out;
assign out[3] = _U583_out;
assign out[2] = _U582_out;
assign out[1] = _U581_out;
assign out[0] = _U580_out;
endmodule

module array_delay_U572 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U573_in;
wire _U573_clk;
wire [15:0] _U573_out;
wire [15:0] _U574_in;
wire _U574_clk;
wire [15:0] _U574_out;
wire [15:0] _U575_in;
wire _U575_clk;
wire [15:0] _U575_out;
wire [15:0] _U576_in;
wire _U576_clk;
wire [15:0] _U576_out;
wire [15:0] _U577_in;
wire _U577_clk;
wire [15:0] _U577_out;
assign _U573_in = in[0];
assign _U573_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U573 (
    .in(_U573_in),
    .clk(_U573_clk),
    .out(_U573_out)
);
assign _U574_in = in[1];
assign _U574_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U574 (
    .in(_U574_in),
    .clk(_U574_clk),
    .out(_U574_out)
);
assign _U575_in = in[2];
assign _U575_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U575 (
    .in(_U575_in),
    .clk(_U575_clk),
    .out(_U575_out)
);
assign _U576_in = in[3];
assign _U576_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U576 (
    .in(_U576_in),
    .clk(_U576_clk),
    .out(_U576_out)
);
assign _U577_in = in[4];
assign _U577_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U577 (
    .in(_U577_in),
    .clk(_U577_clk),
    .out(_U577_out)
);
assign out[4] = _U577_out;
assign out[3] = _U576_out;
assign out[2] = _U575_out;
assign out[1] = _U574_out;
assign out[0] = _U573_out;
endmodule

module array_delay_U565 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U566_in;
wire _U566_clk;
wire [15:0] _U566_out;
wire [15:0] _U567_in;
wire _U567_clk;
wire [15:0] _U567_out;
wire [15:0] _U568_in;
wire _U568_clk;
wire [15:0] _U568_out;
wire [15:0] _U569_in;
wire _U569_clk;
wire [15:0] _U569_out;
wire [15:0] _U570_in;
wire _U570_clk;
wire [15:0] _U570_out;
assign _U566_in = in[0];
assign _U566_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U566 (
    .in(_U566_in),
    .clk(_U566_clk),
    .out(_U566_out)
);
assign _U567_in = in[1];
assign _U567_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U567 (
    .in(_U567_in),
    .clk(_U567_clk),
    .out(_U567_out)
);
assign _U568_in = in[2];
assign _U568_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U568 (
    .in(_U568_in),
    .clk(_U568_clk),
    .out(_U568_out)
);
assign _U569_in = in[3];
assign _U569_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U569 (
    .in(_U569_in),
    .clk(_U569_clk),
    .out(_U569_out)
);
assign _U570_in = in[4];
assign _U570_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U570 (
    .in(_U570_in),
    .clk(_U570_clk),
    .out(_U570_out)
);
assign out[4] = _U570_out;
assign out[3] = _U569_out;
assign out[2] = _U568_out;
assign out[1] = _U567_out;
assign out[0] = _U566_out;
endmodule

module array_delay_U558 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U559_in;
wire _U559_clk;
wire [15:0] _U559_out;
wire [15:0] _U560_in;
wire _U560_clk;
wire [15:0] _U560_out;
wire [15:0] _U561_in;
wire _U561_clk;
wire [15:0] _U561_out;
wire [15:0] _U562_in;
wire _U562_clk;
wire [15:0] _U562_out;
wire [15:0] _U563_in;
wire _U563_clk;
wire [15:0] _U563_out;
assign _U559_in = in[0];
assign _U559_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U559 (
    .in(_U559_in),
    .clk(_U559_clk),
    .out(_U559_out)
);
assign _U560_in = in[1];
assign _U560_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U560 (
    .in(_U560_in),
    .clk(_U560_clk),
    .out(_U560_out)
);
assign _U561_in = in[2];
assign _U561_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U561 (
    .in(_U561_in),
    .clk(_U561_clk),
    .out(_U561_out)
);
assign _U562_in = in[3];
assign _U562_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U562 (
    .in(_U562_in),
    .clk(_U562_clk),
    .out(_U562_out)
);
assign _U563_in = in[4];
assign _U563_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U563 (
    .in(_U563_in),
    .clk(_U563_clk),
    .out(_U563_out)
);
assign out[4] = _U563_out;
assign out[3] = _U562_out;
assign out[2] = _U561_out;
assign out[1] = _U560_out;
assign out[0] = _U559_out;
endmodule

module array_delay_U551 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U552_in;
wire _U552_clk;
wire [15:0] _U552_out;
wire [15:0] _U553_in;
wire _U553_clk;
wire [15:0] _U553_out;
wire [15:0] _U554_in;
wire _U554_clk;
wire [15:0] _U554_out;
wire [15:0] _U555_in;
wire _U555_clk;
wire [15:0] _U555_out;
wire [15:0] _U556_in;
wire _U556_clk;
wire [15:0] _U556_out;
assign _U552_in = in[0];
assign _U552_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U552 (
    .in(_U552_in),
    .clk(_U552_clk),
    .out(_U552_out)
);
assign _U553_in = in[1];
assign _U553_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U553 (
    .in(_U553_in),
    .clk(_U553_clk),
    .out(_U553_out)
);
assign _U554_in = in[2];
assign _U554_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U554 (
    .in(_U554_in),
    .clk(_U554_clk),
    .out(_U554_out)
);
assign _U555_in = in[3];
assign _U555_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U555 (
    .in(_U555_in),
    .clk(_U555_clk),
    .out(_U555_out)
);
assign _U556_in = in[4];
assign _U556_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U556 (
    .in(_U556_in),
    .clk(_U556_clk),
    .out(_U556_out)
);
assign out[4] = _U556_out;
assign out[3] = _U555_out;
assign out[2] = _U554_out;
assign out[1] = _U553_out;
assign out[0] = _U552_out;
endmodule

module array_delay_U544 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U545_in;
wire _U545_clk;
wire [15:0] _U545_out;
wire [15:0] _U546_in;
wire _U546_clk;
wire [15:0] _U546_out;
wire [15:0] _U547_in;
wire _U547_clk;
wire [15:0] _U547_out;
wire [15:0] _U548_in;
wire _U548_clk;
wire [15:0] _U548_out;
wire [15:0] _U549_in;
wire _U549_clk;
wire [15:0] _U549_out;
assign _U545_in = in[0];
assign _U545_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U545 (
    .in(_U545_in),
    .clk(_U545_clk),
    .out(_U545_out)
);
assign _U546_in = in[1];
assign _U546_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U546 (
    .in(_U546_in),
    .clk(_U546_clk),
    .out(_U546_out)
);
assign _U547_in = in[2];
assign _U547_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U547 (
    .in(_U547_in),
    .clk(_U547_clk),
    .out(_U547_out)
);
assign _U548_in = in[3];
assign _U548_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U548 (
    .in(_U548_in),
    .clk(_U548_clk),
    .out(_U548_out)
);
assign _U549_in = in[4];
assign _U549_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U549 (
    .in(_U549_in),
    .clk(_U549_clk),
    .out(_U549_out)
);
assign out[4] = _U549_out;
assign out[3] = _U548_out;
assign out[2] = _U547_out;
assign out[1] = _U546_out;
assign out[0] = _U545_out;
endmodule

module array_delay_U537 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U538_in;
wire _U538_clk;
wire [15:0] _U538_out;
wire [15:0] _U539_in;
wire _U539_clk;
wire [15:0] _U539_out;
wire [15:0] _U540_in;
wire _U540_clk;
wire [15:0] _U540_out;
wire [15:0] _U541_in;
wire _U541_clk;
wire [15:0] _U541_out;
wire [15:0] _U542_in;
wire _U542_clk;
wire [15:0] _U542_out;
assign _U538_in = in[0];
assign _U538_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U538 (
    .in(_U538_in),
    .clk(_U538_clk),
    .out(_U538_out)
);
assign _U539_in = in[1];
assign _U539_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U539 (
    .in(_U539_in),
    .clk(_U539_clk),
    .out(_U539_out)
);
assign _U540_in = in[2];
assign _U540_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U540 (
    .in(_U540_in),
    .clk(_U540_clk),
    .out(_U540_out)
);
assign _U541_in = in[3];
assign _U541_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U541 (
    .in(_U541_in),
    .clk(_U541_clk),
    .out(_U541_out)
);
assign _U542_in = in[4];
assign _U542_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U542 (
    .in(_U542_in),
    .clk(_U542_clk),
    .out(_U542_out)
);
assign out[4] = _U542_out;
assign out[3] = _U541_out;
assign out[2] = _U540_out;
assign out[1] = _U539_out;
assign out[0] = _U538_out;
endmodule

module array_delay_U530 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U531_in;
wire _U531_clk;
wire [15:0] _U531_out;
wire [15:0] _U532_in;
wire _U532_clk;
wire [15:0] _U532_out;
wire [15:0] _U533_in;
wire _U533_clk;
wire [15:0] _U533_out;
wire [15:0] _U534_in;
wire _U534_clk;
wire [15:0] _U534_out;
wire [15:0] _U535_in;
wire _U535_clk;
wire [15:0] _U535_out;
assign _U531_in = in[0];
assign _U531_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U531 (
    .in(_U531_in),
    .clk(_U531_clk),
    .out(_U531_out)
);
assign _U532_in = in[1];
assign _U532_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U532 (
    .in(_U532_in),
    .clk(_U532_clk),
    .out(_U532_out)
);
assign _U533_in = in[2];
assign _U533_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U533 (
    .in(_U533_in),
    .clk(_U533_clk),
    .out(_U533_out)
);
assign _U534_in = in[3];
assign _U534_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U534 (
    .in(_U534_in),
    .clk(_U534_clk),
    .out(_U534_out)
);
assign _U535_in = in[4];
assign _U535_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U535 (
    .in(_U535_in),
    .clk(_U535_clk),
    .out(_U535_out)
);
assign out[4] = _U535_out;
assign out[3] = _U534_out;
assign out[2] = _U533_out;
assign out[1] = _U532_out;
assign out[0] = _U531_out;
endmodule

module array_delay_U523 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U524_in;
wire _U524_clk;
wire [15:0] _U524_out;
wire [15:0] _U525_in;
wire _U525_clk;
wire [15:0] _U525_out;
wire [15:0] _U526_in;
wire _U526_clk;
wire [15:0] _U526_out;
wire [15:0] _U527_in;
wire _U527_clk;
wire [15:0] _U527_out;
wire [15:0] _U528_in;
wire _U528_clk;
wire [15:0] _U528_out;
assign _U524_in = in[0];
assign _U524_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U524 (
    .in(_U524_in),
    .clk(_U524_clk),
    .out(_U524_out)
);
assign _U525_in = in[1];
assign _U525_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U525 (
    .in(_U525_in),
    .clk(_U525_clk),
    .out(_U525_out)
);
assign _U526_in = in[2];
assign _U526_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U526 (
    .in(_U526_in),
    .clk(_U526_clk),
    .out(_U526_out)
);
assign _U527_in = in[3];
assign _U527_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U527 (
    .in(_U527_in),
    .clk(_U527_clk),
    .out(_U527_out)
);
assign _U528_in = in[4];
assign _U528_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U528 (
    .in(_U528_in),
    .clk(_U528_clk),
    .out(_U528_out)
);
assign out[4] = _U528_out;
assign out[3] = _U527_out;
assign out[2] = _U526_out;
assign out[1] = _U525_out;
assign out[0] = _U524_out;
endmodule

module array_delay_U516 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U517_in;
wire _U517_clk;
wire [15:0] _U517_out;
wire [15:0] _U518_in;
wire _U518_clk;
wire [15:0] _U518_out;
wire [15:0] _U519_in;
wire _U519_clk;
wire [15:0] _U519_out;
wire [15:0] _U520_in;
wire _U520_clk;
wire [15:0] _U520_out;
wire [15:0] _U521_in;
wire _U521_clk;
wire [15:0] _U521_out;
assign _U517_in = in[0];
assign _U517_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U517 (
    .in(_U517_in),
    .clk(_U517_clk),
    .out(_U517_out)
);
assign _U518_in = in[1];
assign _U518_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U518 (
    .in(_U518_in),
    .clk(_U518_clk),
    .out(_U518_out)
);
assign _U519_in = in[2];
assign _U519_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U519 (
    .in(_U519_in),
    .clk(_U519_clk),
    .out(_U519_out)
);
assign _U520_in = in[3];
assign _U520_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U520 (
    .in(_U520_in),
    .clk(_U520_clk),
    .out(_U520_out)
);
assign _U521_in = in[4];
assign _U521_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U521 (
    .in(_U521_in),
    .clk(_U521_clk),
    .out(_U521_out)
);
assign out[4] = _U521_out;
assign out[3] = _U520_out;
assign out[2] = _U519_out;
assign out[1] = _U518_out;
assign out[0] = _U517_out;
endmodule

module array_delay_U509 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U510_in;
wire _U510_clk;
wire [15:0] _U510_out;
wire [15:0] _U511_in;
wire _U511_clk;
wire [15:0] _U511_out;
wire [15:0] _U512_in;
wire _U512_clk;
wire [15:0] _U512_out;
wire [15:0] _U513_in;
wire _U513_clk;
wire [15:0] _U513_out;
wire [15:0] _U514_in;
wire _U514_clk;
wire [15:0] _U514_out;
assign _U510_in = in[0];
assign _U510_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U510 (
    .in(_U510_in),
    .clk(_U510_clk),
    .out(_U510_out)
);
assign _U511_in = in[1];
assign _U511_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U511 (
    .in(_U511_in),
    .clk(_U511_clk),
    .out(_U511_out)
);
assign _U512_in = in[2];
assign _U512_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U512 (
    .in(_U512_in),
    .clk(_U512_clk),
    .out(_U512_out)
);
assign _U513_in = in[3];
assign _U513_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U513 (
    .in(_U513_in),
    .clk(_U513_clk),
    .out(_U513_out)
);
assign _U514_in = in[4];
assign _U514_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U514 (
    .in(_U514_in),
    .clk(_U514_clk),
    .out(_U514_out)
);
assign out[4] = _U514_out;
assign out[3] = _U513_out;
assign out[2] = _U512_out;
assign out[1] = _U511_out;
assign out[0] = _U510_out;
endmodule

module array_delay_U502 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U503_in;
wire _U503_clk;
wire [15:0] _U503_out;
wire [15:0] _U504_in;
wire _U504_clk;
wire [15:0] _U504_out;
wire [15:0] _U505_in;
wire _U505_clk;
wire [15:0] _U505_out;
wire [15:0] _U506_in;
wire _U506_clk;
wire [15:0] _U506_out;
wire [15:0] _U507_in;
wire _U507_clk;
wire [15:0] _U507_out;
assign _U503_in = in[0];
assign _U503_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U503 (
    .in(_U503_in),
    .clk(_U503_clk),
    .out(_U503_out)
);
assign _U504_in = in[1];
assign _U504_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U504 (
    .in(_U504_in),
    .clk(_U504_clk),
    .out(_U504_out)
);
assign _U505_in = in[2];
assign _U505_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U505 (
    .in(_U505_in),
    .clk(_U505_clk),
    .out(_U505_out)
);
assign _U506_in = in[3];
assign _U506_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U506 (
    .in(_U506_in),
    .clk(_U506_clk),
    .out(_U506_out)
);
assign _U507_in = in[4];
assign _U507_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U507 (
    .in(_U507_in),
    .clk(_U507_clk),
    .out(_U507_out)
);
assign out[4] = _U507_out;
assign out[3] = _U506_out;
assign out[2] = _U505_out;
assign out[1] = _U504_out;
assign out[0] = _U503_out;
endmodule

module array_delay_U495 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U496_in;
wire _U496_clk;
wire [15:0] _U496_out;
wire [15:0] _U497_in;
wire _U497_clk;
wire [15:0] _U497_out;
wire [15:0] _U498_in;
wire _U498_clk;
wire [15:0] _U498_out;
wire [15:0] _U499_in;
wire _U499_clk;
wire [15:0] _U499_out;
wire [15:0] _U500_in;
wire _U500_clk;
wire [15:0] _U500_out;
assign _U496_in = in[0];
assign _U496_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U496 (
    .in(_U496_in),
    .clk(_U496_clk),
    .out(_U496_out)
);
assign _U497_in = in[1];
assign _U497_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U497 (
    .in(_U497_in),
    .clk(_U497_clk),
    .out(_U497_out)
);
assign _U498_in = in[2];
assign _U498_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U498 (
    .in(_U498_in),
    .clk(_U498_clk),
    .out(_U498_out)
);
assign _U499_in = in[3];
assign _U499_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U499 (
    .in(_U499_in),
    .clk(_U499_clk),
    .out(_U499_out)
);
assign _U500_in = in[4];
assign _U500_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U500 (
    .in(_U500_in),
    .clk(_U500_clk),
    .out(_U500_out)
);
assign out[4] = _U500_out;
assign out[3] = _U499_out;
assign out[2] = _U498_out;
assign out[1] = _U497_out;
assign out[0] = _U496_out;
endmodule

module array_delay_U488 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U489_in;
wire _U489_clk;
wire [15:0] _U489_out;
wire [15:0] _U490_in;
wire _U490_clk;
wire [15:0] _U490_out;
wire [15:0] _U491_in;
wire _U491_clk;
wire [15:0] _U491_out;
wire [15:0] _U492_in;
wire _U492_clk;
wire [15:0] _U492_out;
wire [15:0] _U493_in;
wire _U493_clk;
wire [15:0] _U493_out;
assign _U489_in = in[0];
assign _U489_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U489 (
    .in(_U489_in),
    .clk(_U489_clk),
    .out(_U489_out)
);
assign _U490_in = in[1];
assign _U490_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U490 (
    .in(_U490_in),
    .clk(_U490_clk),
    .out(_U490_out)
);
assign _U491_in = in[2];
assign _U491_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U491 (
    .in(_U491_in),
    .clk(_U491_clk),
    .out(_U491_out)
);
assign _U492_in = in[3];
assign _U492_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U492 (
    .in(_U492_in),
    .clk(_U492_clk),
    .out(_U492_out)
);
assign _U493_in = in[4];
assign _U493_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U493 (
    .in(_U493_in),
    .clk(_U493_clk),
    .out(_U493_out)
);
assign out[4] = _U493_out;
assign out[3] = _U492_out;
assign out[2] = _U491_out;
assign out[1] = _U490_out;
assign out[0] = _U489_out;
endmodule

module array_delay_U481 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U482_in;
wire _U482_clk;
wire [15:0] _U482_out;
wire [15:0] _U483_in;
wire _U483_clk;
wire [15:0] _U483_out;
wire [15:0] _U484_in;
wire _U484_clk;
wire [15:0] _U484_out;
wire [15:0] _U485_in;
wire _U485_clk;
wire [15:0] _U485_out;
wire [15:0] _U486_in;
wire _U486_clk;
wire [15:0] _U486_out;
assign _U482_in = in[0];
assign _U482_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U482 (
    .in(_U482_in),
    .clk(_U482_clk),
    .out(_U482_out)
);
assign _U483_in = in[1];
assign _U483_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U483 (
    .in(_U483_in),
    .clk(_U483_clk),
    .out(_U483_out)
);
assign _U484_in = in[2];
assign _U484_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U484 (
    .in(_U484_in),
    .clk(_U484_clk),
    .out(_U484_out)
);
assign _U485_in = in[3];
assign _U485_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U485 (
    .in(_U485_in),
    .clk(_U485_clk),
    .out(_U485_out)
);
assign _U486_in = in[4];
assign _U486_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U486 (
    .in(_U486_in),
    .clk(_U486_clk),
    .out(_U486_out)
);
assign out[4] = _U486_out;
assign out[3] = _U485_out;
assign out[2] = _U484_out;
assign out[1] = _U483_out;
assign out[0] = _U482_out;
endmodule

module array_delay_U474 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U475_in;
wire _U475_clk;
wire [15:0] _U475_out;
wire [15:0] _U476_in;
wire _U476_clk;
wire [15:0] _U476_out;
wire [15:0] _U477_in;
wire _U477_clk;
wire [15:0] _U477_out;
wire [15:0] _U478_in;
wire _U478_clk;
wire [15:0] _U478_out;
wire [15:0] _U479_in;
wire _U479_clk;
wire [15:0] _U479_out;
assign _U475_in = in[0];
assign _U475_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U475 (
    .in(_U475_in),
    .clk(_U475_clk),
    .out(_U475_out)
);
assign _U476_in = in[1];
assign _U476_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U476 (
    .in(_U476_in),
    .clk(_U476_clk),
    .out(_U476_out)
);
assign _U477_in = in[2];
assign _U477_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U477 (
    .in(_U477_in),
    .clk(_U477_clk),
    .out(_U477_out)
);
assign _U478_in = in[3];
assign _U478_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U478 (
    .in(_U478_in),
    .clk(_U478_clk),
    .out(_U478_out)
);
assign _U479_in = in[4];
assign _U479_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U479 (
    .in(_U479_in),
    .clk(_U479_clk),
    .out(_U479_out)
);
assign out[4] = _U479_out;
assign out[3] = _U478_out;
assign out[2] = _U477_out;
assign out[1] = _U476_out;
assign out[0] = _U475_out;
endmodule

module array_delay_U448 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U449_in;
wire _U449_clk;
wire [15:0] _U449_out;
wire [15:0] _U450_in;
wire _U450_clk;
wire [15:0] _U450_out;
wire [15:0] _U451_in;
wire _U451_clk;
wire [15:0] _U451_out;
wire [15:0] _U452_in;
wire _U452_clk;
wire [15:0] _U452_out;
wire [15:0] _U453_in;
wire _U453_clk;
wire [15:0] _U453_out;
assign _U449_in = in[0];
assign _U449_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U449 (
    .in(_U449_in),
    .clk(_U449_clk),
    .out(_U449_out)
);
assign _U450_in = in[1];
assign _U450_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U450 (
    .in(_U450_in),
    .clk(_U450_clk),
    .out(_U450_out)
);
assign _U451_in = in[2];
assign _U451_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U451 (
    .in(_U451_in),
    .clk(_U451_clk),
    .out(_U451_out)
);
assign _U452_in = in[3];
assign _U452_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U452 (
    .in(_U452_in),
    .clk(_U452_clk),
    .out(_U452_out)
);
assign _U453_in = in[4];
assign _U453_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U453 (
    .in(_U453_in),
    .clk(_U453_clk),
    .out(_U453_out)
);
assign out[4] = _U453_out;
assign out[3] = _U452_out;
assign out[2] = _U451_out;
assign out[1] = _U450_out;
assign out[0] = _U449_out;
endmodule

module array_delay_U441 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U442_in;
wire _U442_clk;
wire [15:0] _U442_out;
wire [15:0] _U443_in;
wire _U443_clk;
wire [15:0] _U443_out;
wire [15:0] _U444_in;
wire _U444_clk;
wire [15:0] _U444_out;
wire [15:0] _U445_in;
wire _U445_clk;
wire [15:0] _U445_out;
wire [15:0] _U446_in;
wire _U446_clk;
wire [15:0] _U446_out;
assign _U442_in = in[0];
assign _U442_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U442 (
    .in(_U442_in),
    .clk(_U442_clk),
    .out(_U442_out)
);
assign _U443_in = in[1];
assign _U443_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U443 (
    .in(_U443_in),
    .clk(_U443_clk),
    .out(_U443_out)
);
assign _U444_in = in[2];
assign _U444_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U444 (
    .in(_U444_in),
    .clk(_U444_clk),
    .out(_U444_out)
);
assign _U445_in = in[3];
assign _U445_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U445 (
    .in(_U445_in),
    .clk(_U445_clk),
    .out(_U445_out)
);
assign _U446_in = in[4];
assign _U446_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U446 (
    .in(_U446_in),
    .clk(_U446_clk),
    .out(_U446_out)
);
assign out[4] = _U446_out;
assign out[3] = _U445_out;
assign out[2] = _U444_out;
assign out[1] = _U443_out;
assign out[0] = _U442_out;
endmodule

module array_delay_U2280 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2281_in;
wire _U2281_clk;
wire [15:0] _U2281_out;
wire [15:0] _U2282_in;
wire _U2282_clk;
wire [15:0] _U2282_out;
wire [15:0] _U2283_in;
wire _U2283_clk;
wire [15:0] _U2283_out;
assign _U2281_in = in[0];
assign _U2281_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2281 (
    .in(_U2281_in),
    .clk(_U2281_clk),
    .out(_U2281_out)
);
assign _U2282_in = in[1];
assign _U2282_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2282 (
    .in(_U2282_in),
    .clk(_U2282_clk),
    .out(_U2282_out)
);
assign _U2283_in = in[2];
assign _U2283_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2283 (
    .in(_U2283_in),
    .clk(_U2283_clk),
    .out(_U2283_out)
);
assign out[2] = _U2283_out;
assign out[1] = _U2282_out;
assign out[0] = _U2281_out;
endmodule

module array_delay_U2275 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2276_in;
wire _U2276_clk;
wire [15:0] _U2276_out;
wire [15:0] _U2277_in;
wire _U2277_clk;
wire [15:0] _U2277_out;
wire [15:0] _U2278_in;
wire _U2278_clk;
wire [15:0] _U2278_out;
assign _U2276_in = in[0];
assign _U2276_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2276 (
    .in(_U2276_in),
    .clk(_U2276_clk),
    .out(_U2276_out)
);
assign _U2277_in = in[1];
assign _U2277_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2277 (
    .in(_U2277_in),
    .clk(_U2277_clk),
    .out(_U2277_out)
);
assign _U2278_in = in[2];
assign _U2278_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2278 (
    .in(_U2278_in),
    .clk(_U2278_clk),
    .out(_U2278_out)
);
assign out[2] = _U2278_out;
assign out[1] = _U2277_out;
assign out[0] = _U2276_out;
endmodule

module array_delay_U2266 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2267_in;
wire _U2267_clk;
wire [15:0] _U2267_out;
wire [15:0] _U2268_in;
wire _U2268_clk;
wire [15:0] _U2268_out;
wire [15:0] _U2269_in;
wire _U2269_clk;
wire [15:0] _U2269_out;
assign _U2267_in = in[0];
assign _U2267_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2267 (
    .in(_U2267_in),
    .clk(_U2267_clk),
    .out(_U2267_out)
);
assign _U2268_in = in[1];
assign _U2268_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2268 (
    .in(_U2268_in),
    .clk(_U2268_clk),
    .out(_U2268_out)
);
assign _U2269_in = in[2];
assign _U2269_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2269 (
    .in(_U2269_in),
    .clk(_U2269_clk),
    .out(_U2269_out)
);
assign out[2] = _U2269_out;
assign out[1] = _U2268_out;
assign out[0] = _U2267_out;
endmodule

module array_delay_U2261 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2262_in;
wire _U2262_clk;
wire [15:0] _U2262_out;
wire [15:0] _U2263_in;
wire _U2263_clk;
wire [15:0] _U2263_out;
wire [15:0] _U2264_in;
wire _U2264_clk;
wire [15:0] _U2264_out;
assign _U2262_in = in[0];
assign _U2262_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2262 (
    .in(_U2262_in),
    .clk(_U2262_clk),
    .out(_U2262_out)
);
assign _U2263_in = in[1];
assign _U2263_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2263 (
    .in(_U2263_in),
    .clk(_U2263_clk),
    .out(_U2263_out)
);
assign _U2264_in = in[2];
assign _U2264_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2264 (
    .in(_U2264_in),
    .clk(_U2264_clk),
    .out(_U2264_out)
);
assign out[2] = _U2264_out;
assign out[1] = _U2263_out;
assign out[0] = _U2262_out;
endmodule

module array_delay_U2233 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2234_in;
wire _U2234_clk;
wire [15:0] _U2234_out;
wire [15:0] _U2235_in;
wire _U2235_clk;
wire [15:0] _U2235_out;
wire [15:0] _U2236_in;
wire _U2236_clk;
wire [15:0] _U2236_out;
assign _U2234_in = in[0];
assign _U2234_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2234 (
    .in(_U2234_in),
    .clk(_U2234_clk),
    .out(_U2234_out)
);
assign _U2235_in = in[1];
assign _U2235_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2235 (
    .in(_U2235_in),
    .clk(_U2235_clk),
    .out(_U2235_out)
);
assign _U2236_in = in[2];
assign _U2236_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2236 (
    .in(_U2236_in),
    .clk(_U2236_clk),
    .out(_U2236_out)
);
assign out[2] = _U2236_out;
assign out[1] = _U2235_out;
assign out[0] = _U2234_out;
endmodule

module array_delay_U2228 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2229_in;
wire _U2229_clk;
wire [15:0] _U2229_out;
wire [15:0] _U2230_in;
wire _U2230_clk;
wire [15:0] _U2230_out;
wire [15:0] _U2231_in;
wire _U2231_clk;
wire [15:0] _U2231_out;
assign _U2229_in = in[0];
assign _U2229_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2229 (
    .in(_U2229_in),
    .clk(_U2229_clk),
    .out(_U2229_out)
);
assign _U2230_in = in[1];
assign _U2230_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2230 (
    .in(_U2230_in),
    .clk(_U2230_clk),
    .out(_U2230_out)
);
assign _U2231_in = in[2];
assign _U2231_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2231 (
    .in(_U2231_in),
    .clk(_U2231_clk),
    .out(_U2231_out)
);
assign out[2] = _U2231_out;
assign out[1] = _U2230_out;
assign out[0] = _U2229_out;
endmodule

module array_delay_U2219 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2220_in;
wire _U2220_clk;
wire [15:0] _U2220_out;
wire [15:0] _U2221_in;
wire _U2221_clk;
wire [15:0] _U2221_out;
wire [15:0] _U2222_in;
wire _U2222_clk;
wire [15:0] _U2222_out;
assign _U2220_in = in[0];
assign _U2220_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2220 (
    .in(_U2220_in),
    .clk(_U2220_clk),
    .out(_U2220_out)
);
assign _U2221_in = in[1];
assign _U2221_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2221 (
    .in(_U2221_in),
    .clk(_U2221_clk),
    .out(_U2221_out)
);
assign _U2222_in = in[2];
assign _U2222_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2222 (
    .in(_U2222_in),
    .clk(_U2222_clk),
    .out(_U2222_out)
);
assign out[2] = _U2222_out;
assign out[1] = _U2221_out;
assign out[0] = _U2220_out;
endmodule

module array_delay_U2214 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2215_in;
wire _U2215_clk;
wire [15:0] _U2215_out;
wire [15:0] _U2216_in;
wire _U2216_clk;
wire [15:0] _U2216_out;
wire [15:0] _U2217_in;
wire _U2217_clk;
wire [15:0] _U2217_out;
assign _U2215_in = in[0];
assign _U2215_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2215 (
    .in(_U2215_in),
    .clk(_U2215_clk),
    .out(_U2215_out)
);
assign _U2216_in = in[1];
assign _U2216_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2216 (
    .in(_U2216_in),
    .clk(_U2216_clk),
    .out(_U2216_out)
);
assign _U2217_in = in[2];
assign _U2217_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2217 (
    .in(_U2217_in),
    .clk(_U2217_clk),
    .out(_U2217_out)
);
assign out[2] = _U2217_out;
assign out[1] = _U2216_out;
assign out[0] = _U2215_out;
endmodule

module array_delay_U2186 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2187_in;
wire _U2187_clk;
wire [15:0] _U2187_out;
wire [15:0] _U2188_in;
wire _U2188_clk;
wire [15:0] _U2188_out;
wire [15:0] _U2189_in;
wire _U2189_clk;
wire [15:0] _U2189_out;
assign _U2187_in = in[0];
assign _U2187_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2187 (
    .in(_U2187_in),
    .clk(_U2187_clk),
    .out(_U2187_out)
);
assign _U2188_in = in[1];
assign _U2188_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2188 (
    .in(_U2188_in),
    .clk(_U2188_clk),
    .out(_U2188_out)
);
assign _U2189_in = in[2];
assign _U2189_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2189 (
    .in(_U2189_in),
    .clk(_U2189_clk),
    .out(_U2189_out)
);
assign out[2] = _U2189_out;
assign out[1] = _U2188_out;
assign out[0] = _U2187_out;
endmodule

module array_delay_U2181 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2182_in;
wire _U2182_clk;
wire [15:0] _U2182_out;
wire [15:0] _U2183_in;
wire _U2183_clk;
wire [15:0] _U2183_out;
wire [15:0] _U2184_in;
wire _U2184_clk;
wire [15:0] _U2184_out;
assign _U2182_in = in[0];
assign _U2182_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2182 (
    .in(_U2182_in),
    .clk(_U2182_clk),
    .out(_U2182_out)
);
assign _U2183_in = in[1];
assign _U2183_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2183 (
    .in(_U2183_in),
    .clk(_U2183_clk),
    .out(_U2183_out)
);
assign _U2184_in = in[2];
assign _U2184_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2184 (
    .in(_U2184_in),
    .clk(_U2184_clk),
    .out(_U2184_out)
);
assign out[2] = _U2184_out;
assign out[1] = _U2183_out;
assign out[0] = _U2182_out;
endmodule

module array_delay_U2172 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2173_in;
wire _U2173_clk;
wire [15:0] _U2173_out;
wire [15:0] _U2174_in;
wire _U2174_clk;
wire [15:0] _U2174_out;
wire [15:0] _U2175_in;
wire _U2175_clk;
wire [15:0] _U2175_out;
assign _U2173_in = in[0];
assign _U2173_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2173 (
    .in(_U2173_in),
    .clk(_U2173_clk),
    .out(_U2173_out)
);
assign _U2174_in = in[1];
assign _U2174_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2174 (
    .in(_U2174_in),
    .clk(_U2174_clk),
    .out(_U2174_out)
);
assign _U2175_in = in[2];
assign _U2175_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2175 (
    .in(_U2175_in),
    .clk(_U2175_clk),
    .out(_U2175_out)
);
assign out[2] = _U2175_out;
assign out[1] = _U2174_out;
assign out[0] = _U2173_out;
endmodule

module array_delay_U2167 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2168_in;
wire _U2168_clk;
wire [15:0] _U2168_out;
wire [15:0] _U2169_in;
wire _U2169_clk;
wire [15:0] _U2169_out;
wire [15:0] _U2170_in;
wire _U2170_clk;
wire [15:0] _U2170_out;
assign _U2168_in = in[0];
assign _U2168_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2168 (
    .in(_U2168_in),
    .clk(_U2168_clk),
    .out(_U2168_out)
);
assign _U2169_in = in[1];
assign _U2169_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2169 (
    .in(_U2169_in),
    .clk(_U2169_clk),
    .out(_U2169_out)
);
assign _U2170_in = in[2];
assign _U2170_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2170 (
    .in(_U2170_in),
    .clk(_U2170_clk),
    .out(_U2170_out)
);
assign out[2] = _U2170_out;
assign out[1] = _U2169_out;
assign out[0] = _U2168_out;
endmodule

module array_delay_U2139 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2140_in;
wire _U2140_clk;
wire [15:0] _U2140_out;
wire [15:0] _U2141_in;
wire _U2141_clk;
wire [15:0] _U2141_out;
wire [15:0] _U2142_in;
wire _U2142_clk;
wire [15:0] _U2142_out;
assign _U2140_in = in[0];
assign _U2140_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2140 (
    .in(_U2140_in),
    .clk(_U2140_clk),
    .out(_U2140_out)
);
assign _U2141_in = in[1];
assign _U2141_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2141 (
    .in(_U2141_in),
    .clk(_U2141_clk),
    .out(_U2141_out)
);
assign _U2142_in = in[2];
assign _U2142_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2142 (
    .in(_U2142_in),
    .clk(_U2142_clk),
    .out(_U2142_out)
);
assign out[2] = _U2142_out;
assign out[1] = _U2141_out;
assign out[0] = _U2140_out;
endmodule

module array_delay_U2134 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2135_in;
wire _U2135_clk;
wire [15:0] _U2135_out;
wire [15:0] _U2136_in;
wire _U2136_clk;
wire [15:0] _U2136_out;
wire [15:0] _U2137_in;
wire _U2137_clk;
wire [15:0] _U2137_out;
assign _U2135_in = in[0];
assign _U2135_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2135 (
    .in(_U2135_in),
    .clk(_U2135_clk),
    .out(_U2135_out)
);
assign _U2136_in = in[1];
assign _U2136_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2136 (
    .in(_U2136_in),
    .clk(_U2136_clk),
    .out(_U2136_out)
);
assign _U2137_in = in[2];
assign _U2137_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2137 (
    .in(_U2137_in),
    .clk(_U2137_clk),
    .out(_U2137_out)
);
assign out[2] = _U2137_out;
assign out[1] = _U2136_out;
assign out[0] = _U2135_out;
endmodule

module array_delay_U2125 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2126_in;
wire _U2126_clk;
wire [15:0] _U2126_out;
wire [15:0] _U2127_in;
wire _U2127_clk;
wire [15:0] _U2127_out;
wire [15:0] _U2128_in;
wire _U2128_clk;
wire [15:0] _U2128_out;
assign _U2126_in = in[0];
assign _U2126_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2126 (
    .in(_U2126_in),
    .clk(_U2126_clk),
    .out(_U2126_out)
);
assign _U2127_in = in[1];
assign _U2127_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2127 (
    .in(_U2127_in),
    .clk(_U2127_clk),
    .out(_U2127_out)
);
assign _U2128_in = in[2];
assign _U2128_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2128 (
    .in(_U2128_in),
    .clk(_U2128_clk),
    .out(_U2128_out)
);
assign out[2] = _U2128_out;
assign out[1] = _U2127_out;
assign out[0] = _U2126_out;
endmodule

module array_delay_U2120 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2121_in;
wire _U2121_clk;
wire [15:0] _U2121_out;
wire [15:0] _U2122_in;
wire _U2122_clk;
wire [15:0] _U2122_out;
wire [15:0] _U2123_in;
wire _U2123_clk;
wire [15:0] _U2123_out;
assign _U2121_in = in[0];
assign _U2121_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2121 (
    .in(_U2121_in),
    .clk(_U2121_clk),
    .out(_U2121_out)
);
assign _U2122_in = in[1];
assign _U2122_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2122 (
    .in(_U2122_in),
    .clk(_U2122_clk),
    .out(_U2122_out)
);
assign _U2123_in = in[2];
assign _U2123_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2123 (
    .in(_U2123_in),
    .clk(_U2123_clk),
    .out(_U2123_out)
);
assign out[2] = _U2123_out;
assign out[1] = _U2122_out;
assign out[0] = _U2121_out;
endmodule

module array_delay_U2092 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2093_in;
wire _U2093_clk;
wire [15:0] _U2093_out;
wire [15:0] _U2094_in;
wire _U2094_clk;
wire [15:0] _U2094_out;
wire [15:0] _U2095_in;
wire _U2095_clk;
wire [15:0] _U2095_out;
assign _U2093_in = in[0];
assign _U2093_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2093 (
    .in(_U2093_in),
    .clk(_U2093_clk),
    .out(_U2093_out)
);
assign _U2094_in = in[1];
assign _U2094_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2094 (
    .in(_U2094_in),
    .clk(_U2094_clk),
    .out(_U2094_out)
);
assign _U2095_in = in[2];
assign _U2095_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2095 (
    .in(_U2095_in),
    .clk(_U2095_clk),
    .out(_U2095_out)
);
assign out[2] = _U2095_out;
assign out[1] = _U2094_out;
assign out[0] = _U2093_out;
endmodule

module array_delay_U2087 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2088_in;
wire _U2088_clk;
wire [15:0] _U2088_out;
wire [15:0] _U2089_in;
wire _U2089_clk;
wire [15:0] _U2089_out;
wire [15:0] _U2090_in;
wire _U2090_clk;
wire [15:0] _U2090_out;
assign _U2088_in = in[0];
assign _U2088_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2088 (
    .in(_U2088_in),
    .clk(_U2088_clk),
    .out(_U2088_out)
);
assign _U2089_in = in[1];
assign _U2089_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2089 (
    .in(_U2089_in),
    .clk(_U2089_clk),
    .out(_U2089_out)
);
assign _U2090_in = in[2];
assign _U2090_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2090 (
    .in(_U2090_in),
    .clk(_U2090_clk),
    .out(_U2090_out)
);
assign out[2] = _U2090_out;
assign out[1] = _U2089_out;
assign out[0] = _U2088_out;
endmodule

module array_delay_U2078 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2079_in;
wire _U2079_clk;
wire [15:0] _U2079_out;
wire [15:0] _U2080_in;
wire _U2080_clk;
wire [15:0] _U2080_out;
wire [15:0] _U2081_in;
wire _U2081_clk;
wire [15:0] _U2081_out;
assign _U2079_in = in[0];
assign _U2079_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2079 (
    .in(_U2079_in),
    .clk(_U2079_clk),
    .out(_U2079_out)
);
assign _U2080_in = in[1];
assign _U2080_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2080 (
    .in(_U2080_in),
    .clk(_U2080_clk),
    .out(_U2080_out)
);
assign _U2081_in = in[2];
assign _U2081_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2081 (
    .in(_U2081_in),
    .clk(_U2081_clk),
    .out(_U2081_out)
);
assign out[2] = _U2081_out;
assign out[1] = _U2080_out;
assign out[0] = _U2079_out;
endmodule

module array_delay_U2073 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2074_in;
wire _U2074_clk;
wire [15:0] _U2074_out;
wire [15:0] _U2075_in;
wire _U2075_clk;
wire [15:0] _U2075_out;
wire [15:0] _U2076_in;
wire _U2076_clk;
wire [15:0] _U2076_out;
assign _U2074_in = in[0];
assign _U2074_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2074 (
    .in(_U2074_in),
    .clk(_U2074_clk),
    .out(_U2074_out)
);
assign _U2075_in = in[1];
assign _U2075_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2075 (
    .in(_U2075_in),
    .clk(_U2075_clk),
    .out(_U2075_out)
);
assign _U2076_in = in[2];
assign _U2076_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2076 (
    .in(_U2076_in),
    .clk(_U2076_clk),
    .out(_U2076_out)
);
assign out[2] = _U2076_out;
assign out[1] = _U2075_out;
assign out[0] = _U2074_out;
endmodule

module array_delay_U2045 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2046_in;
wire _U2046_clk;
wire [15:0] _U2046_out;
wire [15:0] _U2047_in;
wire _U2047_clk;
wire [15:0] _U2047_out;
wire [15:0] _U2048_in;
wire _U2048_clk;
wire [15:0] _U2048_out;
assign _U2046_in = in[0];
assign _U2046_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2046 (
    .in(_U2046_in),
    .clk(_U2046_clk),
    .out(_U2046_out)
);
assign _U2047_in = in[1];
assign _U2047_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2047 (
    .in(_U2047_in),
    .clk(_U2047_clk),
    .out(_U2047_out)
);
assign _U2048_in = in[2];
assign _U2048_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2048 (
    .in(_U2048_in),
    .clk(_U2048_clk),
    .out(_U2048_out)
);
assign out[2] = _U2048_out;
assign out[1] = _U2047_out;
assign out[0] = _U2046_out;
endmodule

module array_delay_U2040 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2041_in;
wire _U2041_clk;
wire [15:0] _U2041_out;
wire [15:0] _U2042_in;
wire _U2042_clk;
wire [15:0] _U2042_out;
wire [15:0] _U2043_in;
wire _U2043_clk;
wire [15:0] _U2043_out;
assign _U2041_in = in[0];
assign _U2041_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2041 (
    .in(_U2041_in),
    .clk(_U2041_clk),
    .out(_U2041_out)
);
assign _U2042_in = in[1];
assign _U2042_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2042 (
    .in(_U2042_in),
    .clk(_U2042_clk),
    .out(_U2042_out)
);
assign _U2043_in = in[2];
assign _U2043_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2043 (
    .in(_U2043_in),
    .clk(_U2043_clk),
    .out(_U2043_out)
);
assign out[2] = _U2043_out;
assign out[1] = _U2042_out;
assign out[0] = _U2041_out;
endmodule

module array_delay_U2031 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2032_in;
wire _U2032_clk;
wire [15:0] _U2032_out;
wire [15:0] _U2033_in;
wire _U2033_clk;
wire [15:0] _U2033_out;
wire [15:0] _U2034_in;
wire _U2034_clk;
wire [15:0] _U2034_out;
assign _U2032_in = in[0];
assign _U2032_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2032 (
    .in(_U2032_in),
    .clk(_U2032_clk),
    .out(_U2032_out)
);
assign _U2033_in = in[1];
assign _U2033_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2033 (
    .in(_U2033_in),
    .clk(_U2033_clk),
    .out(_U2033_out)
);
assign _U2034_in = in[2];
assign _U2034_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2034 (
    .in(_U2034_in),
    .clk(_U2034_clk),
    .out(_U2034_out)
);
assign out[2] = _U2034_out;
assign out[1] = _U2033_out;
assign out[0] = _U2032_out;
endmodule

module array_delay_U2026 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U2027_in;
wire _U2027_clk;
wire [15:0] _U2027_out;
wire [15:0] _U2028_in;
wire _U2028_clk;
wire [15:0] _U2028_out;
wire [15:0] _U2029_in;
wire _U2029_clk;
wire [15:0] _U2029_out;
assign _U2027_in = in[0];
assign _U2027_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2027 (
    .in(_U2027_in),
    .clk(_U2027_clk),
    .out(_U2027_out)
);
assign _U2028_in = in[1];
assign _U2028_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2028 (
    .in(_U2028_in),
    .clk(_U2028_clk),
    .out(_U2028_out)
);
assign _U2029_in = in[2];
assign _U2029_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2029 (
    .in(_U2029_in),
    .clk(_U2029_clk),
    .out(_U2029_out)
);
assign out[2] = _U2029_out;
assign out[1] = _U2028_out;
assign out[0] = _U2027_out;
endmodule

module array_delay_U1998 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1999_in;
wire _U1999_clk;
wire [15:0] _U1999_out;
wire [15:0] _U2000_in;
wire _U2000_clk;
wire [15:0] _U2000_out;
wire [15:0] _U2001_in;
wire _U2001_clk;
wire [15:0] _U2001_out;
assign _U1999_in = in[0];
assign _U1999_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1999 (
    .in(_U1999_in),
    .clk(_U1999_clk),
    .out(_U1999_out)
);
assign _U2000_in = in[1];
assign _U2000_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2000 (
    .in(_U2000_in),
    .clk(_U2000_clk),
    .out(_U2000_out)
);
assign _U2001_in = in[2];
assign _U2001_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U2001 (
    .in(_U2001_in),
    .clk(_U2001_clk),
    .out(_U2001_out)
);
assign out[2] = _U2001_out;
assign out[1] = _U2000_out;
assign out[0] = _U1999_out;
endmodule

module array_delay_U1993 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1994_in;
wire _U1994_clk;
wire [15:0] _U1994_out;
wire [15:0] _U1995_in;
wire _U1995_clk;
wire [15:0] _U1995_out;
wire [15:0] _U1996_in;
wire _U1996_clk;
wire [15:0] _U1996_out;
assign _U1994_in = in[0];
assign _U1994_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1994 (
    .in(_U1994_in),
    .clk(_U1994_clk),
    .out(_U1994_out)
);
assign _U1995_in = in[1];
assign _U1995_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1995 (
    .in(_U1995_in),
    .clk(_U1995_clk),
    .out(_U1995_out)
);
assign _U1996_in = in[2];
assign _U1996_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1996 (
    .in(_U1996_in),
    .clk(_U1996_clk),
    .out(_U1996_out)
);
assign out[2] = _U1996_out;
assign out[1] = _U1995_out;
assign out[0] = _U1994_out;
endmodule

module array_delay_U1984 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1985_in;
wire _U1985_clk;
wire [15:0] _U1985_out;
wire [15:0] _U1986_in;
wire _U1986_clk;
wire [15:0] _U1986_out;
wire [15:0] _U1987_in;
wire _U1987_clk;
wire [15:0] _U1987_out;
assign _U1985_in = in[0];
assign _U1985_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1985 (
    .in(_U1985_in),
    .clk(_U1985_clk),
    .out(_U1985_out)
);
assign _U1986_in = in[1];
assign _U1986_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1986 (
    .in(_U1986_in),
    .clk(_U1986_clk),
    .out(_U1986_out)
);
assign _U1987_in = in[2];
assign _U1987_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1987 (
    .in(_U1987_in),
    .clk(_U1987_clk),
    .out(_U1987_out)
);
assign out[2] = _U1987_out;
assign out[1] = _U1986_out;
assign out[0] = _U1985_out;
endmodule

module array_delay_U1979 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1980_in;
wire _U1980_clk;
wire [15:0] _U1980_out;
wire [15:0] _U1981_in;
wire _U1981_clk;
wire [15:0] _U1981_out;
wire [15:0] _U1982_in;
wire _U1982_clk;
wire [15:0] _U1982_out;
assign _U1980_in = in[0];
assign _U1980_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1980 (
    .in(_U1980_in),
    .clk(_U1980_clk),
    .out(_U1980_out)
);
assign _U1981_in = in[1];
assign _U1981_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1981 (
    .in(_U1981_in),
    .clk(_U1981_clk),
    .out(_U1981_out)
);
assign _U1982_in = in[2];
assign _U1982_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1982 (
    .in(_U1982_in),
    .clk(_U1982_clk),
    .out(_U1982_out)
);
assign out[2] = _U1982_out;
assign out[1] = _U1981_out;
assign out[0] = _U1980_out;
endmodule

module array_delay_U1951 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1952_in;
wire _U1952_clk;
wire [15:0] _U1952_out;
wire [15:0] _U1953_in;
wire _U1953_clk;
wire [15:0] _U1953_out;
wire [15:0] _U1954_in;
wire _U1954_clk;
wire [15:0] _U1954_out;
assign _U1952_in = in[0];
assign _U1952_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1952 (
    .in(_U1952_in),
    .clk(_U1952_clk),
    .out(_U1952_out)
);
assign _U1953_in = in[1];
assign _U1953_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1953 (
    .in(_U1953_in),
    .clk(_U1953_clk),
    .out(_U1953_out)
);
assign _U1954_in = in[2];
assign _U1954_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1954 (
    .in(_U1954_in),
    .clk(_U1954_clk),
    .out(_U1954_out)
);
assign out[2] = _U1954_out;
assign out[1] = _U1953_out;
assign out[0] = _U1952_out;
endmodule

module array_delay_U1946 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1947_in;
wire _U1947_clk;
wire [15:0] _U1947_out;
wire [15:0] _U1948_in;
wire _U1948_clk;
wire [15:0] _U1948_out;
wire [15:0] _U1949_in;
wire _U1949_clk;
wire [15:0] _U1949_out;
assign _U1947_in = in[0];
assign _U1947_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1947 (
    .in(_U1947_in),
    .clk(_U1947_clk),
    .out(_U1947_out)
);
assign _U1948_in = in[1];
assign _U1948_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1948 (
    .in(_U1948_in),
    .clk(_U1948_clk),
    .out(_U1948_out)
);
assign _U1949_in = in[2];
assign _U1949_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1949 (
    .in(_U1949_in),
    .clk(_U1949_clk),
    .out(_U1949_out)
);
assign out[2] = _U1949_out;
assign out[1] = _U1948_out;
assign out[0] = _U1947_out;
endmodule

module array_delay_U1937 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1938_in;
wire _U1938_clk;
wire [15:0] _U1938_out;
wire [15:0] _U1939_in;
wire _U1939_clk;
wire [15:0] _U1939_out;
wire [15:0] _U1940_in;
wire _U1940_clk;
wire [15:0] _U1940_out;
assign _U1938_in = in[0];
assign _U1938_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1938 (
    .in(_U1938_in),
    .clk(_U1938_clk),
    .out(_U1938_out)
);
assign _U1939_in = in[1];
assign _U1939_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1939 (
    .in(_U1939_in),
    .clk(_U1939_clk),
    .out(_U1939_out)
);
assign _U1940_in = in[2];
assign _U1940_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1940 (
    .in(_U1940_in),
    .clk(_U1940_clk),
    .out(_U1940_out)
);
assign out[2] = _U1940_out;
assign out[1] = _U1939_out;
assign out[0] = _U1938_out;
endmodule

module array_delay_U1932 (
    input clk,
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
wire [15:0] _U1933_in;
wire _U1933_clk;
wire [15:0] _U1933_out;
wire [15:0] _U1934_in;
wire _U1934_clk;
wire [15:0] _U1934_out;
wire [15:0] _U1935_in;
wire _U1935_clk;
wire [15:0] _U1935_out;
assign _U1933_in = in[0];
assign _U1933_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1933 (
    .in(_U1933_in),
    .clk(_U1933_clk),
    .out(_U1933_out)
);
assign _U1934_in = in[1];
assign _U1934_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1934 (
    .in(_U1934_in),
    .clk(_U1934_clk),
    .out(_U1934_out)
);
assign _U1935_in = in[2];
assign _U1935_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1935 (
    .in(_U1935_in),
    .clk(_U1935_clk),
    .out(_U1935_out)
);
assign out[2] = _U1935_out;
assign out[1] = _U1934_out;
assign out[0] = _U1933_out;
endmodule

module array_delay_U1902 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1903_in;
wire _U1903_clk;
wire [15:0] _U1903_out;
wire [15:0] _U1904_in;
wire _U1904_clk;
wire [15:0] _U1904_out;
wire [15:0] _U1905_in;
wire _U1905_clk;
wire [15:0] _U1905_out;
wire [15:0] _U1906_in;
wire _U1906_clk;
wire [15:0] _U1906_out;
wire [15:0] _U1907_in;
wire _U1907_clk;
wire [15:0] _U1907_out;
assign _U1903_in = in[0];
assign _U1903_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1903 (
    .in(_U1903_in),
    .clk(_U1903_clk),
    .out(_U1903_out)
);
assign _U1904_in = in[1];
assign _U1904_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1904 (
    .in(_U1904_in),
    .clk(_U1904_clk),
    .out(_U1904_out)
);
assign _U1905_in = in[2];
assign _U1905_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1905 (
    .in(_U1905_in),
    .clk(_U1905_clk),
    .out(_U1905_out)
);
assign _U1906_in = in[3];
assign _U1906_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1906 (
    .in(_U1906_in),
    .clk(_U1906_clk),
    .out(_U1906_out)
);
assign _U1907_in = in[4];
assign _U1907_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1907 (
    .in(_U1907_in),
    .clk(_U1907_clk),
    .out(_U1907_out)
);
assign out[4] = _U1907_out;
assign out[3] = _U1906_out;
assign out[2] = _U1905_out;
assign out[1] = _U1904_out;
assign out[0] = _U1903_out;
endmodule

module array_delay_U1895 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1896_in;
wire _U1896_clk;
wire [15:0] _U1896_out;
wire [15:0] _U1897_in;
wire _U1897_clk;
wire [15:0] _U1897_out;
wire [15:0] _U1898_in;
wire _U1898_clk;
wire [15:0] _U1898_out;
wire [15:0] _U1899_in;
wire _U1899_clk;
wire [15:0] _U1899_out;
wire [15:0] _U1900_in;
wire _U1900_clk;
wire [15:0] _U1900_out;
assign _U1896_in = in[0];
assign _U1896_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1896 (
    .in(_U1896_in),
    .clk(_U1896_clk),
    .out(_U1896_out)
);
assign _U1897_in = in[1];
assign _U1897_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1897 (
    .in(_U1897_in),
    .clk(_U1897_clk),
    .out(_U1897_out)
);
assign _U1898_in = in[2];
assign _U1898_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1898 (
    .in(_U1898_in),
    .clk(_U1898_clk),
    .out(_U1898_out)
);
assign _U1899_in = in[3];
assign _U1899_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1899 (
    .in(_U1899_in),
    .clk(_U1899_clk),
    .out(_U1899_out)
);
assign _U1900_in = in[4];
assign _U1900_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1900 (
    .in(_U1900_in),
    .clk(_U1900_clk),
    .out(_U1900_out)
);
assign out[4] = _U1900_out;
assign out[3] = _U1899_out;
assign out[2] = _U1898_out;
assign out[1] = _U1897_out;
assign out[0] = _U1896_out;
endmodule

module array_delay_U1888 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1889_in;
wire _U1889_clk;
wire [15:0] _U1889_out;
wire [15:0] _U1890_in;
wire _U1890_clk;
wire [15:0] _U1890_out;
wire [15:0] _U1891_in;
wire _U1891_clk;
wire [15:0] _U1891_out;
wire [15:0] _U1892_in;
wire _U1892_clk;
wire [15:0] _U1892_out;
wire [15:0] _U1893_in;
wire _U1893_clk;
wire [15:0] _U1893_out;
assign _U1889_in = in[0];
assign _U1889_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1889 (
    .in(_U1889_in),
    .clk(_U1889_clk),
    .out(_U1889_out)
);
assign _U1890_in = in[1];
assign _U1890_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1890 (
    .in(_U1890_in),
    .clk(_U1890_clk),
    .out(_U1890_out)
);
assign _U1891_in = in[2];
assign _U1891_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1891 (
    .in(_U1891_in),
    .clk(_U1891_clk),
    .out(_U1891_out)
);
assign _U1892_in = in[3];
assign _U1892_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1892 (
    .in(_U1892_in),
    .clk(_U1892_clk),
    .out(_U1892_out)
);
assign _U1893_in = in[4];
assign _U1893_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1893 (
    .in(_U1893_in),
    .clk(_U1893_clk),
    .out(_U1893_out)
);
assign out[4] = _U1893_out;
assign out[3] = _U1892_out;
assign out[2] = _U1891_out;
assign out[1] = _U1890_out;
assign out[0] = _U1889_out;
endmodule

module array_delay_U1881 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1882_in;
wire _U1882_clk;
wire [15:0] _U1882_out;
wire [15:0] _U1883_in;
wire _U1883_clk;
wire [15:0] _U1883_out;
wire [15:0] _U1884_in;
wire _U1884_clk;
wire [15:0] _U1884_out;
wire [15:0] _U1885_in;
wire _U1885_clk;
wire [15:0] _U1885_out;
wire [15:0] _U1886_in;
wire _U1886_clk;
wire [15:0] _U1886_out;
assign _U1882_in = in[0];
assign _U1882_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1882 (
    .in(_U1882_in),
    .clk(_U1882_clk),
    .out(_U1882_out)
);
assign _U1883_in = in[1];
assign _U1883_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1883 (
    .in(_U1883_in),
    .clk(_U1883_clk),
    .out(_U1883_out)
);
assign _U1884_in = in[2];
assign _U1884_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1884 (
    .in(_U1884_in),
    .clk(_U1884_clk),
    .out(_U1884_out)
);
assign _U1885_in = in[3];
assign _U1885_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1885 (
    .in(_U1885_in),
    .clk(_U1885_clk),
    .out(_U1885_out)
);
assign _U1886_in = in[4];
assign _U1886_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1886 (
    .in(_U1886_in),
    .clk(_U1886_clk),
    .out(_U1886_out)
);
assign out[4] = _U1886_out;
assign out[3] = _U1885_out;
assign out[2] = _U1884_out;
assign out[1] = _U1883_out;
assign out[0] = _U1882_out;
endmodule

module array_delay_U1874 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1875_in;
wire _U1875_clk;
wire [15:0] _U1875_out;
wire [15:0] _U1876_in;
wire _U1876_clk;
wire [15:0] _U1876_out;
wire [15:0] _U1877_in;
wire _U1877_clk;
wire [15:0] _U1877_out;
wire [15:0] _U1878_in;
wire _U1878_clk;
wire [15:0] _U1878_out;
wire [15:0] _U1879_in;
wire _U1879_clk;
wire [15:0] _U1879_out;
assign _U1875_in = in[0];
assign _U1875_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1875 (
    .in(_U1875_in),
    .clk(_U1875_clk),
    .out(_U1875_out)
);
assign _U1876_in = in[1];
assign _U1876_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1876 (
    .in(_U1876_in),
    .clk(_U1876_clk),
    .out(_U1876_out)
);
assign _U1877_in = in[2];
assign _U1877_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1877 (
    .in(_U1877_in),
    .clk(_U1877_clk),
    .out(_U1877_out)
);
assign _U1878_in = in[3];
assign _U1878_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1878 (
    .in(_U1878_in),
    .clk(_U1878_clk),
    .out(_U1878_out)
);
assign _U1879_in = in[4];
assign _U1879_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1879 (
    .in(_U1879_in),
    .clk(_U1879_clk),
    .out(_U1879_out)
);
assign out[4] = _U1879_out;
assign out[3] = _U1878_out;
assign out[2] = _U1877_out;
assign out[1] = _U1876_out;
assign out[0] = _U1875_out;
endmodule

module array_delay_U1867 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1868_in;
wire _U1868_clk;
wire [15:0] _U1868_out;
wire [15:0] _U1869_in;
wire _U1869_clk;
wire [15:0] _U1869_out;
wire [15:0] _U1870_in;
wire _U1870_clk;
wire [15:0] _U1870_out;
wire [15:0] _U1871_in;
wire _U1871_clk;
wire [15:0] _U1871_out;
wire [15:0] _U1872_in;
wire _U1872_clk;
wire [15:0] _U1872_out;
assign _U1868_in = in[0];
assign _U1868_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1868 (
    .in(_U1868_in),
    .clk(_U1868_clk),
    .out(_U1868_out)
);
assign _U1869_in = in[1];
assign _U1869_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1869 (
    .in(_U1869_in),
    .clk(_U1869_clk),
    .out(_U1869_out)
);
assign _U1870_in = in[2];
assign _U1870_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1870 (
    .in(_U1870_in),
    .clk(_U1870_clk),
    .out(_U1870_out)
);
assign _U1871_in = in[3];
assign _U1871_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1871 (
    .in(_U1871_in),
    .clk(_U1871_clk),
    .out(_U1871_out)
);
assign _U1872_in = in[4];
assign _U1872_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1872 (
    .in(_U1872_in),
    .clk(_U1872_clk),
    .out(_U1872_out)
);
assign out[4] = _U1872_out;
assign out[3] = _U1871_out;
assign out[2] = _U1870_out;
assign out[1] = _U1869_out;
assign out[0] = _U1868_out;
endmodule

module array_delay_U1860 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1861_in;
wire _U1861_clk;
wire [15:0] _U1861_out;
wire [15:0] _U1862_in;
wire _U1862_clk;
wire [15:0] _U1862_out;
wire [15:0] _U1863_in;
wire _U1863_clk;
wire [15:0] _U1863_out;
wire [15:0] _U1864_in;
wire _U1864_clk;
wire [15:0] _U1864_out;
wire [15:0] _U1865_in;
wire _U1865_clk;
wire [15:0] _U1865_out;
assign _U1861_in = in[0];
assign _U1861_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1861 (
    .in(_U1861_in),
    .clk(_U1861_clk),
    .out(_U1861_out)
);
assign _U1862_in = in[1];
assign _U1862_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1862 (
    .in(_U1862_in),
    .clk(_U1862_clk),
    .out(_U1862_out)
);
assign _U1863_in = in[2];
assign _U1863_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1863 (
    .in(_U1863_in),
    .clk(_U1863_clk),
    .out(_U1863_out)
);
assign _U1864_in = in[3];
assign _U1864_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1864 (
    .in(_U1864_in),
    .clk(_U1864_clk),
    .out(_U1864_out)
);
assign _U1865_in = in[4];
assign _U1865_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1865 (
    .in(_U1865_in),
    .clk(_U1865_clk),
    .out(_U1865_out)
);
assign out[4] = _U1865_out;
assign out[3] = _U1864_out;
assign out[2] = _U1863_out;
assign out[1] = _U1862_out;
assign out[0] = _U1861_out;
endmodule

module array_delay_U1853 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1854_in;
wire _U1854_clk;
wire [15:0] _U1854_out;
wire [15:0] _U1855_in;
wire _U1855_clk;
wire [15:0] _U1855_out;
wire [15:0] _U1856_in;
wire _U1856_clk;
wire [15:0] _U1856_out;
wire [15:0] _U1857_in;
wire _U1857_clk;
wire [15:0] _U1857_out;
wire [15:0] _U1858_in;
wire _U1858_clk;
wire [15:0] _U1858_out;
assign _U1854_in = in[0];
assign _U1854_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1854 (
    .in(_U1854_in),
    .clk(_U1854_clk),
    .out(_U1854_out)
);
assign _U1855_in = in[1];
assign _U1855_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1855 (
    .in(_U1855_in),
    .clk(_U1855_clk),
    .out(_U1855_out)
);
assign _U1856_in = in[2];
assign _U1856_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1856 (
    .in(_U1856_in),
    .clk(_U1856_clk),
    .out(_U1856_out)
);
assign _U1857_in = in[3];
assign _U1857_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1857 (
    .in(_U1857_in),
    .clk(_U1857_clk),
    .out(_U1857_out)
);
assign _U1858_in = in[4];
assign _U1858_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1858 (
    .in(_U1858_in),
    .clk(_U1858_clk),
    .out(_U1858_out)
);
assign out[4] = _U1858_out;
assign out[3] = _U1857_out;
assign out[2] = _U1856_out;
assign out[1] = _U1855_out;
assign out[0] = _U1854_out;
endmodule

module array_delay_U1846 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1847_in;
wire _U1847_clk;
wire [15:0] _U1847_out;
wire [15:0] _U1848_in;
wire _U1848_clk;
wire [15:0] _U1848_out;
wire [15:0] _U1849_in;
wire _U1849_clk;
wire [15:0] _U1849_out;
wire [15:0] _U1850_in;
wire _U1850_clk;
wire [15:0] _U1850_out;
wire [15:0] _U1851_in;
wire _U1851_clk;
wire [15:0] _U1851_out;
assign _U1847_in = in[0];
assign _U1847_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1847 (
    .in(_U1847_in),
    .clk(_U1847_clk),
    .out(_U1847_out)
);
assign _U1848_in = in[1];
assign _U1848_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1848 (
    .in(_U1848_in),
    .clk(_U1848_clk),
    .out(_U1848_out)
);
assign _U1849_in = in[2];
assign _U1849_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1849 (
    .in(_U1849_in),
    .clk(_U1849_clk),
    .out(_U1849_out)
);
assign _U1850_in = in[3];
assign _U1850_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1850 (
    .in(_U1850_in),
    .clk(_U1850_clk),
    .out(_U1850_out)
);
assign _U1851_in = in[4];
assign _U1851_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1851 (
    .in(_U1851_in),
    .clk(_U1851_clk),
    .out(_U1851_out)
);
assign out[4] = _U1851_out;
assign out[3] = _U1850_out;
assign out[2] = _U1849_out;
assign out[1] = _U1848_out;
assign out[0] = _U1847_out;
endmodule

module array_delay_U1839 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1840_in;
wire _U1840_clk;
wire [15:0] _U1840_out;
wire [15:0] _U1841_in;
wire _U1841_clk;
wire [15:0] _U1841_out;
wire [15:0] _U1842_in;
wire _U1842_clk;
wire [15:0] _U1842_out;
wire [15:0] _U1843_in;
wire _U1843_clk;
wire [15:0] _U1843_out;
wire [15:0] _U1844_in;
wire _U1844_clk;
wire [15:0] _U1844_out;
assign _U1840_in = in[0];
assign _U1840_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1840 (
    .in(_U1840_in),
    .clk(_U1840_clk),
    .out(_U1840_out)
);
assign _U1841_in = in[1];
assign _U1841_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1841 (
    .in(_U1841_in),
    .clk(_U1841_clk),
    .out(_U1841_out)
);
assign _U1842_in = in[2];
assign _U1842_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1842 (
    .in(_U1842_in),
    .clk(_U1842_clk),
    .out(_U1842_out)
);
assign _U1843_in = in[3];
assign _U1843_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1843 (
    .in(_U1843_in),
    .clk(_U1843_clk),
    .out(_U1843_out)
);
assign _U1844_in = in[4];
assign _U1844_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1844 (
    .in(_U1844_in),
    .clk(_U1844_clk),
    .out(_U1844_out)
);
assign out[4] = _U1844_out;
assign out[3] = _U1843_out;
assign out[2] = _U1842_out;
assign out[1] = _U1841_out;
assign out[0] = _U1840_out;
endmodule

module array_delay_U1832 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1833_in;
wire _U1833_clk;
wire [15:0] _U1833_out;
wire [15:0] _U1834_in;
wire _U1834_clk;
wire [15:0] _U1834_out;
wire [15:0] _U1835_in;
wire _U1835_clk;
wire [15:0] _U1835_out;
wire [15:0] _U1836_in;
wire _U1836_clk;
wire [15:0] _U1836_out;
wire [15:0] _U1837_in;
wire _U1837_clk;
wire [15:0] _U1837_out;
assign _U1833_in = in[0];
assign _U1833_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1833 (
    .in(_U1833_in),
    .clk(_U1833_clk),
    .out(_U1833_out)
);
assign _U1834_in = in[1];
assign _U1834_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1834 (
    .in(_U1834_in),
    .clk(_U1834_clk),
    .out(_U1834_out)
);
assign _U1835_in = in[2];
assign _U1835_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1835 (
    .in(_U1835_in),
    .clk(_U1835_clk),
    .out(_U1835_out)
);
assign _U1836_in = in[3];
assign _U1836_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1836 (
    .in(_U1836_in),
    .clk(_U1836_clk),
    .out(_U1836_out)
);
assign _U1837_in = in[4];
assign _U1837_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1837 (
    .in(_U1837_in),
    .clk(_U1837_clk),
    .out(_U1837_out)
);
assign out[4] = _U1837_out;
assign out[3] = _U1836_out;
assign out[2] = _U1835_out;
assign out[1] = _U1834_out;
assign out[0] = _U1833_out;
endmodule

module array_delay_U1825 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1826_in;
wire _U1826_clk;
wire [15:0] _U1826_out;
wire [15:0] _U1827_in;
wire _U1827_clk;
wire [15:0] _U1827_out;
wire [15:0] _U1828_in;
wire _U1828_clk;
wire [15:0] _U1828_out;
wire [15:0] _U1829_in;
wire _U1829_clk;
wire [15:0] _U1829_out;
wire [15:0] _U1830_in;
wire _U1830_clk;
wire [15:0] _U1830_out;
assign _U1826_in = in[0];
assign _U1826_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1826 (
    .in(_U1826_in),
    .clk(_U1826_clk),
    .out(_U1826_out)
);
assign _U1827_in = in[1];
assign _U1827_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1827 (
    .in(_U1827_in),
    .clk(_U1827_clk),
    .out(_U1827_out)
);
assign _U1828_in = in[2];
assign _U1828_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1828 (
    .in(_U1828_in),
    .clk(_U1828_clk),
    .out(_U1828_out)
);
assign _U1829_in = in[3];
assign _U1829_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1829 (
    .in(_U1829_in),
    .clk(_U1829_clk),
    .out(_U1829_out)
);
assign _U1830_in = in[4];
assign _U1830_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1830 (
    .in(_U1830_in),
    .clk(_U1830_clk),
    .out(_U1830_out)
);
assign out[4] = _U1830_out;
assign out[3] = _U1829_out;
assign out[2] = _U1828_out;
assign out[1] = _U1827_out;
assign out[0] = _U1826_out;
endmodule

module array_delay_U1818 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1819_in;
wire _U1819_clk;
wire [15:0] _U1819_out;
wire [15:0] _U1820_in;
wire _U1820_clk;
wire [15:0] _U1820_out;
wire [15:0] _U1821_in;
wire _U1821_clk;
wire [15:0] _U1821_out;
wire [15:0] _U1822_in;
wire _U1822_clk;
wire [15:0] _U1822_out;
wire [15:0] _U1823_in;
wire _U1823_clk;
wire [15:0] _U1823_out;
assign _U1819_in = in[0];
assign _U1819_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1819 (
    .in(_U1819_in),
    .clk(_U1819_clk),
    .out(_U1819_out)
);
assign _U1820_in = in[1];
assign _U1820_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1820 (
    .in(_U1820_in),
    .clk(_U1820_clk),
    .out(_U1820_out)
);
assign _U1821_in = in[2];
assign _U1821_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1821 (
    .in(_U1821_in),
    .clk(_U1821_clk),
    .out(_U1821_out)
);
assign _U1822_in = in[3];
assign _U1822_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1822 (
    .in(_U1822_in),
    .clk(_U1822_clk),
    .out(_U1822_out)
);
assign _U1823_in = in[4];
assign _U1823_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1823 (
    .in(_U1823_in),
    .clk(_U1823_clk),
    .out(_U1823_out)
);
assign out[4] = _U1823_out;
assign out[3] = _U1822_out;
assign out[2] = _U1821_out;
assign out[1] = _U1820_out;
assign out[0] = _U1819_out;
endmodule

module array_delay_U1811 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1812_in;
wire _U1812_clk;
wire [15:0] _U1812_out;
wire [15:0] _U1813_in;
wire _U1813_clk;
wire [15:0] _U1813_out;
wire [15:0] _U1814_in;
wire _U1814_clk;
wire [15:0] _U1814_out;
wire [15:0] _U1815_in;
wire _U1815_clk;
wire [15:0] _U1815_out;
wire [15:0] _U1816_in;
wire _U1816_clk;
wire [15:0] _U1816_out;
assign _U1812_in = in[0];
assign _U1812_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1812 (
    .in(_U1812_in),
    .clk(_U1812_clk),
    .out(_U1812_out)
);
assign _U1813_in = in[1];
assign _U1813_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1813 (
    .in(_U1813_in),
    .clk(_U1813_clk),
    .out(_U1813_out)
);
assign _U1814_in = in[2];
assign _U1814_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1814 (
    .in(_U1814_in),
    .clk(_U1814_clk),
    .out(_U1814_out)
);
assign _U1815_in = in[3];
assign _U1815_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1815 (
    .in(_U1815_in),
    .clk(_U1815_clk),
    .out(_U1815_out)
);
assign _U1816_in = in[4];
assign _U1816_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1816 (
    .in(_U1816_in),
    .clk(_U1816_clk),
    .out(_U1816_out)
);
assign out[4] = _U1816_out;
assign out[3] = _U1815_out;
assign out[2] = _U1814_out;
assign out[1] = _U1813_out;
assign out[0] = _U1812_out;
endmodule

module array_delay_U1804 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1805_in;
wire _U1805_clk;
wire [15:0] _U1805_out;
wire [15:0] _U1806_in;
wire _U1806_clk;
wire [15:0] _U1806_out;
wire [15:0] _U1807_in;
wire _U1807_clk;
wire [15:0] _U1807_out;
wire [15:0] _U1808_in;
wire _U1808_clk;
wire [15:0] _U1808_out;
wire [15:0] _U1809_in;
wire _U1809_clk;
wire [15:0] _U1809_out;
assign _U1805_in = in[0];
assign _U1805_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1805 (
    .in(_U1805_in),
    .clk(_U1805_clk),
    .out(_U1805_out)
);
assign _U1806_in = in[1];
assign _U1806_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1806 (
    .in(_U1806_in),
    .clk(_U1806_clk),
    .out(_U1806_out)
);
assign _U1807_in = in[2];
assign _U1807_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1807 (
    .in(_U1807_in),
    .clk(_U1807_clk),
    .out(_U1807_out)
);
assign _U1808_in = in[3];
assign _U1808_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1808 (
    .in(_U1808_in),
    .clk(_U1808_clk),
    .out(_U1808_out)
);
assign _U1809_in = in[4];
assign _U1809_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1809 (
    .in(_U1809_in),
    .clk(_U1809_clk),
    .out(_U1809_out)
);
assign out[4] = _U1809_out;
assign out[3] = _U1808_out;
assign out[2] = _U1807_out;
assign out[1] = _U1806_out;
assign out[0] = _U1805_out;
endmodule

module array_delay_U1797 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1798_in;
wire _U1798_clk;
wire [15:0] _U1798_out;
wire [15:0] _U1799_in;
wire _U1799_clk;
wire [15:0] _U1799_out;
wire [15:0] _U1800_in;
wire _U1800_clk;
wire [15:0] _U1800_out;
wire [15:0] _U1801_in;
wire _U1801_clk;
wire [15:0] _U1801_out;
wire [15:0] _U1802_in;
wire _U1802_clk;
wire [15:0] _U1802_out;
assign _U1798_in = in[0];
assign _U1798_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1798 (
    .in(_U1798_in),
    .clk(_U1798_clk),
    .out(_U1798_out)
);
assign _U1799_in = in[1];
assign _U1799_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1799 (
    .in(_U1799_in),
    .clk(_U1799_clk),
    .out(_U1799_out)
);
assign _U1800_in = in[2];
assign _U1800_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1800 (
    .in(_U1800_in),
    .clk(_U1800_clk),
    .out(_U1800_out)
);
assign _U1801_in = in[3];
assign _U1801_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1801 (
    .in(_U1801_in),
    .clk(_U1801_clk),
    .out(_U1801_out)
);
assign _U1802_in = in[4];
assign _U1802_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1802 (
    .in(_U1802_in),
    .clk(_U1802_clk),
    .out(_U1802_out)
);
assign out[4] = _U1802_out;
assign out[3] = _U1801_out;
assign out[2] = _U1800_out;
assign out[1] = _U1799_out;
assign out[0] = _U1798_out;
endmodule

module array_delay_U1790 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1791_in;
wire _U1791_clk;
wire [15:0] _U1791_out;
wire [15:0] _U1792_in;
wire _U1792_clk;
wire [15:0] _U1792_out;
wire [15:0] _U1793_in;
wire _U1793_clk;
wire [15:0] _U1793_out;
wire [15:0] _U1794_in;
wire _U1794_clk;
wire [15:0] _U1794_out;
wire [15:0] _U1795_in;
wire _U1795_clk;
wire [15:0] _U1795_out;
assign _U1791_in = in[0];
assign _U1791_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1791 (
    .in(_U1791_in),
    .clk(_U1791_clk),
    .out(_U1791_out)
);
assign _U1792_in = in[1];
assign _U1792_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1792 (
    .in(_U1792_in),
    .clk(_U1792_clk),
    .out(_U1792_out)
);
assign _U1793_in = in[2];
assign _U1793_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1793 (
    .in(_U1793_in),
    .clk(_U1793_clk),
    .out(_U1793_out)
);
assign _U1794_in = in[3];
assign _U1794_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1794 (
    .in(_U1794_in),
    .clk(_U1794_clk),
    .out(_U1794_out)
);
assign _U1795_in = in[4];
assign _U1795_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1795 (
    .in(_U1795_in),
    .clk(_U1795_clk),
    .out(_U1795_out)
);
assign out[4] = _U1795_out;
assign out[3] = _U1794_out;
assign out[2] = _U1793_out;
assign out[1] = _U1792_out;
assign out[0] = _U1791_out;
endmodule

module array_delay_U1764 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1765_in;
wire _U1765_clk;
wire [15:0] _U1765_out;
wire [15:0] _U1766_in;
wire _U1766_clk;
wire [15:0] _U1766_out;
wire [15:0] _U1767_in;
wire _U1767_clk;
wire [15:0] _U1767_out;
wire [15:0] _U1768_in;
wire _U1768_clk;
wire [15:0] _U1768_out;
wire [15:0] _U1769_in;
wire _U1769_clk;
wire [15:0] _U1769_out;
assign _U1765_in = in[0];
assign _U1765_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1765 (
    .in(_U1765_in),
    .clk(_U1765_clk),
    .out(_U1765_out)
);
assign _U1766_in = in[1];
assign _U1766_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1766 (
    .in(_U1766_in),
    .clk(_U1766_clk),
    .out(_U1766_out)
);
assign _U1767_in = in[2];
assign _U1767_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1767 (
    .in(_U1767_in),
    .clk(_U1767_clk),
    .out(_U1767_out)
);
assign _U1768_in = in[3];
assign _U1768_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1768 (
    .in(_U1768_in),
    .clk(_U1768_clk),
    .out(_U1768_out)
);
assign _U1769_in = in[4];
assign _U1769_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1769 (
    .in(_U1769_in),
    .clk(_U1769_clk),
    .out(_U1769_out)
);
assign out[4] = _U1769_out;
assign out[3] = _U1768_out;
assign out[2] = _U1767_out;
assign out[1] = _U1766_out;
assign out[0] = _U1765_out;
endmodule

module array_delay_U1757 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1758_in;
wire _U1758_clk;
wire [15:0] _U1758_out;
wire [15:0] _U1759_in;
wire _U1759_clk;
wire [15:0] _U1759_out;
wire [15:0] _U1760_in;
wire _U1760_clk;
wire [15:0] _U1760_out;
wire [15:0] _U1761_in;
wire _U1761_clk;
wire [15:0] _U1761_out;
wire [15:0] _U1762_in;
wire _U1762_clk;
wire [15:0] _U1762_out;
assign _U1758_in = in[0];
assign _U1758_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1758 (
    .in(_U1758_in),
    .clk(_U1758_clk),
    .out(_U1758_out)
);
assign _U1759_in = in[1];
assign _U1759_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1759 (
    .in(_U1759_in),
    .clk(_U1759_clk),
    .out(_U1759_out)
);
assign _U1760_in = in[2];
assign _U1760_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1760 (
    .in(_U1760_in),
    .clk(_U1760_clk),
    .out(_U1760_out)
);
assign _U1761_in = in[3];
assign _U1761_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1761 (
    .in(_U1761_in),
    .clk(_U1761_clk),
    .out(_U1761_out)
);
assign _U1762_in = in[4];
assign _U1762_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1762 (
    .in(_U1762_in),
    .clk(_U1762_clk),
    .out(_U1762_out)
);
assign out[4] = _U1762_out;
assign out[3] = _U1761_out;
assign out[2] = _U1760_out;
assign out[1] = _U1759_out;
assign out[0] = _U1758_out;
endmodule

module array_delay_U1714 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1715_in;
wire _U1715_clk;
wire [15:0] _U1715_out;
wire [15:0] _U1716_in;
wire _U1716_clk;
wire [15:0] _U1716_out;
wire [15:0] _U1717_in;
wire _U1717_clk;
wire [15:0] _U1717_out;
wire [15:0] _U1718_in;
wire _U1718_clk;
wire [15:0] _U1718_out;
wire [15:0] _U1719_in;
wire _U1719_clk;
wire [15:0] _U1719_out;
assign _U1715_in = in[0];
assign _U1715_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1715 (
    .in(_U1715_in),
    .clk(_U1715_clk),
    .out(_U1715_out)
);
assign _U1716_in = in[1];
assign _U1716_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1716 (
    .in(_U1716_in),
    .clk(_U1716_clk),
    .out(_U1716_out)
);
assign _U1717_in = in[2];
assign _U1717_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1717 (
    .in(_U1717_in),
    .clk(_U1717_clk),
    .out(_U1717_out)
);
assign _U1718_in = in[3];
assign _U1718_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1718 (
    .in(_U1718_in),
    .clk(_U1718_clk),
    .out(_U1718_out)
);
assign _U1719_in = in[4];
assign _U1719_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1719 (
    .in(_U1719_in),
    .clk(_U1719_clk),
    .out(_U1719_out)
);
assign out[4] = _U1719_out;
assign out[3] = _U1718_out;
assign out[2] = _U1717_out;
assign out[1] = _U1716_out;
assign out[0] = _U1715_out;
endmodule

module array_delay_U1707 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1708_in;
wire _U1708_clk;
wire [15:0] _U1708_out;
wire [15:0] _U1709_in;
wire _U1709_clk;
wire [15:0] _U1709_out;
wire [15:0] _U1710_in;
wire _U1710_clk;
wire [15:0] _U1710_out;
wire [15:0] _U1711_in;
wire _U1711_clk;
wire [15:0] _U1711_out;
wire [15:0] _U1712_in;
wire _U1712_clk;
wire [15:0] _U1712_out;
assign _U1708_in = in[0];
assign _U1708_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1708 (
    .in(_U1708_in),
    .clk(_U1708_clk),
    .out(_U1708_out)
);
assign _U1709_in = in[1];
assign _U1709_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1709 (
    .in(_U1709_in),
    .clk(_U1709_clk),
    .out(_U1709_out)
);
assign _U1710_in = in[2];
assign _U1710_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1710 (
    .in(_U1710_in),
    .clk(_U1710_clk),
    .out(_U1710_out)
);
assign _U1711_in = in[3];
assign _U1711_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1711 (
    .in(_U1711_in),
    .clk(_U1711_clk),
    .out(_U1711_out)
);
assign _U1712_in = in[4];
assign _U1712_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1712 (
    .in(_U1712_in),
    .clk(_U1712_clk),
    .out(_U1712_out)
);
assign out[4] = _U1712_out;
assign out[3] = _U1711_out;
assign out[2] = _U1710_out;
assign out[1] = _U1709_out;
assign out[0] = _U1708_out;
endmodule

module array_delay_U1700 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1701_in;
wire _U1701_clk;
wire [15:0] _U1701_out;
wire [15:0] _U1702_in;
wire _U1702_clk;
wire [15:0] _U1702_out;
wire [15:0] _U1703_in;
wire _U1703_clk;
wire [15:0] _U1703_out;
wire [15:0] _U1704_in;
wire _U1704_clk;
wire [15:0] _U1704_out;
wire [15:0] _U1705_in;
wire _U1705_clk;
wire [15:0] _U1705_out;
assign _U1701_in = in[0];
assign _U1701_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1701 (
    .in(_U1701_in),
    .clk(_U1701_clk),
    .out(_U1701_out)
);
assign _U1702_in = in[1];
assign _U1702_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1702 (
    .in(_U1702_in),
    .clk(_U1702_clk),
    .out(_U1702_out)
);
assign _U1703_in = in[2];
assign _U1703_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1703 (
    .in(_U1703_in),
    .clk(_U1703_clk),
    .out(_U1703_out)
);
assign _U1704_in = in[3];
assign _U1704_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1704 (
    .in(_U1704_in),
    .clk(_U1704_clk),
    .out(_U1704_out)
);
assign _U1705_in = in[4];
assign _U1705_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1705 (
    .in(_U1705_in),
    .clk(_U1705_clk),
    .out(_U1705_out)
);
assign out[4] = _U1705_out;
assign out[3] = _U1704_out;
assign out[2] = _U1703_out;
assign out[1] = _U1702_out;
assign out[0] = _U1701_out;
endmodule

module array_delay_U1693 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1694_in;
wire _U1694_clk;
wire [15:0] _U1694_out;
wire [15:0] _U1695_in;
wire _U1695_clk;
wire [15:0] _U1695_out;
wire [15:0] _U1696_in;
wire _U1696_clk;
wire [15:0] _U1696_out;
wire [15:0] _U1697_in;
wire _U1697_clk;
wire [15:0] _U1697_out;
wire [15:0] _U1698_in;
wire _U1698_clk;
wire [15:0] _U1698_out;
assign _U1694_in = in[0];
assign _U1694_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1694 (
    .in(_U1694_in),
    .clk(_U1694_clk),
    .out(_U1694_out)
);
assign _U1695_in = in[1];
assign _U1695_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1695 (
    .in(_U1695_in),
    .clk(_U1695_clk),
    .out(_U1695_out)
);
assign _U1696_in = in[2];
assign _U1696_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1696 (
    .in(_U1696_in),
    .clk(_U1696_clk),
    .out(_U1696_out)
);
assign _U1697_in = in[3];
assign _U1697_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1697 (
    .in(_U1697_in),
    .clk(_U1697_clk),
    .out(_U1697_out)
);
assign _U1698_in = in[4];
assign _U1698_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1698 (
    .in(_U1698_in),
    .clk(_U1698_clk),
    .out(_U1698_out)
);
assign out[4] = _U1698_out;
assign out[3] = _U1697_out;
assign out[2] = _U1696_out;
assign out[1] = _U1695_out;
assign out[0] = _U1694_out;
endmodule

module array_delay_U1686 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1687_in;
wire _U1687_clk;
wire [15:0] _U1687_out;
wire [15:0] _U1688_in;
wire _U1688_clk;
wire [15:0] _U1688_out;
wire [15:0] _U1689_in;
wire _U1689_clk;
wire [15:0] _U1689_out;
wire [15:0] _U1690_in;
wire _U1690_clk;
wire [15:0] _U1690_out;
wire [15:0] _U1691_in;
wire _U1691_clk;
wire [15:0] _U1691_out;
assign _U1687_in = in[0];
assign _U1687_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1687 (
    .in(_U1687_in),
    .clk(_U1687_clk),
    .out(_U1687_out)
);
assign _U1688_in = in[1];
assign _U1688_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1688 (
    .in(_U1688_in),
    .clk(_U1688_clk),
    .out(_U1688_out)
);
assign _U1689_in = in[2];
assign _U1689_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1689 (
    .in(_U1689_in),
    .clk(_U1689_clk),
    .out(_U1689_out)
);
assign _U1690_in = in[3];
assign _U1690_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1690 (
    .in(_U1690_in),
    .clk(_U1690_clk),
    .out(_U1690_out)
);
assign _U1691_in = in[4];
assign _U1691_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1691 (
    .in(_U1691_in),
    .clk(_U1691_clk),
    .out(_U1691_out)
);
assign out[4] = _U1691_out;
assign out[3] = _U1690_out;
assign out[2] = _U1689_out;
assign out[1] = _U1688_out;
assign out[0] = _U1687_out;
endmodule

module array_delay_U1679 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1680_in;
wire _U1680_clk;
wire [15:0] _U1680_out;
wire [15:0] _U1681_in;
wire _U1681_clk;
wire [15:0] _U1681_out;
wire [15:0] _U1682_in;
wire _U1682_clk;
wire [15:0] _U1682_out;
wire [15:0] _U1683_in;
wire _U1683_clk;
wire [15:0] _U1683_out;
wire [15:0] _U1684_in;
wire _U1684_clk;
wire [15:0] _U1684_out;
assign _U1680_in = in[0];
assign _U1680_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1680 (
    .in(_U1680_in),
    .clk(_U1680_clk),
    .out(_U1680_out)
);
assign _U1681_in = in[1];
assign _U1681_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1681 (
    .in(_U1681_in),
    .clk(_U1681_clk),
    .out(_U1681_out)
);
assign _U1682_in = in[2];
assign _U1682_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1682 (
    .in(_U1682_in),
    .clk(_U1682_clk),
    .out(_U1682_out)
);
assign _U1683_in = in[3];
assign _U1683_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1683 (
    .in(_U1683_in),
    .clk(_U1683_clk),
    .out(_U1683_out)
);
assign _U1684_in = in[4];
assign _U1684_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1684 (
    .in(_U1684_in),
    .clk(_U1684_clk),
    .out(_U1684_out)
);
assign out[4] = _U1684_out;
assign out[3] = _U1683_out;
assign out[2] = _U1682_out;
assign out[1] = _U1681_out;
assign out[0] = _U1680_out;
endmodule

module array_delay_U1672 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1673_in;
wire _U1673_clk;
wire [15:0] _U1673_out;
wire [15:0] _U1674_in;
wire _U1674_clk;
wire [15:0] _U1674_out;
wire [15:0] _U1675_in;
wire _U1675_clk;
wire [15:0] _U1675_out;
wire [15:0] _U1676_in;
wire _U1676_clk;
wire [15:0] _U1676_out;
wire [15:0] _U1677_in;
wire _U1677_clk;
wire [15:0] _U1677_out;
assign _U1673_in = in[0];
assign _U1673_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1673 (
    .in(_U1673_in),
    .clk(_U1673_clk),
    .out(_U1673_out)
);
assign _U1674_in = in[1];
assign _U1674_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1674 (
    .in(_U1674_in),
    .clk(_U1674_clk),
    .out(_U1674_out)
);
assign _U1675_in = in[2];
assign _U1675_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1675 (
    .in(_U1675_in),
    .clk(_U1675_clk),
    .out(_U1675_out)
);
assign _U1676_in = in[3];
assign _U1676_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1676 (
    .in(_U1676_in),
    .clk(_U1676_clk),
    .out(_U1676_out)
);
assign _U1677_in = in[4];
assign _U1677_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1677 (
    .in(_U1677_in),
    .clk(_U1677_clk),
    .out(_U1677_out)
);
assign out[4] = _U1677_out;
assign out[3] = _U1676_out;
assign out[2] = _U1675_out;
assign out[1] = _U1674_out;
assign out[0] = _U1673_out;
endmodule

module array_delay_U1665 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1666_in;
wire _U1666_clk;
wire [15:0] _U1666_out;
wire [15:0] _U1667_in;
wire _U1667_clk;
wire [15:0] _U1667_out;
wire [15:0] _U1668_in;
wire _U1668_clk;
wire [15:0] _U1668_out;
wire [15:0] _U1669_in;
wire _U1669_clk;
wire [15:0] _U1669_out;
wire [15:0] _U1670_in;
wire _U1670_clk;
wire [15:0] _U1670_out;
assign _U1666_in = in[0];
assign _U1666_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1666 (
    .in(_U1666_in),
    .clk(_U1666_clk),
    .out(_U1666_out)
);
assign _U1667_in = in[1];
assign _U1667_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1667 (
    .in(_U1667_in),
    .clk(_U1667_clk),
    .out(_U1667_out)
);
assign _U1668_in = in[2];
assign _U1668_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1668 (
    .in(_U1668_in),
    .clk(_U1668_clk),
    .out(_U1668_out)
);
assign _U1669_in = in[3];
assign _U1669_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1669 (
    .in(_U1669_in),
    .clk(_U1669_clk),
    .out(_U1669_out)
);
assign _U1670_in = in[4];
assign _U1670_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1670 (
    .in(_U1670_in),
    .clk(_U1670_clk),
    .out(_U1670_out)
);
assign out[4] = _U1670_out;
assign out[3] = _U1669_out;
assign out[2] = _U1668_out;
assign out[1] = _U1667_out;
assign out[0] = _U1666_out;
endmodule

module array_delay_U1658 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1659_in;
wire _U1659_clk;
wire [15:0] _U1659_out;
wire [15:0] _U1660_in;
wire _U1660_clk;
wire [15:0] _U1660_out;
wire [15:0] _U1661_in;
wire _U1661_clk;
wire [15:0] _U1661_out;
wire [15:0] _U1662_in;
wire _U1662_clk;
wire [15:0] _U1662_out;
wire [15:0] _U1663_in;
wire _U1663_clk;
wire [15:0] _U1663_out;
assign _U1659_in = in[0];
assign _U1659_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1659 (
    .in(_U1659_in),
    .clk(_U1659_clk),
    .out(_U1659_out)
);
assign _U1660_in = in[1];
assign _U1660_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1660 (
    .in(_U1660_in),
    .clk(_U1660_clk),
    .out(_U1660_out)
);
assign _U1661_in = in[2];
assign _U1661_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1661 (
    .in(_U1661_in),
    .clk(_U1661_clk),
    .out(_U1661_out)
);
assign _U1662_in = in[3];
assign _U1662_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1662 (
    .in(_U1662_in),
    .clk(_U1662_clk),
    .out(_U1662_out)
);
assign _U1663_in = in[4];
assign _U1663_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1663 (
    .in(_U1663_in),
    .clk(_U1663_clk),
    .out(_U1663_out)
);
assign out[4] = _U1663_out;
assign out[3] = _U1662_out;
assign out[2] = _U1661_out;
assign out[1] = _U1660_out;
assign out[0] = _U1659_out;
endmodule

module array_delay_U1651 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1652_in;
wire _U1652_clk;
wire [15:0] _U1652_out;
wire [15:0] _U1653_in;
wire _U1653_clk;
wire [15:0] _U1653_out;
wire [15:0] _U1654_in;
wire _U1654_clk;
wire [15:0] _U1654_out;
wire [15:0] _U1655_in;
wire _U1655_clk;
wire [15:0] _U1655_out;
wire [15:0] _U1656_in;
wire _U1656_clk;
wire [15:0] _U1656_out;
assign _U1652_in = in[0];
assign _U1652_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1652 (
    .in(_U1652_in),
    .clk(_U1652_clk),
    .out(_U1652_out)
);
assign _U1653_in = in[1];
assign _U1653_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1653 (
    .in(_U1653_in),
    .clk(_U1653_clk),
    .out(_U1653_out)
);
assign _U1654_in = in[2];
assign _U1654_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1654 (
    .in(_U1654_in),
    .clk(_U1654_clk),
    .out(_U1654_out)
);
assign _U1655_in = in[3];
assign _U1655_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1655 (
    .in(_U1655_in),
    .clk(_U1655_clk),
    .out(_U1655_out)
);
assign _U1656_in = in[4];
assign _U1656_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1656 (
    .in(_U1656_in),
    .clk(_U1656_clk),
    .out(_U1656_out)
);
assign out[4] = _U1656_out;
assign out[3] = _U1655_out;
assign out[2] = _U1654_out;
assign out[1] = _U1653_out;
assign out[0] = _U1652_out;
endmodule

module array_delay_U1644 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1645_in;
wire _U1645_clk;
wire [15:0] _U1645_out;
wire [15:0] _U1646_in;
wire _U1646_clk;
wire [15:0] _U1646_out;
wire [15:0] _U1647_in;
wire _U1647_clk;
wire [15:0] _U1647_out;
wire [15:0] _U1648_in;
wire _U1648_clk;
wire [15:0] _U1648_out;
wire [15:0] _U1649_in;
wire _U1649_clk;
wire [15:0] _U1649_out;
assign _U1645_in = in[0];
assign _U1645_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1645 (
    .in(_U1645_in),
    .clk(_U1645_clk),
    .out(_U1645_out)
);
assign _U1646_in = in[1];
assign _U1646_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1646 (
    .in(_U1646_in),
    .clk(_U1646_clk),
    .out(_U1646_out)
);
assign _U1647_in = in[2];
assign _U1647_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1647 (
    .in(_U1647_in),
    .clk(_U1647_clk),
    .out(_U1647_out)
);
assign _U1648_in = in[3];
assign _U1648_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1648 (
    .in(_U1648_in),
    .clk(_U1648_clk),
    .out(_U1648_out)
);
assign _U1649_in = in[4];
assign _U1649_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1649 (
    .in(_U1649_in),
    .clk(_U1649_clk),
    .out(_U1649_out)
);
assign out[4] = _U1649_out;
assign out[3] = _U1648_out;
assign out[2] = _U1647_out;
assign out[1] = _U1646_out;
assign out[0] = _U1645_out;
endmodule

module array_delay_U1637 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1638_in;
wire _U1638_clk;
wire [15:0] _U1638_out;
wire [15:0] _U1639_in;
wire _U1639_clk;
wire [15:0] _U1639_out;
wire [15:0] _U1640_in;
wire _U1640_clk;
wire [15:0] _U1640_out;
wire [15:0] _U1641_in;
wire _U1641_clk;
wire [15:0] _U1641_out;
wire [15:0] _U1642_in;
wire _U1642_clk;
wire [15:0] _U1642_out;
assign _U1638_in = in[0];
assign _U1638_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1638 (
    .in(_U1638_in),
    .clk(_U1638_clk),
    .out(_U1638_out)
);
assign _U1639_in = in[1];
assign _U1639_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1639 (
    .in(_U1639_in),
    .clk(_U1639_clk),
    .out(_U1639_out)
);
assign _U1640_in = in[2];
assign _U1640_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1640 (
    .in(_U1640_in),
    .clk(_U1640_clk),
    .out(_U1640_out)
);
assign _U1641_in = in[3];
assign _U1641_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1641 (
    .in(_U1641_in),
    .clk(_U1641_clk),
    .out(_U1641_out)
);
assign _U1642_in = in[4];
assign _U1642_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1642 (
    .in(_U1642_in),
    .clk(_U1642_clk),
    .out(_U1642_out)
);
assign out[4] = _U1642_out;
assign out[3] = _U1641_out;
assign out[2] = _U1640_out;
assign out[1] = _U1639_out;
assign out[0] = _U1638_out;
endmodule

module array_delay_U1630 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1631_in;
wire _U1631_clk;
wire [15:0] _U1631_out;
wire [15:0] _U1632_in;
wire _U1632_clk;
wire [15:0] _U1632_out;
wire [15:0] _U1633_in;
wire _U1633_clk;
wire [15:0] _U1633_out;
wire [15:0] _U1634_in;
wire _U1634_clk;
wire [15:0] _U1634_out;
wire [15:0] _U1635_in;
wire _U1635_clk;
wire [15:0] _U1635_out;
assign _U1631_in = in[0];
assign _U1631_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1631 (
    .in(_U1631_in),
    .clk(_U1631_clk),
    .out(_U1631_out)
);
assign _U1632_in = in[1];
assign _U1632_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1632 (
    .in(_U1632_in),
    .clk(_U1632_clk),
    .out(_U1632_out)
);
assign _U1633_in = in[2];
assign _U1633_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1633 (
    .in(_U1633_in),
    .clk(_U1633_clk),
    .out(_U1633_out)
);
assign _U1634_in = in[3];
assign _U1634_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1634 (
    .in(_U1634_in),
    .clk(_U1634_clk),
    .out(_U1634_out)
);
assign _U1635_in = in[4];
assign _U1635_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1635 (
    .in(_U1635_in),
    .clk(_U1635_clk),
    .out(_U1635_out)
);
assign out[4] = _U1635_out;
assign out[3] = _U1634_out;
assign out[2] = _U1633_out;
assign out[1] = _U1632_out;
assign out[0] = _U1631_out;
endmodule

module array_delay_U1623 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1624_in;
wire _U1624_clk;
wire [15:0] _U1624_out;
wire [15:0] _U1625_in;
wire _U1625_clk;
wire [15:0] _U1625_out;
wire [15:0] _U1626_in;
wire _U1626_clk;
wire [15:0] _U1626_out;
wire [15:0] _U1627_in;
wire _U1627_clk;
wire [15:0] _U1627_out;
wire [15:0] _U1628_in;
wire _U1628_clk;
wire [15:0] _U1628_out;
assign _U1624_in = in[0];
assign _U1624_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1624 (
    .in(_U1624_in),
    .clk(_U1624_clk),
    .out(_U1624_out)
);
assign _U1625_in = in[1];
assign _U1625_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1625 (
    .in(_U1625_in),
    .clk(_U1625_clk),
    .out(_U1625_out)
);
assign _U1626_in = in[2];
assign _U1626_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1626 (
    .in(_U1626_in),
    .clk(_U1626_clk),
    .out(_U1626_out)
);
assign _U1627_in = in[3];
assign _U1627_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1627 (
    .in(_U1627_in),
    .clk(_U1627_clk),
    .out(_U1627_out)
);
assign _U1628_in = in[4];
assign _U1628_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1628 (
    .in(_U1628_in),
    .clk(_U1628_clk),
    .out(_U1628_out)
);
assign out[4] = _U1628_out;
assign out[3] = _U1627_out;
assign out[2] = _U1626_out;
assign out[1] = _U1625_out;
assign out[0] = _U1624_out;
endmodule

module array_delay_U1616 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1617_in;
wire _U1617_clk;
wire [15:0] _U1617_out;
wire [15:0] _U1618_in;
wire _U1618_clk;
wire [15:0] _U1618_out;
wire [15:0] _U1619_in;
wire _U1619_clk;
wire [15:0] _U1619_out;
wire [15:0] _U1620_in;
wire _U1620_clk;
wire [15:0] _U1620_out;
wire [15:0] _U1621_in;
wire _U1621_clk;
wire [15:0] _U1621_out;
assign _U1617_in = in[0];
assign _U1617_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1617 (
    .in(_U1617_in),
    .clk(_U1617_clk),
    .out(_U1617_out)
);
assign _U1618_in = in[1];
assign _U1618_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1618 (
    .in(_U1618_in),
    .clk(_U1618_clk),
    .out(_U1618_out)
);
assign _U1619_in = in[2];
assign _U1619_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1619 (
    .in(_U1619_in),
    .clk(_U1619_clk),
    .out(_U1619_out)
);
assign _U1620_in = in[3];
assign _U1620_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1620 (
    .in(_U1620_in),
    .clk(_U1620_clk),
    .out(_U1620_out)
);
assign _U1621_in = in[4];
assign _U1621_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1621 (
    .in(_U1621_in),
    .clk(_U1621_clk),
    .out(_U1621_out)
);
assign out[4] = _U1621_out;
assign out[3] = _U1620_out;
assign out[2] = _U1619_out;
assign out[1] = _U1618_out;
assign out[0] = _U1617_out;
endmodule

module array_delay_U1609 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1610_in;
wire _U1610_clk;
wire [15:0] _U1610_out;
wire [15:0] _U1611_in;
wire _U1611_clk;
wire [15:0] _U1611_out;
wire [15:0] _U1612_in;
wire _U1612_clk;
wire [15:0] _U1612_out;
wire [15:0] _U1613_in;
wire _U1613_clk;
wire [15:0] _U1613_out;
wire [15:0] _U1614_in;
wire _U1614_clk;
wire [15:0] _U1614_out;
assign _U1610_in = in[0];
assign _U1610_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1610 (
    .in(_U1610_in),
    .clk(_U1610_clk),
    .out(_U1610_out)
);
assign _U1611_in = in[1];
assign _U1611_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1611 (
    .in(_U1611_in),
    .clk(_U1611_clk),
    .out(_U1611_out)
);
assign _U1612_in = in[2];
assign _U1612_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1612 (
    .in(_U1612_in),
    .clk(_U1612_clk),
    .out(_U1612_out)
);
assign _U1613_in = in[3];
assign _U1613_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1613 (
    .in(_U1613_in),
    .clk(_U1613_clk),
    .out(_U1613_out)
);
assign _U1614_in = in[4];
assign _U1614_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1614 (
    .in(_U1614_in),
    .clk(_U1614_clk),
    .out(_U1614_out)
);
assign out[4] = _U1614_out;
assign out[3] = _U1613_out;
assign out[2] = _U1612_out;
assign out[1] = _U1611_out;
assign out[0] = _U1610_out;
endmodule

module array_delay_U1602 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1603_in;
wire _U1603_clk;
wire [15:0] _U1603_out;
wire [15:0] _U1604_in;
wire _U1604_clk;
wire [15:0] _U1604_out;
wire [15:0] _U1605_in;
wire _U1605_clk;
wire [15:0] _U1605_out;
wire [15:0] _U1606_in;
wire _U1606_clk;
wire [15:0] _U1606_out;
wire [15:0] _U1607_in;
wire _U1607_clk;
wire [15:0] _U1607_out;
assign _U1603_in = in[0];
assign _U1603_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1603 (
    .in(_U1603_in),
    .clk(_U1603_clk),
    .out(_U1603_out)
);
assign _U1604_in = in[1];
assign _U1604_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1604 (
    .in(_U1604_in),
    .clk(_U1604_clk),
    .out(_U1604_out)
);
assign _U1605_in = in[2];
assign _U1605_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1605 (
    .in(_U1605_in),
    .clk(_U1605_clk),
    .out(_U1605_out)
);
assign _U1606_in = in[3];
assign _U1606_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1606 (
    .in(_U1606_in),
    .clk(_U1606_clk),
    .out(_U1606_out)
);
assign _U1607_in = in[4];
assign _U1607_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1607 (
    .in(_U1607_in),
    .clk(_U1607_clk),
    .out(_U1607_out)
);
assign out[4] = _U1607_out;
assign out[3] = _U1606_out;
assign out[2] = _U1605_out;
assign out[1] = _U1604_out;
assign out[0] = _U1603_out;
endmodule

module array_delay_U1576 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1577_in;
wire _U1577_clk;
wire [15:0] _U1577_out;
wire [15:0] _U1578_in;
wire _U1578_clk;
wire [15:0] _U1578_out;
wire [15:0] _U1579_in;
wire _U1579_clk;
wire [15:0] _U1579_out;
wire [15:0] _U1580_in;
wire _U1580_clk;
wire [15:0] _U1580_out;
wire [15:0] _U1581_in;
wire _U1581_clk;
wire [15:0] _U1581_out;
assign _U1577_in = in[0];
assign _U1577_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1577 (
    .in(_U1577_in),
    .clk(_U1577_clk),
    .out(_U1577_out)
);
assign _U1578_in = in[1];
assign _U1578_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1578 (
    .in(_U1578_in),
    .clk(_U1578_clk),
    .out(_U1578_out)
);
assign _U1579_in = in[2];
assign _U1579_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1579 (
    .in(_U1579_in),
    .clk(_U1579_clk),
    .out(_U1579_out)
);
assign _U1580_in = in[3];
assign _U1580_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1580 (
    .in(_U1580_in),
    .clk(_U1580_clk),
    .out(_U1580_out)
);
assign _U1581_in = in[4];
assign _U1581_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1581 (
    .in(_U1581_in),
    .clk(_U1581_clk),
    .out(_U1581_out)
);
assign out[4] = _U1581_out;
assign out[3] = _U1580_out;
assign out[2] = _U1579_out;
assign out[1] = _U1578_out;
assign out[0] = _U1577_out;
endmodule

module array_delay_U1569 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1570_in;
wire _U1570_clk;
wire [15:0] _U1570_out;
wire [15:0] _U1571_in;
wire _U1571_clk;
wire [15:0] _U1571_out;
wire [15:0] _U1572_in;
wire _U1572_clk;
wire [15:0] _U1572_out;
wire [15:0] _U1573_in;
wire _U1573_clk;
wire [15:0] _U1573_out;
wire [15:0] _U1574_in;
wire _U1574_clk;
wire [15:0] _U1574_out;
assign _U1570_in = in[0];
assign _U1570_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1570 (
    .in(_U1570_in),
    .clk(_U1570_clk),
    .out(_U1570_out)
);
assign _U1571_in = in[1];
assign _U1571_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1571 (
    .in(_U1571_in),
    .clk(_U1571_clk),
    .out(_U1571_out)
);
assign _U1572_in = in[2];
assign _U1572_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1572 (
    .in(_U1572_in),
    .clk(_U1572_clk),
    .out(_U1572_out)
);
assign _U1573_in = in[3];
assign _U1573_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1573 (
    .in(_U1573_in),
    .clk(_U1573_clk),
    .out(_U1573_out)
);
assign _U1574_in = in[4];
assign _U1574_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1574 (
    .in(_U1574_in),
    .clk(_U1574_clk),
    .out(_U1574_out)
);
assign out[4] = _U1574_out;
assign out[3] = _U1573_out;
assign out[2] = _U1572_out;
assign out[1] = _U1571_out;
assign out[0] = _U1570_out;
endmodule

module array_delay_U1526 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1527_in;
wire _U1527_clk;
wire [15:0] _U1527_out;
wire [15:0] _U1528_in;
wire _U1528_clk;
wire [15:0] _U1528_out;
wire [15:0] _U1529_in;
wire _U1529_clk;
wire [15:0] _U1529_out;
wire [15:0] _U1530_in;
wire _U1530_clk;
wire [15:0] _U1530_out;
wire [15:0] _U1531_in;
wire _U1531_clk;
wire [15:0] _U1531_out;
assign _U1527_in = in[0];
assign _U1527_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1527 (
    .in(_U1527_in),
    .clk(_U1527_clk),
    .out(_U1527_out)
);
assign _U1528_in = in[1];
assign _U1528_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1528 (
    .in(_U1528_in),
    .clk(_U1528_clk),
    .out(_U1528_out)
);
assign _U1529_in = in[2];
assign _U1529_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1529 (
    .in(_U1529_in),
    .clk(_U1529_clk),
    .out(_U1529_out)
);
assign _U1530_in = in[3];
assign _U1530_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1530 (
    .in(_U1530_in),
    .clk(_U1530_clk),
    .out(_U1530_out)
);
assign _U1531_in = in[4];
assign _U1531_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1531 (
    .in(_U1531_in),
    .clk(_U1531_clk),
    .out(_U1531_out)
);
assign out[4] = _U1531_out;
assign out[3] = _U1530_out;
assign out[2] = _U1529_out;
assign out[1] = _U1528_out;
assign out[0] = _U1527_out;
endmodule

module array_delay_U1519 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1520_in;
wire _U1520_clk;
wire [15:0] _U1520_out;
wire [15:0] _U1521_in;
wire _U1521_clk;
wire [15:0] _U1521_out;
wire [15:0] _U1522_in;
wire _U1522_clk;
wire [15:0] _U1522_out;
wire [15:0] _U1523_in;
wire _U1523_clk;
wire [15:0] _U1523_out;
wire [15:0] _U1524_in;
wire _U1524_clk;
wire [15:0] _U1524_out;
assign _U1520_in = in[0];
assign _U1520_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1520 (
    .in(_U1520_in),
    .clk(_U1520_clk),
    .out(_U1520_out)
);
assign _U1521_in = in[1];
assign _U1521_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1521 (
    .in(_U1521_in),
    .clk(_U1521_clk),
    .out(_U1521_out)
);
assign _U1522_in = in[2];
assign _U1522_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1522 (
    .in(_U1522_in),
    .clk(_U1522_clk),
    .out(_U1522_out)
);
assign _U1523_in = in[3];
assign _U1523_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1523 (
    .in(_U1523_in),
    .clk(_U1523_clk),
    .out(_U1523_out)
);
assign _U1524_in = in[4];
assign _U1524_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1524 (
    .in(_U1524_in),
    .clk(_U1524_clk),
    .out(_U1524_out)
);
assign out[4] = _U1524_out;
assign out[3] = _U1523_out;
assign out[2] = _U1522_out;
assign out[1] = _U1521_out;
assign out[0] = _U1520_out;
endmodule

module array_delay_U1512 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1513_in;
wire _U1513_clk;
wire [15:0] _U1513_out;
wire [15:0] _U1514_in;
wire _U1514_clk;
wire [15:0] _U1514_out;
wire [15:0] _U1515_in;
wire _U1515_clk;
wire [15:0] _U1515_out;
wire [15:0] _U1516_in;
wire _U1516_clk;
wire [15:0] _U1516_out;
wire [15:0] _U1517_in;
wire _U1517_clk;
wire [15:0] _U1517_out;
assign _U1513_in = in[0];
assign _U1513_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1513 (
    .in(_U1513_in),
    .clk(_U1513_clk),
    .out(_U1513_out)
);
assign _U1514_in = in[1];
assign _U1514_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1514 (
    .in(_U1514_in),
    .clk(_U1514_clk),
    .out(_U1514_out)
);
assign _U1515_in = in[2];
assign _U1515_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1515 (
    .in(_U1515_in),
    .clk(_U1515_clk),
    .out(_U1515_out)
);
assign _U1516_in = in[3];
assign _U1516_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1516 (
    .in(_U1516_in),
    .clk(_U1516_clk),
    .out(_U1516_out)
);
assign _U1517_in = in[4];
assign _U1517_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1517 (
    .in(_U1517_in),
    .clk(_U1517_clk),
    .out(_U1517_out)
);
assign out[4] = _U1517_out;
assign out[3] = _U1516_out;
assign out[2] = _U1515_out;
assign out[1] = _U1514_out;
assign out[0] = _U1513_out;
endmodule

module array_delay_U1505 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1506_in;
wire _U1506_clk;
wire [15:0] _U1506_out;
wire [15:0] _U1507_in;
wire _U1507_clk;
wire [15:0] _U1507_out;
wire [15:0] _U1508_in;
wire _U1508_clk;
wire [15:0] _U1508_out;
wire [15:0] _U1509_in;
wire _U1509_clk;
wire [15:0] _U1509_out;
wire [15:0] _U1510_in;
wire _U1510_clk;
wire [15:0] _U1510_out;
assign _U1506_in = in[0];
assign _U1506_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1506 (
    .in(_U1506_in),
    .clk(_U1506_clk),
    .out(_U1506_out)
);
assign _U1507_in = in[1];
assign _U1507_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1507 (
    .in(_U1507_in),
    .clk(_U1507_clk),
    .out(_U1507_out)
);
assign _U1508_in = in[2];
assign _U1508_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1508 (
    .in(_U1508_in),
    .clk(_U1508_clk),
    .out(_U1508_out)
);
assign _U1509_in = in[3];
assign _U1509_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1509 (
    .in(_U1509_in),
    .clk(_U1509_clk),
    .out(_U1509_out)
);
assign _U1510_in = in[4];
assign _U1510_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1510 (
    .in(_U1510_in),
    .clk(_U1510_clk),
    .out(_U1510_out)
);
assign out[4] = _U1510_out;
assign out[3] = _U1509_out;
assign out[2] = _U1508_out;
assign out[1] = _U1507_out;
assign out[0] = _U1506_out;
endmodule

module array_delay_U1498 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1499_in;
wire _U1499_clk;
wire [15:0] _U1499_out;
wire [15:0] _U1500_in;
wire _U1500_clk;
wire [15:0] _U1500_out;
wire [15:0] _U1501_in;
wire _U1501_clk;
wire [15:0] _U1501_out;
wire [15:0] _U1502_in;
wire _U1502_clk;
wire [15:0] _U1502_out;
wire [15:0] _U1503_in;
wire _U1503_clk;
wire [15:0] _U1503_out;
assign _U1499_in = in[0];
assign _U1499_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1499 (
    .in(_U1499_in),
    .clk(_U1499_clk),
    .out(_U1499_out)
);
assign _U1500_in = in[1];
assign _U1500_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1500 (
    .in(_U1500_in),
    .clk(_U1500_clk),
    .out(_U1500_out)
);
assign _U1501_in = in[2];
assign _U1501_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1501 (
    .in(_U1501_in),
    .clk(_U1501_clk),
    .out(_U1501_out)
);
assign _U1502_in = in[3];
assign _U1502_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1502 (
    .in(_U1502_in),
    .clk(_U1502_clk),
    .out(_U1502_out)
);
assign _U1503_in = in[4];
assign _U1503_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1503 (
    .in(_U1503_in),
    .clk(_U1503_clk),
    .out(_U1503_out)
);
assign out[4] = _U1503_out;
assign out[3] = _U1502_out;
assign out[2] = _U1501_out;
assign out[1] = _U1500_out;
assign out[0] = _U1499_out;
endmodule

module array_delay_U1491 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1492_in;
wire _U1492_clk;
wire [15:0] _U1492_out;
wire [15:0] _U1493_in;
wire _U1493_clk;
wire [15:0] _U1493_out;
wire [15:0] _U1494_in;
wire _U1494_clk;
wire [15:0] _U1494_out;
wire [15:0] _U1495_in;
wire _U1495_clk;
wire [15:0] _U1495_out;
wire [15:0] _U1496_in;
wire _U1496_clk;
wire [15:0] _U1496_out;
assign _U1492_in = in[0];
assign _U1492_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1492 (
    .in(_U1492_in),
    .clk(_U1492_clk),
    .out(_U1492_out)
);
assign _U1493_in = in[1];
assign _U1493_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1493 (
    .in(_U1493_in),
    .clk(_U1493_clk),
    .out(_U1493_out)
);
assign _U1494_in = in[2];
assign _U1494_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1494 (
    .in(_U1494_in),
    .clk(_U1494_clk),
    .out(_U1494_out)
);
assign _U1495_in = in[3];
assign _U1495_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1495 (
    .in(_U1495_in),
    .clk(_U1495_clk),
    .out(_U1495_out)
);
assign _U1496_in = in[4];
assign _U1496_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1496 (
    .in(_U1496_in),
    .clk(_U1496_clk),
    .out(_U1496_out)
);
assign out[4] = _U1496_out;
assign out[3] = _U1495_out;
assign out[2] = _U1494_out;
assign out[1] = _U1493_out;
assign out[0] = _U1492_out;
endmodule

module array_delay_U1484 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1485_in;
wire _U1485_clk;
wire [15:0] _U1485_out;
wire [15:0] _U1486_in;
wire _U1486_clk;
wire [15:0] _U1486_out;
wire [15:0] _U1487_in;
wire _U1487_clk;
wire [15:0] _U1487_out;
wire [15:0] _U1488_in;
wire _U1488_clk;
wire [15:0] _U1488_out;
wire [15:0] _U1489_in;
wire _U1489_clk;
wire [15:0] _U1489_out;
assign _U1485_in = in[0];
assign _U1485_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1485 (
    .in(_U1485_in),
    .clk(_U1485_clk),
    .out(_U1485_out)
);
assign _U1486_in = in[1];
assign _U1486_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1486 (
    .in(_U1486_in),
    .clk(_U1486_clk),
    .out(_U1486_out)
);
assign _U1487_in = in[2];
assign _U1487_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1487 (
    .in(_U1487_in),
    .clk(_U1487_clk),
    .out(_U1487_out)
);
assign _U1488_in = in[3];
assign _U1488_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1488 (
    .in(_U1488_in),
    .clk(_U1488_clk),
    .out(_U1488_out)
);
assign _U1489_in = in[4];
assign _U1489_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1489 (
    .in(_U1489_in),
    .clk(_U1489_clk),
    .out(_U1489_out)
);
assign out[4] = _U1489_out;
assign out[3] = _U1488_out;
assign out[2] = _U1487_out;
assign out[1] = _U1486_out;
assign out[0] = _U1485_out;
endmodule

module array_delay_U1477 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1478_in;
wire _U1478_clk;
wire [15:0] _U1478_out;
wire [15:0] _U1479_in;
wire _U1479_clk;
wire [15:0] _U1479_out;
wire [15:0] _U1480_in;
wire _U1480_clk;
wire [15:0] _U1480_out;
wire [15:0] _U1481_in;
wire _U1481_clk;
wire [15:0] _U1481_out;
wire [15:0] _U1482_in;
wire _U1482_clk;
wire [15:0] _U1482_out;
assign _U1478_in = in[0];
assign _U1478_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1478 (
    .in(_U1478_in),
    .clk(_U1478_clk),
    .out(_U1478_out)
);
assign _U1479_in = in[1];
assign _U1479_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1479 (
    .in(_U1479_in),
    .clk(_U1479_clk),
    .out(_U1479_out)
);
assign _U1480_in = in[2];
assign _U1480_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1480 (
    .in(_U1480_in),
    .clk(_U1480_clk),
    .out(_U1480_out)
);
assign _U1481_in = in[3];
assign _U1481_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1481 (
    .in(_U1481_in),
    .clk(_U1481_clk),
    .out(_U1481_out)
);
assign _U1482_in = in[4];
assign _U1482_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1482 (
    .in(_U1482_in),
    .clk(_U1482_clk),
    .out(_U1482_out)
);
assign out[4] = _U1482_out;
assign out[3] = _U1481_out;
assign out[2] = _U1480_out;
assign out[1] = _U1479_out;
assign out[0] = _U1478_out;
endmodule

module array_delay_U1470 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1471_in;
wire _U1471_clk;
wire [15:0] _U1471_out;
wire [15:0] _U1472_in;
wire _U1472_clk;
wire [15:0] _U1472_out;
wire [15:0] _U1473_in;
wire _U1473_clk;
wire [15:0] _U1473_out;
wire [15:0] _U1474_in;
wire _U1474_clk;
wire [15:0] _U1474_out;
wire [15:0] _U1475_in;
wire _U1475_clk;
wire [15:0] _U1475_out;
assign _U1471_in = in[0];
assign _U1471_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1471 (
    .in(_U1471_in),
    .clk(_U1471_clk),
    .out(_U1471_out)
);
assign _U1472_in = in[1];
assign _U1472_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1472 (
    .in(_U1472_in),
    .clk(_U1472_clk),
    .out(_U1472_out)
);
assign _U1473_in = in[2];
assign _U1473_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1473 (
    .in(_U1473_in),
    .clk(_U1473_clk),
    .out(_U1473_out)
);
assign _U1474_in = in[3];
assign _U1474_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1474 (
    .in(_U1474_in),
    .clk(_U1474_clk),
    .out(_U1474_out)
);
assign _U1475_in = in[4];
assign _U1475_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1475 (
    .in(_U1475_in),
    .clk(_U1475_clk),
    .out(_U1475_out)
);
assign out[4] = _U1475_out;
assign out[3] = _U1474_out;
assign out[2] = _U1473_out;
assign out[1] = _U1472_out;
assign out[0] = _U1471_out;
endmodule

module array_delay_U1463 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1464_in;
wire _U1464_clk;
wire [15:0] _U1464_out;
wire [15:0] _U1465_in;
wire _U1465_clk;
wire [15:0] _U1465_out;
wire [15:0] _U1466_in;
wire _U1466_clk;
wire [15:0] _U1466_out;
wire [15:0] _U1467_in;
wire _U1467_clk;
wire [15:0] _U1467_out;
wire [15:0] _U1468_in;
wire _U1468_clk;
wire [15:0] _U1468_out;
assign _U1464_in = in[0];
assign _U1464_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1464 (
    .in(_U1464_in),
    .clk(_U1464_clk),
    .out(_U1464_out)
);
assign _U1465_in = in[1];
assign _U1465_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1465 (
    .in(_U1465_in),
    .clk(_U1465_clk),
    .out(_U1465_out)
);
assign _U1466_in = in[2];
assign _U1466_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1466 (
    .in(_U1466_in),
    .clk(_U1466_clk),
    .out(_U1466_out)
);
assign _U1467_in = in[3];
assign _U1467_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1467 (
    .in(_U1467_in),
    .clk(_U1467_clk),
    .out(_U1467_out)
);
assign _U1468_in = in[4];
assign _U1468_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1468 (
    .in(_U1468_in),
    .clk(_U1468_clk),
    .out(_U1468_out)
);
assign out[4] = _U1468_out;
assign out[3] = _U1467_out;
assign out[2] = _U1466_out;
assign out[1] = _U1465_out;
assign out[0] = _U1464_out;
endmodule

module array_delay_U1456 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1457_in;
wire _U1457_clk;
wire [15:0] _U1457_out;
wire [15:0] _U1458_in;
wire _U1458_clk;
wire [15:0] _U1458_out;
wire [15:0] _U1459_in;
wire _U1459_clk;
wire [15:0] _U1459_out;
wire [15:0] _U1460_in;
wire _U1460_clk;
wire [15:0] _U1460_out;
wire [15:0] _U1461_in;
wire _U1461_clk;
wire [15:0] _U1461_out;
assign _U1457_in = in[0];
assign _U1457_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1457 (
    .in(_U1457_in),
    .clk(_U1457_clk),
    .out(_U1457_out)
);
assign _U1458_in = in[1];
assign _U1458_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1458 (
    .in(_U1458_in),
    .clk(_U1458_clk),
    .out(_U1458_out)
);
assign _U1459_in = in[2];
assign _U1459_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1459 (
    .in(_U1459_in),
    .clk(_U1459_clk),
    .out(_U1459_out)
);
assign _U1460_in = in[3];
assign _U1460_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1460 (
    .in(_U1460_in),
    .clk(_U1460_clk),
    .out(_U1460_out)
);
assign _U1461_in = in[4];
assign _U1461_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1461 (
    .in(_U1461_in),
    .clk(_U1461_clk),
    .out(_U1461_out)
);
assign out[4] = _U1461_out;
assign out[3] = _U1460_out;
assign out[2] = _U1459_out;
assign out[1] = _U1458_out;
assign out[0] = _U1457_out;
endmodule

module array_delay_U1449 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1450_in;
wire _U1450_clk;
wire [15:0] _U1450_out;
wire [15:0] _U1451_in;
wire _U1451_clk;
wire [15:0] _U1451_out;
wire [15:0] _U1452_in;
wire _U1452_clk;
wire [15:0] _U1452_out;
wire [15:0] _U1453_in;
wire _U1453_clk;
wire [15:0] _U1453_out;
wire [15:0] _U1454_in;
wire _U1454_clk;
wire [15:0] _U1454_out;
assign _U1450_in = in[0];
assign _U1450_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1450 (
    .in(_U1450_in),
    .clk(_U1450_clk),
    .out(_U1450_out)
);
assign _U1451_in = in[1];
assign _U1451_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1451 (
    .in(_U1451_in),
    .clk(_U1451_clk),
    .out(_U1451_out)
);
assign _U1452_in = in[2];
assign _U1452_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1452 (
    .in(_U1452_in),
    .clk(_U1452_clk),
    .out(_U1452_out)
);
assign _U1453_in = in[3];
assign _U1453_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1453 (
    .in(_U1453_in),
    .clk(_U1453_clk),
    .out(_U1453_out)
);
assign _U1454_in = in[4];
assign _U1454_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1454 (
    .in(_U1454_in),
    .clk(_U1454_clk),
    .out(_U1454_out)
);
assign out[4] = _U1454_out;
assign out[3] = _U1453_out;
assign out[2] = _U1452_out;
assign out[1] = _U1451_out;
assign out[0] = _U1450_out;
endmodule

module array_delay_U1442 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1443_in;
wire _U1443_clk;
wire [15:0] _U1443_out;
wire [15:0] _U1444_in;
wire _U1444_clk;
wire [15:0] _U1444_out;
wire [15:0] _U1445_in;
wire _U1445_clk;
wire [15:0] _U1445_out;
wire [15:0] _U1446_in;
wire _U1446_clk;
wire [15:0] _U1446_out;
wire [15:0] _U1447_in;
wire _U1447_clk;
wire [15:0] _U1447_out;
assign _U1443_in = in[0];
assign _U1443_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1443 (
    .in(_U1443_in),
    .clk(_U1443_clk),
    .out(_U1443_out)
);
assign _U1444_in = in[1];
assign _U1444_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1444 (
    .in(_U1444_in),
    .clk(_U1444_clk),
    .out(_U1444_out)
);
assign _U1445_in = in[2];
assign _U1445_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1445 (
    .in(_U1445_in),
    .clk(_U1445_clk),
    .out(_U1445_out)
);
assign _U1446_in = in[3];
assign _U1446_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1446 (
    .in(_U1446_in),
    .clk(_U1446_clk),
    .out(_U1446_out)
);
assign _U1447_in = in[4];
assign _U1447_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1447 (
    .in(_U1447_in),
    .clk(_U1447_clk),
    .out(_U1447_out)
);
assign out[4] = _U1447_out;
assign out[3] = _U1446_out;
assign out[2] = _U1445_out;
assign out[1] = _U1444_out;
assign out[0] = _U1443_out;
endmodule

module array_delay_U1435 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1436_in;
wire _U1436_clk;
wire [15:0] _U1436_out;
wire [15:0] _U1437_in;
wire _U1437_clk;
wire [15:0] _U1437_out;
wire [15:0] _U1438_in;
wire _U1438_clk;
wire [15:0] _U1438_out;
wire [15:0] _U1439_in;
wire _U1439_clk;
wire [15:0] _U1439_out;
wire [15:0] _U1440_in;
wire _U1440_clk;
wire [15:0] _U1440_out;
assign _U1436_in = in[0];
assign _U1436_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1436 (
    .in(_U1436_in),
    .clk(_U1436_clk),
    .out(_U1436_out)
);
assign _U1437_in = in[1];
assign _U1437_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1437 (
    .in(_U1437_in),
    .clk(_U1437_clk),
    .out(_U1437_out)
);
assign _U1438_in = in[2];
assign _U1438_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1438 (
    .in(_U1438_in),
    .clk(_U1438_clk),
    .out(_U1438_out)
);
assign _U1439_in = in[3];
assign _U1439_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1439 (
    .in(_U1439_in),
    .clk(_U1439_clk),
    .out(_U1439_out)
);
assign _U1440_in = in[4];
assign _U1440_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1440 (
    .in(_U1440_in),
    .clk(_U1440_clk),
    .out(_U1440_out)
);
assign out[4] = _U1440_out;
assign out[3] = _U1439_out;
assign out[2] = _U1438_out;
assign out[1] = _U1437_out;
assign out[0] = _U1436_out;
endmodule

module array_delay_U1428 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1429_in;
wire _U1429_clk;
wire [15:0] _U1429_out;
wire [15:0] _U1430_in;
wire _U1430_clk;
wire [15:0] _U1430_out;
wire [15:0] _U1431_in;
wire _U1431_clk;
wire [15:0] _U1431_out;
wire [15:0] _U1432_in;
wire _U1432_clk;
wire [15:0] _U1432_out;
wire [15:0] _U1433_in;
wire _U1433_clk;
wire [15:0] _U1433_out;
assign _U1429_in = in[0];
assign _U1429_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1429 (
    .in(_U1429_in),
    .clk(_U1429_clk),
    .out(_U1429_out)
);
assign _U1430_in = in[1];
assign _U1430_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1430 (
    .in(_U1430_in),
    .clk(_U1430_clk),
    .out(_U1430_out)
);
assign _U1431_in = in[2];
assign _U1431_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1431 (
    .in(_U1431_in),
    .clk(_U1431_clk),
    .out(_U1431_out)
);
assign _U1432_in = in[3];
assign _U1432_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1432 (
    .in(_U1432_in),
    .clk(_U1432_clk),
    .out(_U1432_out)
);
assign _U1433_in = in[4];
assign _U1433_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1433 (
    .in(_U1433_in),
    .clk(_U1433_clk),
    .out(_U1433_out)
);
assign out[4] = _U1433_out;
assign out[3] = _U1432_out;
assign out[2] = _U1431_out;
assign out[1] = _U1430_out;
assign out[0] = _U1429_out;
endmodule

module array_delay_U1421 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1422_in;
wire _U1422_clk;
wire [15:0] _U1422_out;
wire [15:0] _U1423_in;
wire _U1423_clk;
wire [15:0] _U1423_out;
wire [15:0] _U1424_in;
wire _U1424_clk;
wire [15:0] _U1424_out;
wire [15:0] _U1425_in;
wire _U1425_clk;
wire [15:0] _U1425_out;
wire [15:0] _U1426_in;
wire _U1426_clk;
wire [15:0] _U1426_out;
assign _U1422_in = in[0];
assign _U1422_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1422 (
    .in(_U1422_in),
    .clk(_U1422_clk),
    .out(_U1422_out)
);
assign _U1423_in = in[1];
assign _U1423_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1423 (
    .in(_U1423_in),
    .clk(_U1423_clk),
    .out(_U1423_out)
);
assign _U1424_in = in[2];
assign _U1424_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1424 (
    .in(_U1424_in),
    .clk(_U1424_clk),
    .out(_U1424_out)
);
assign _U1425_in = in[3];
assign _U1425_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1425 (
    .in(_U1425_in),
    .clk(_U1425_clk),
    .out(_U1425_out)
);
assign _U1426_in = in[4];
assign _U1426_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1426 (
    .in(_U1426_in),
    .clk(_U1426_clk),
    .out(_U1426_out)
);
assign out[4] = _U1426_out;
assign out[3] = _U1425_out;
assign out[2] = _U1424_out;
assign out[1] = _U1423_out;
assign out[0] = _U1422_out;
endmodule

module array_delay_U1414 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1415_in;
wire _U1415_clk;
wire [15:0] _U1415_out;
wire [15:0] _U1416_in;
wire _U1416_clk;
wire [15:0] _U1416_out;
wire [15:0] _U1417_in;
wire _U1417_clk;
wire [15:0] _U1417_out;
wire [15:0] _U1418_in;
wire _U1418_clk;
wire [15:0] _U1418_out;
wire [15:0] _U1419_in;
wire _U1419_clk;
wire [15:0] _U1419_out;
assign _U1415_in = in[0];
assign _U1415_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1415 (
    .in(_U1415_in),
    .clk(_U1415_clk),
    .out(_U1415_out)
);
assign _U1416_in = in[1];
assign _U1416_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1416 (
    .in(_U1416_in),
    .clk(_U1416_clk),
    .out(_U1416_out)
);
assign _U1417_in = in[2];
assign _U1417_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1417 (
    .in(_U1417_in),
    .clk(_U1417_clk),
    .out(_U1417_out)
);
assign _U1418_in = in[3];
assign _U1418_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1418 (
    .in(_U1418_in),
    .clk(_U1418_clk),
    .out(_U1418_out)
);
assign _U1419_in = in[4];
assign _U1419_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1419 (
    .in(_U1419_in),
    .clk(_U1419_clk),
    .out(_U1419_out)
);
assign out[4] = _U1419_out;
assign out[3] = _U1418_out;
assign out[2] = _U1417_out;
assign out[1] = _U1416_out;
assign out[0] = _U1415_out;
endmodule

module array_delay_U1388 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1389_in;
wire _U1389_clk;
wire [15:0] _U1389_out;
wire [15:0] _U1390_in;
wire _U1390_clk;
wire [15:0] _U1390_out;
wire [15:0] _U1391_in;
wire _U1391_clk;
wire [15:0] _U1391_out;
wire [15:0] _U1392_in;
wire _U1392_clk;
wire [15:0] _U1392_out;
wire [15:0] _U1393_in;
wire _U1393_clk;
wire [15:0] _U1393_out;
assign _U1389_in = in[0];
assign _U1389_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1389 (
    .in(_U1389_in),
    .clk(_U1389_clk),
    .out(_U1389_out)
);
assign _U1390_in = in[1];
assign _U1390_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1390 (
    .in(_U1390_in),
    .clk(_U1390_clk),
    .out(_U1390_out)
);
assign _U1391_in = in[2];
assign _U1391_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1391 (
    .in(_U1391_in),
    .clk(_U1391_clk),
    .out(_U1391_out)
);
assign _U1392_in = in[3];
assign _U1392_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1392 (
    .in(_U1392_in),
    .clk(_U1392_clk),
    .out(_U1392_out)
);
assign _U1393_in = in[4];
assign _U1393_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1393 (
    .in(_U1393_in),
    .clk(_U1393_clk),
    .out(_U1393_out)
);
assign out[4] = _U1393_out;
assign out[3] = _U1392_out;
assign out[2] = _U1391_out;
assign out[1] = _U1390_out;
assign out[0] = _U1389_out;
endmodule

module array_delay_U1381 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1382_in;
wire _U1382_clk;
wire [15:0] _U1382_out;
wire [15:0] _U1383_in;
wire _U1383_clk;
wire [15:0] _U1383_out;
wire [15:0] _U1384_in;
wire _U1384_clk;
wire [15:0] _U1384_out;
wire [15:0] _U1385_in;
wire _U1385_clk;
wire [15:0] _U1385_out;
wire [15:0] _U1386_in;
wire _U1386_clk;
wire [15:0] _U1386_out;
assign _U1382_in = in[0];
assign _U1382_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1382 (
    .in(_U1382_in),
    .clk(_U1382_clk),
    .out(_U1382_out)
);
assign _U1383_in = in[1];
assign _U1383_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1383 (
    .in(_U1383_in),
    .clk(_U1383_clk),
    .out(_U1383_out)
);
assign _U1384_in = in[2];
assign _U1384_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1384 (
    .in(_U1384_in),
    .clk(_U1384_clk),
    .out(_U1384_out)
);
assign _U1385_in = in[3];
assign _U1385_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1385 (
    .in(_U1385_in),
    .clk(_U1385_clk),
    .out(_U1385_out)
);
assign _U1386_in = in[4];
assign _U1386_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1386 (
    .in(_U1386_in),
    .clk(_U1386_clk),
    .out(_U1386_out)
);
assign out[4] = _U1386_out;
assign out[3] = _U1385_out;
assign out[2] = _U1384_out;
assign out[1] = _U1383_out;
assign out[0] = _U1382_out;
endmodule

module array_delay_U1338 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1339_in;
wire _U1339_clk;
wire [15:0] _U1339_out;
wire [15:0] _U1340_in;
wire _U1340_clk;
wire [15:0] _U1340_out;
wire [15:0] _U1341_in;
wire _U1341_clk;
wire [15:0] _U1341_out;
wire [15:0] _U1342_in;
wire _U1342_clk;
wire [15:0] _U1342_out;
wire [15:0] _U1343_in;
wire _U1343_clk;
wire [15:0] _U1343_out;
assign _U1339_in = in[0];
assign _U1339_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1339 (
    .in(_U1339_in),
    .clk(_U1339_clk),
    .out(_U1339_out)
);
assign _U1340_in = in[1];
assign _U1340_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1340 (
    .in(_U1340_in),
    .clk(_U1340_clk),
    .out(_U1340_out)
);
assign _U1341_in = in[2];
assign _U1341_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1341 (
    .in(_U1341_in),
    .clk(_U1341_clk),
    .out(_U1341_out)
);
assign _U1342_in = in[3];
assign _U1342_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1342 (
    .in(_U1342_in),
    .clk(_U1342_clk),
    .out(_U1342_out)
);
assign _U1343_in = in[4];
assign _U1343_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1343 (
    .in(_U1343_in),
    .clk(_U1343_clk),
    .out(_U1343_out)
);
assign out[4] = _U1343_out;
assign out[3] = _U1342_out;
assign out[2] = _U1341_out;
assign out[1] = _U1340_out;
assign out[0] = _U1339_out;
endmodule

module array_delay_U1331 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1332_in;
wire _U1332_clk;
wire [15:0] _U1332_out;
wire [15:0] _U1333_in;
wire _U1333_clk;
wire [15:0] _U1333_out;
wire [15:0] _U1334_in;
wire _U1334_clk;
wire [15:0] _U1334_out;
wire [15:0] _U1335_in;
wire _U1335_clk;
wire [15:0] _U1335_out;
wire [15:0] _U1336_in;
wire _U1336_clk;
wire [15:0] _U1336_out;
assign _U1332_in = in[0];
assign _U1332_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1332 (
    .in(_U1332_in),
    .clk(_U1332_clk),
    .out(_U1332_out)
);
assign _U1333_in = in[1];
assign _U1333_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1333 (
    .in(_U1333_in),
    .clk(_U1333_clk),
    .out(_U1333_out)
);
assign _U1334_in = in[2];
assign _U1334_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1334 (
    .in(_U1334_in),
    .clk(_U1334_clk),
    .out(_U1334_out)
);
assign _U1335_in = in[3];
assign _U1335_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1335 (
    .in(_U1335_in),
    .clk(_U1335_clk),
    .out(_U1335_out)
);
assign _U1336_in = in[4];
assign _U1336_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1336 (
    .in(_U1336_in),
    .clk(_U1336_clk),
    .out(_U1336_out)
);
assign out[4] = _U1336_out;
assign out[3] = _U1335_out;
assign out[2] = _U1334_out;
assign out[1] = _U1333_out;
assign out[0] = _U1332_out;
endmodule

module array_delay_U1324 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1325_in;
wire _U1325_clk;
wire [15:0] _U1325_out;
wire [15:0] _U1326_in;
wire _U1326_clk;
wire [15:0] _U1326_out;
wire [15:0] _U1327_in;
wire _U1327_clk;
wire [15:0] _U1327_out;
wire [15:0] _U1328_in;
wire _U1328_clk;
wire [15:0] _U1328_out;
wire [15:0] _U1329_in;
wire _U1329_clk;
wire [15:0] _U1329_out;
assign _U1325_in = in[0];
assign _U1325_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1325 (
    .in(_U1325_in),
    .clk(_U1325_clk),
    .out(_U1325_out)
);
assign _U1326_in = in[1];
assign _U1326_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1326 (
    .in(_U1326_in),
    .clk(_U1326_clk),
    .out(_U1326_out)
);
assign _U1327_in = in[2];
assign _U1327_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1327 (
    .in(_U1327_in),
    .clk(_U1327_clk),
    .out(_U1327_out)
);
assign _U1328_in = in[3];
assign _U1328_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1328 (
    .in(_U1328_in),
    .clk(_U1328_clk),
    .out(_U1328_out)
);
assign _U1329_in = in[4];
assign _U1329_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1329 (
    .in(_U1329_in),
    .clk(_U1329_clk),
    .out(_U1329_out)
);
assign out[4] = _U1329_out;
assign out[3] = _U1328_out;
assign out[2] = _U1327_out;
assign out[1] = _U1326_out;
assign out[0] = _U1325_out;
endmodule

module array_delay_U1317 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1318_in;
wire _U1318_clk;
wire [15:0] _U1318_out;
wire [15:0] _U1319_in;
wire _U1319_clk;
wire [15:0] _U1319_out;
wire [15:0] _U1320_in;
wire _U1320_clk;
wire [15:0] _U1320_out;
wire [15:0] _U1321_in;
wire _U1321_clk;
wire [15:0] _U1321_out;
wire [15:0] _U1322_in;
wire _U1322_clk;
wire [15:0] _U1322_out;
assign _U1318_in = in[0];
assign _U1318_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1318 (
    .in(_U1318_in),
    .clk(_U1318_clk),
    .out(_U1318_out)
);
assign _U1319_in = in[1];
assign _U1319_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1319 (
    .in(_U1319_in),
    .clk(_U1319_clk),
    .out(_U1319_out)
);
assign _U1320_in = in[2];
assign _U1320_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1320 (
    .in(_U1320_in),
    .clk(_U1320_clk),
    .out(_U1320_out)
);
assign _U1321_in = in[3];
assign _U1321_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1321 (
    .in(_U1321_in),
    .clk(_U1321_clk),
    .out(_U1321_out)
);
assign _U1322_in = in[4];
assign _U1322_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1322 (
    .in(_U1322_in),
    .clk(_U1322_clk),
    .out(_U1322_out)
);
assign out[4] = _U1322_out;
assign out[3] = _U1321_out;
assign out[2] = _U1320_out;
assign out[1] = _U1319_out;
assign out[0] = _U1318_out;
endmodule

module array_delay_U1310 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1311_in;
wire _U1311_clk;
wire [15:0] _U1311_out;
wire [15:0] _U1312_in;
wire _U1312_clk;
wire [15:0] _U1312_out;
wire [15:0] _U1313_in;
wire _U1313_clk;
wire [15:0] _U1313_out;
wire [15:0] _U1314_in;
wire _U1314_clk;
wire [15:0] _U1314_out;
wire [15:0] _U1315_in;
wire _U1315_clk;
wire [15:0] _U1315_out;
assign _U1311_in = in[0];
assign _U1311_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1311 (
    .in(_U1311_in),
    .clk(_U1311_clk),
    .out(_U1311_out)
);
assign _U1312_in = in[1];
assign _U1312_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1312 (
    .in(_U1312_in),
    .clk(_U1312_clk),
    .out(_U1312_out)
);
assign _U1313_in = in[2];
assign _U1313_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1313 (
    .in(_U1313_in),
    .clk(_U1313_clk),
    .out(_U1313_out)
);
assign _U1314_in = in[3];
assign _U1314_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1314 (
    .in(_U1314_in),
    .clk(_U1314_clk),
    .out(_U1314_out)
);
assign _U1315_in = in[4];
assign _U1315_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1315 (
    .in(_U1315_in),
    .clk(_U1315_clk),
    .out(_U1315_out)
);
assign out[4] = _U1315_out;
assign out[3] = _U1314_out;
assign out[2] = _U1313_out;
assign out[1] = _U1312_out;
assign out[0] = _U1311_out;
endmodule

module array_delay_U1303 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1304_in;
wire _U1304_clk;
wire [15:0] _U1304_out;
wire [15:0] _U1305_in;
wire _U1305_clk;
wire [15:0] _U1305_out;
wire [15:0] _U1306_in;
wire _U1306_clk;
wire [15:0] _U1306_out;
wire [15:0] _U1307_in;
wire _U1307_clk;
wire [15:0] _U1307_out;
wire [15:0] _U1308_in;
wire _U1308_clk;
wire [15:0] _U1308_out;
assign _U1304_in = in[0];
assign _U1304_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1304 (
    .in(_U1304_in),
    .clk(_U1304_clk),
    .out(_U1304_out)
);
assign _U1305_in = in[1];
assign _U1305_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1305 (
    .in(_U1305_in),
    .clk(_U1305_clk),
    .out(_U1305_out)
);
assign _U1306_in = in[2];
assign _U1306_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1306 (
    .in(_U1306_in),
    .clk(_U1306_clk),
    .out(_U1306_out)
);
assign _U1307_in = in[3];
assign _U1307_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1307 (
    .in(_U1307_in),
    .clk(_U1307_clk),
    .out(_U1307_out)
);
assign _U1308_in = in[4];
assign _U1308_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1308 (
    .in(_U1308_in),
    .clk(_U1308_clk),
    .out(_U1308_out)
);
assign out[4] = _U1308_out;
assign out[3] = _U1307_out;
assign out[2] = _U1306_out;
assign out[1] = _U1305_out;
assign out[0] = _U1304_out;
endmodule

module array_delay_U1296 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1297_in;
wire _U1297_clk;
wire [15:0] _U1297_out;
wire [15:0] _U1298_in;
wire _U1298_clk;
wire [15:0] _U1298_out;
wire [15:0] _U1299_in;
wire _U1299_clk;
wire [15:0] _U1299_out;
wire [15:0] _U1300_in;
wire _U1300_clk;
wire [15:0] _U1300_out;
wire [15:0] _U1301_in;
wire _U1301_clk;
wire [15:0] _U1301_out;
assign _U1297_in = in[0];
assign _U1297_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1297 (
    .in(_U1297_in),
    .clk(_U1297_clk),
    .out(_U1297_out)
);
assign _U1298_in = in[1];
assign _U1298_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1298 (
    .in(_U1298_in),
    .clk(_U1298_clk),
    .out(_U1298_out)
);
assign _U1299_in = in[2];
assign _U1299_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1299 (
    .in(_U1299_in),
    .clk(_U1299_clk),
    .out(_U1299_out)
);
assign _U1300_in = in[3];
assign _U1300_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1300 (
    .in(_U1300_in),
    .clk(_U1300_clk),
    .out(_U1300_out)
);
assign _U1301_in = in[4];
assign _U1301_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1301 (
    .in(_U1301_in),
    .clk(_U1301_clk),
    .out(_U1301_out)
);
assign out[4] = _U1301_out;
assign out[3] = _U1300_out;
assign out[2] = _U1299_out;
assign out[1] = _U1298_out;
assign out[0] = _U1297_out;
endmodule

module array_delay_U1289 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1290_in;
wire _U1290_clk;
wire [15:0] _U1290_out;
wire [15:0] _U1291_in;
wire _U1291_clk;
wire [15:0] _U1291_out;
wire [15:0] _U1292_in;
wire _U1292_clk;
wire [15:0] _U1292_out;
wire [15:0] _U1293_in;
wire _U1293_clk;
wire [15:0] _U1293_out;
wire [15:0] _U1294_in;
wire _U1294_clk;
wire [15:0] _U1294_out;
assign _U1290_in = in[0];
assign _U1290_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1290 (
    .in(_U1290_in),
    .clk(_U1290_clk),
    .out(_U1290_out)
);
assign _U1291_in = in[1];
assign _U1291_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1291 (
    .in(_U1291_in),
    .clk(_U1291_clk),
    .out(_U1291_out)
);
assign _U1292_in = in[2];
assign _U1292_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1292 (
    .in(_U1292_in),
    .clk(_U1292_clk),
    .out(_U1292_out)
);
assign _U1293_in = in[3];
assign _U1293_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1293 (
    .in(_U1293_in),
    .clk(_U1293_clk),
    .out(_U1293_out)
);
assign _U1294_in = in[4];
assign _U1294_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1294 (
    .in(_U1294_in),
    .clk(_U1294_clk),
    .out(_U1294_out)
);
assign out[4] = _U1294_out;
assign out[3] = _U1293_out;
assign out[2] = _U1292_out;
assign out[1] = _U1291_out;
assign out[0] = _U1290_out;
endmodule

module array_delay_U1282 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1283_in;
wire _U1283_clk;
wire [15:0] _U1283_out;
wire [15:0] _U1284_in;
wire _U1284_clk;
wire [15:0] _U1284_out;
wire [15:0] _U1285_in;
wire _U1285_clk;
wire [15:0] _U1285_out;
wire [15:0] _U1286_in;
wire _U1286_clk;
wire [15:0] _U1286_out;
wire [15:0] _U1287_in;
wire _U1287_clk;
wire [15:0] _U1287_out;
assign _U1283_in = in[0];
assign _U1283_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1283 (
    .in(_U1283_in),
    .clk(_U1283_clk),
    .out(_U1283_out)
);
assign _U1284_in = in[1];
assign _U1284_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1284 (
    .in(_U1284_in),
    .clk(_U1284_clk),
    .out(_U1284_out)
);
assign _U1285_in = in[2];
assign _U1285_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1285 (
    .in(_U1285_in),
    .clk(_U1285_clk),
    .out(_U1285_out)
);
assign _U1286_in = in[3];
assign _U1286_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1286 (
    .in(_U1286_in),
    .clk(_U1286_clk),
    .out(_U1286_out)
);
assign _U1287_in = in[4];
assign _U1287_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1287 (
    .in(_U1287_in),
    .clk(_U1287_clk),
    .out(_U1287_out)
);
assign out[4] = _U1287_out;
assign out[3] = _U1286_out;
assign out[2] = _U1285_out;
assign out[1] = _U1284_out;
assign out[0] = _U1283_out;
endmodule

module array_delay_U1275 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1276_in;
wire _U1276_clk;
wire [15:0] _U1276_out;
wire [15:0] _U1277_in;
wire _U1277_clk;
wire [15:0] _U1277_out;
wire [15:0] _U1278_in;
wire _U1278_clk;
wire [15:0] _U1278_out;
wire [15:0] _U1279_in;
wire _U1279_clk;
wire [15:0] _U1279_out;
wire [15:0] _U1280_in;
wire _U1280_clk;
wire [15:0] _U1280_out;
assign _U1276_in = in[0];
assign _U1276_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1276 (
    .in(_U1276_in),
    .clk(_U1276_clk),
    .out(_U1276_out)
);
assign _U1277_in = in[1];
assign _U1277_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1277 (
    .in(_U1277_in),
    .clk(_U1277_clk),
    .out(_U1277_out)
);
assign _U1278_in = in[2];
assign _U1278_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1278 (
    .in(_U1278_in),
    .clk(_U1278_clk),
    .out(_U1278_out)
);
assign _U1279_in = in[3];
assign _U1279_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1279 (
    .in(_U1279_in),
    .clk(_U1279_clk),
    .out(_U1279_out)
);
assign _U1280_in = in[4];
assign _U1280_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1280 (
    .in(_U1280_in),
    .clk(_U1280_clk),
    .out(_U1280_out)
);
assign out[4] = _U1280_out;
assign out[3] = _U1279_out;
assign out[2] = _U1278_out;
assign out[1] = _U1277_out;
assign out[0] = _U1276_out;
endmodule

module array_delay_U1268 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1269_in;
wire _U1269_clk;
wire [15:0] _U1269_out;
wire [15:0] _U1270_in;
wire _U1270_clk;
wire [15:0] _U1270_out;
wire [15:0] _U1271_in;
wire _U1271_clk;
wire [15:0] _U1271_out;
wire [15:0] _U1272_in;
wire _U1272_clk;
wire [15:0] _U1272_out;
wire [15:0] _U1273_in;
wire _U1273_clk;
wire [15:0] _U1273_out;
assign _U1269_in = in[0];
assign _U1269_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1269 (
    .in(_U1269_in),
    .clk(_U1269_clk),
    .out(_U1269_out)
);
assign _U1270_in = in[1];
assign _U1270_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1270 (
    .in(_U1270_in),
    .clk(_U1270_clk),
    .out(_U1270_out)
);
assign _U1271_in = in[2];
assign _U1271_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1271 (
    .in(_U1271_in),
    .clk(_U1271_clk),
    .out(_U1271_out)
);
assign _U1272_in = in[3];
assign _U1272_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1272 (
    .in(_U1272_in),
    .clk(_U1272_clk),
    .out(_U1272_out)
);
assign _U1273_in = in[4];
assign _U1273_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1273 (
    .in(_U1273_in),
    .clk(_U1273_clk),
    .out(_U1273_out)
);
assign out[4] = _U1273_out;
assign out[3] = _U1272_out;
assign out[2] = _U1271_out;
assign out[1] = _U1270_out;
assign out[0] = _U1269_out;
endmodule

module array_delay_U1261 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1262_in;
wire _U1262_clk;
wire [15:0] _U1262_out;
wire [15:0] _U1263_in;
wire _U1263_clk;
wire [15:0] _U1263_out;
wire [15:0] _U1264_in;
wire _U1264_clk;
wire [15:0] _U1264_out;
wire [15:0] _U1265_in;
wire _U1265_clk;
wire [15:0] _U1265_out;
wire [15:0] _U1266_in;
wire _U1266_clk;
wire [15:0] _U1266_out;
assign _U1262_in = in[0];
assign _U1262_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1262 (
    .in(_U1262_in),
    .clk(_U1262_clk),
    .out(_U1262_out)
);
assign _U1263_in = in[1];
assign _U1263_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1263 (
    .in(_U1263_in),
    .clk(_U1263_clk),
    .out(_U1263_out)
);
assign _U1264_in = in[2];
assign _U1264_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1264 (
    .in(_U1264_in),
    .clk(_U1264_clk),
    .out(_U1264_out)
);
assign _U1265_in = in[3];
assign _U1265_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1265 (
    .in(_U1265_in),
    .clk(_U1265_clk),
    .out(_U1265_out)
);
assign _U1266_in = in[4];
assign _U1266_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1266 (
    .in(_U1266_in),
    .clk(_U1266_clk),
    .out(_U1266_out)
);
assign out[4] = _U1266_out;
assign out[3] = _U1265_out;
assign out[2] = _U1264_out;
assign out[1] = _U1263_out;
assign out[0] = _U1262_out;
endmodule

module array_delay_U1254 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1255_in;
wire _U1255_clk;
wire [15:0] _U1255_out;
wire [15:0] _U1256_in;
wire _U1256_clk;
wire [15:0] _U1256_out;
wire [15:0] _U1257_in;
wire _U1257_clk;
wire [15:0] _U1257_out;
wire [15:0] _U1258_in;
wire _U1258_clk;
wire [15:0] _U1258_out;
wire [15:0] _U1259_in;
wire _U1259_clk;
wire [15:0] _U1259_out;
assign _U1255_in = in[0];
assign _U1255_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1255 (
    .in(_U1255_in),
    .clk(_U1255_clk),
    .out(_U1255_out)
);
assign _U1256_in = in[1];
assign _U1256_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1256 (
    .in(_U1256_in),
    .clk(_U1256_clk),
    .out(_U1256_out)
);
assign _U1257_in = in[2];
assign _U1257_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1257 (
    .in(_U1257_in),
    .clk(_U1257_clk),
    .out(_U1257_out)
);
assign _U1258_in = in[3];
assign _U1258_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1258 (
    .in(_U1258_in),
    .clk(_U1258_clk),
    .out(_U1258_out)
);
assign _U1259_in = in[4];
assign _U1259_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1259 (
    .in(_U1259_in),
    .clk(_U1259_clk),
    .out(_U1259_out)
);
assign out[4] = _U1259_out;
assign out[3] = _U1258_out;
assign out[2] = _U1257_out;
assign out[1] = _U1256_out;
assign out[0] = _U1255_out;
endmodule

module array_delay_U1247 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1248_in;
wire _U1248_clk;
wire [15:0] _U1248_out;
wire [15:0] _U1249_in;
wire _U1249_clk;
wire [15:0] _U1249_out;
wire [15:0] _U1250_in;
wire _U1250_clk;
wire [15:0] _U1250_out;
wire [15:0] _U1251_in;
wire _U1251_clk;
wire [15:0] _U1251_out;
wire [15:0] _U1252_in;
wire _U1252_clk;
wire [15:0] _U1252_out;
assign _U1248_in = in[0];
assign _U1248_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1248 (
    .in(_U1248_in),
    .clk(_U1248_clk),
    .out(_U1248_out)
);
assign _U1249_in = in[1];
assign _U1249_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1249 (
    .in(_U1249_in),
    .clk(_U1249_clk),
    .out(_U1249_out)
);
assign _U1250_in = in[2];
assign _U1250_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1250 (
    .in(_U1250_in),
    .clk(_U1250_clk),
    .out(_U1250_out)
);
assign _U1251_in = in[3];
assign _U1251_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1251 (
    .in(_U1251_in),
    .clk(_U1251_clk),
    .out(_U1251_out)
);
assign _U1252_in = in[4];
assign _U1252_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1252 (
    .in(_U1252_in),
    .clk(_U1252_clk),
    .out(_U1252_out)
);
assign out[4] = _U1252_out;
assign out[3] = _U1251_out;
assign out[2] = _U1250_out;
assign out[1] = _U1249_out;
assign out[0] = _U1248_out;
endmodule

module array_delay_U1240 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1241_in;
wire _U1241_clk;
wire [15:0] _U1241_out;
wire [15:0] _U1242_in;
wire _U1242_clk;
wire [15:0] _U1242_out;
wire [15:0] _U1243_in;
wire _U1243_clk;
wire [15:0] _U1243_out;
wire [15:0] _U1244_in;
wire _U1244_clk;
wire [15:0] _U1244_out;
wire [15:0] _U1245_in;
wire _U1245_clk;
wire [15:0] _U1245_out;
assign _U1241_in = in[0];
assign _U1241_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1241 (
    .in(_U1241_in),
    .clk(_U1241_clk),
    .out(_U1241_out)
);
assign _U1242_in = in[1];
assign _U1242_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1242 (
    .in(_U1242_in),
    .clk(_U1242_clk),
    .out(_U1242_out)
);
assign _U1243_in = in[2];
assign _U1243_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1243 (
    .in(_U1243_in),
    .clk(_U1243_clk),
    .out(_U1243_out)
);
assign _U1244_in = in[3];
assign _U1244_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1244 (
    .in(_U1244_in),
    .clk(_U1244_clk),
    .out(_U1244_out)
);
assign _U1245_in = in[4];
assign _U1245_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1245 (
    .in(_U1245_in),
    .clk(_U1245_clk),
    .out(_U1245_out)
);
assign out[4] = _U1245_out;
assign out[3] = _U1244_out;
assign out[2] = _U1243_out;
assign out[1] = _U1242_out;
assign out[0] = _U1241_out;
endmodule

module array_delay_U1233 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1234_in;
wire _U1234_clk;
wire [15:0] _U1234_out;
wire [15:0] _U1235_in;
wire _U1235_clk;
wire [15:0] _U1235_out;
wire [15:0] _U1236_in;
wire _U1236_clk;
wire [15:0] _U1236_out;
wire [15:0] _U1237_in;
wire _U1237_clk;
wire [15:0] _U1237_out;
wire [15:0] _U1238_in;
wire _U1238_clk;
wire [15:0] _U1238_out;
assign _U1234_in = in[0];
assign _U1234_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1234 (
    .in(_U1234_in),
    .clk(_U1234_clk),
    .out(_U1234_out)
);
assign _U1235_in = in[1];
assign _U1235_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1235 (
    .in(_U1235_in),
    .clk(_U1235_clk),
    .out(_U1235_out)
);
assign _U1236_in = in[2];
assign _U1236_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1236 (
    .in(_U1236_in),
    .clk(_U1236_clk),
    .out(_U1236_out)
);
assign _U1237_in = in[3];
assign _U1237_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1237 (
    .in(_U1237_in),
    .clk(_U1237_clk),
    .out(_U1237_out)
);
assign _U1238_in = in[4];
assign _U1238_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1238 (
    .in(_U1238_in),
    .clk(_U1238_clk),
    .out(_U1238_out)
);
assign out[4] = _U1238_out;
assign out[3] = _U1237_out;
assign out[2] = _U1236_out;
assign out[1] = _U1235_out;
assign out[0] = _U1234_out;
endmodule

module array_delay_U1226 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1227_in;
wire _U1227_clk;
wire [15:0] _U1227_out;
wire [15:0] _U1228_in;
wire _U1228_clk;
wire [15:0] _U1228_out;
wire [15:0] _U1229_in;
wire _U1229_clk;
wire [15:0] _U1229_out;
wire [15:0] _U1230_in;
wire _U1230_clk;
wire [15:0] _U1230_out;
wire [15:0] _U1231_in;
wire _U1231_clk;
wire [15:0] _U1231_out;
assign _U1227_in = in[0];
assign _U1227_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1227 (
    .in(_U1227_in),
    .clk(_U1227_clk),
    .out(_U1227_out)
);
assign _U1228_in = in[1];
assign _U1228_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1228 (
    .in(_U1228_in),
    .clk(_U1228_clk),
    .out(_U1228_out)
);
assign _U1229_in = in[2];
assign _U1229_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1229 (
    .in(_U1229_in),
    .clk(_U1229_clk),
    .out(_U1229_out)
);
assign _U1230_in = in[3];
assign _U1230_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1230 (
    .in(_U1230_in),
    .clk(_U1230_clk),
    .out(_U1230_out)
);
assign _U1231_in = in[4];
assign _U1231_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1231 (
    .in(_U1231_in),
    .clk(_U1231_clk),
    .out(_U1231_out)
);
assign out[4] = _U1231_out;
assign out[3] = _U1230_out;
assign out[2] = _U1229_out;
assign out[1] = _U1228_out;
assign out[0] = _U1227_out;
endmodule

module array_delay_U1200 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1201_in;
wire _U1201_clk;
wire [15:0] _U1201_out;
wire [15:0] _U1202_in;
wire _U1202_clk;
wire [15:0] _U1202_out;
wire [15:0] _U1203_in;
wire _U1203_clk;
wire [15:0] _U1203_out;
wire [15:0] _U1204_in;
wire _U1204_clk;
wire [15:0] _U1204_out;
wire [15:0] _U1205_in;
wire _U1205_clk;
wire [15:0] _U1205_out;
assign _U1201_in = in[0];
assign _U1201_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1201 (
    .in(_U1201_in),
    .clk(_U1201_clk),
    .out(_U1201_out)
);
assign _U1202_in = in[1];
assign _U1202_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1202 (
    .in(_U1202_in),
    .clk(_U1202_clk),
    .out(_U1202_out)
);
assign _U1203_in = in[2];
assign _U1203_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1203 (
    .in(_U1203_in),
    .clk(_U1203_clk),
    .out(_U1203_out)
);
assign _U1204_in = in[3];
assign _U1204_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1204 (
    .in(_U1204_in),
    .clk(_U1204_clk),
    .out(_U1204_out)
);
assign _U1205_in = in[4];
assign _U1205_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1205 (
    .in(_U1205_in),
    .clk(_U1205_clk),
    .out(_U1205_out)
);
assign out[4] = _U1205_out;
assign out[3] = _U1204_out;
assign out[2] = _U1203_out;
assign out[1] = _U1202_out;
assign out[0] = _U1201_out;
endmodule

module array_delay_U1193 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1194_in;
wire _U1194_clk;
wire [15:0] _U1194_out;
wire [15:0] _U1195_in;
wire _U1195_clk;
wire [15:0] _U1195_out;
wire [15:0] _U1196_in;
wire _U1196_clk;
wire [15:0] _U1196_out;
wire [15:0] _U1197_in;
wire _U1197_clk;
wire [15:0] _U1197_out;
wire [15:0] _U1198_in;
wire _U1198_clk;
wire [15:0] _U1198_out;
assign _U1194_in = in[0];
assign _U1194_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1194 (
    .in(_U1194_in),
    .clk(_U1194_clk),
    .out(_U1194_out)
);
assign _U1195_in = in[1];
assign _U1195_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1195 (
    .in(_U1195_in),
    .clk(_U1195_clk),
    .out(_U1195_out)
);
assign _U1196_in = in[2];
assign _U1196_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1196 (
    .in(_U1196_in),
    .clk(_U1196_clk),
    .out(_U1196_out)
);
assign _U1197_in = in[3];
assign _U1197_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1197 (
    .in(_U1197_in),
    .clk(_U1197_clk),
    .out(_U1197_out)
);
assign _U1198_in = in[4];
assign _U1198_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1198 (
    .in(_U1198_in),
    .clk(_U1198_clk),
    .out(_U1198_out)
);
assign out[4] = _U1198_out;
assign out[3] = _U1197_out;
assign out[2] = _U1196_out;
assign out[1] = _U1195_out;
assign out[0] = _U1194_out;
endmodule

module array_delay_U1150 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1151_in;
wire _U1151_clk;
wire [15:0] _U1151_out;
wire [15:0] _U1152_in;
wire _U1152_clk;
wire [15:0] _U1152_out;
wire [15:0] _U1153_in;
wire _U1153_clk;
wire [15:0] _U1153_out;
wire [15:0] _U1154_in;
wire _U1154_clk;
wire [15:0] _U1154_out;
wire [15:0] _U1155_in;
wire _U1155_clk;
wire [15:0] _U1155_out;
assign _U1151_in = in[0];
assign _U1151_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1151 (
    .in(_U1151_in),
    .clk(_U1151_clk),
    .out(_U1151_out)
);
assign _U1152_in = in[1];
assign _U1152_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1152 (
    .in(_U1152_in),
    .clk(_U1152_clk),
    .out(_U1152_out)
);
assign _U1153_in = in[2];
assign _U1153_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1153 (
    .in(_U1153_in),
    .clk(_U1153_clk),
    .out(_U1153_out)
);
assign _U1154_in = in[3];
assign _U1154_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1154 (
    .in(_U1154_in),
    .clk(_U1154_clk),
    .out(_U1154_out)
);
assign _U1155_in = in[4];
assign _U1155_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1155 (
    .in(_U1155_in),
    .clk(_U1155_clk),
    .out(_U1155_out)
);
assign out[4] = _U1155_out;
assign out[3] = _U1154_out;
assign out[2] = _U1153_out;
assign out[1] = _U1152_out;
assign out[0] = _U1151_out;
endmodule

module array_delay_U1143 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1144_in;
wire _U1144_clk;
wire [15:0] _U1144_out;
wire [15:0] _U1145_in;
wire _U1145_clk;
wire [15:0] _U1145_out;
wire [15:0] _U1146_in;
wire _U1146_clk;
wire [15:0] _U1146_out;
wire [15:0] _U1147_in;
wire _U1147_clk;
wire [15:0] _U1147_out;
wire [15:0] _U1148_in;
wire _U1148_clk;
wire [15:0] _U1148_out;
assign _U1144_in = in[0];
assign _U1144_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1144 (
    .in(_U1144_in),
    .clk(_U1144_clk),
    .out(_U1144_out)
);
assign _U1145_in = in[1];
assign _U1145_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1145 (
    .in(_U1145_in),
    .clk(_U1145_clk),
    .out(_U1145_out)
);
assign _U1146_in = in[2];
assign _U1146_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1146 (
    .in(_U1146_in),
    .clk(_U1146_clk),
    .out(_U1146_out)
);
assign _U1147_in = in[3];
assign _U1147_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1147 (
    .in(_U1147_in),
    .clk(_U1147_clk),
    .out(_U1147_out)
);
assign _U1148_in = in[4];
assign _U1148_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1148 (
    .in(_U1148_in),
    .clk(_U1148_clk),
    .out(_U1148_out)
);
assign out[4] = _U1148_out;
assign out[3] = _U1147_out;
assign out[2] = _U1146_out;
assign out[1] = _U1145_out;
assign out[0] = _U1144_out;
endmodule

module array_delay_U1136 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1137_in;
wire _U1137_clk;
wire [15:0] _U1137_out;
wire [15:0] _U1138_in;
wire _U1138_clk;
wire [15:0] _U1138_out;
wire [15:0] _U1139_in;
wire _U1139_clk;
wire [15:0] _U1139_out;
wire [15:0] _U1140_in;
wire _U1140_clk;
wire [15:0] _U1140_out;
wire [15:0] _U1141_in;
wire _U1141_clk;
wire [15:0] _U1141_out;
assign _U1137_in = in[0];
assign _U1137_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1137 (
    .in(_U1137_in),
    .clk(_U1137_clk),
    .out(_U1137_out)
);
assign _U1138_in = in[1];
assign _U1138_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1138 (
    .in(_U1138_in),
    .clk(_U1138_clk),
    .out(_U1138_out)
);
assign _U1139_in = in[2];
assign _U1139_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1139 (
    .in(_U1139_in),
    .clk(_U1139_clk),
    .out(_U1139_out)
);
assign _U1140_in = in[3];
assign _U1140_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1140 (
    .in(_U1140_in),
    .clk(_U1140_clk),
    .out(_U1140_out)
);
assign _U1141_in = in[4];
assign _U1141_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1141 (
    .in(_U1141_in),
    .clk(_U1141_clk),
    .out(_U1141_out)
);
assign out[4] = _U1141_out;
assign out[3] = _U1140_out;
assign out[2] = _U1139_out;
assign out[1] = _U1138_out;
assign out[0] = _U1137_out;
endmodule

module array_delay_U1129 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1130_in;
wire _U1130_clk;
wire [15:0] _U1130_out;
wire [15:0] _U1131_in;
wire _U1131_clk;
wire [15:0] _U1131_out;
wire [15:0] _U1132_in;
wire _U1132_clk;
wire [15:0] _U1132_out;
wire [15:0] _U1133_in;
wire _U1133_clk;
wire [15:0] _U1133_out;
wire [15:0] _U1134_in;
wire _U1134_clk;
wire [15:0] _U1134_out;
assign _U1130_in = in[0];
assign _U1130_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1130 (
    .in(_U1130_in),
    .clk(_U1130_clk),
    .out(_U1130_out)
);
assign _U1131_in = in[1];
assign _U1131_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1131 (
    .in(_U1131_in),
    .clk(_U1131_clk),
    .out(_U1131_out)
);
assign _U1132_in = in[2];
assign _U1132_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1132 (
    .in(_U1132_in),
    .clk(_U1132_clk),
    .out(_U1132_out)
);
assign _U1133_in = in[3];
assign _U1133_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1133 (
    .in(_U1133_in),
    .clk(_U1133_clk),
    .out(_U1133_out)
);
assign _U1134_in = in[4];
assign _U1134_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1134 (
    .in(_U1134_in),
    .clk(_U1134_clk),
    .out(_U1134_out)
);
assign out[4] = _U1134_out;
assign out[3] = _U1133_out;
assign out[2] = _U1132_out;
assign out[1] = _U1131_out;
assign out[0] = _U1130_out;
endmodule

module array_delay_U1122 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1123_in;
wire _U1123_clk;
wire [15:0] _U1123_out;
wire [15:0] _U1124_in;
wire _U1124_clk;
wire [15:0] _U1124_out;
wire [15:0] _U1125_in;
wire _U1125_clk;
wire [15:0] _U1125_out;
wire [15:0] _U1126_in;
wire _U1126_clk;
wire [15:0] _U1126_out;
wire [15:0] _U1127_in;
wire _U1127_clk;
wire [15:0] _U1127_out;
assign _U1123_in = in[0];
assign _U1123_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1123 (
    .in(_U1123_in),
    .clk(_U1123_clk),
    .out(_U1123_out)
);
assign _U1124_in = in[1];
assign _U1124_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1124 (
    .in(_U1124_in),
    .clk(_U1124_clk),
    .out(_U1124_out)
);
assign _U1125_in = in[2];
assign _U1125_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1125 (
    .in(_U1125_in),
    .clk(_U1125_clk),
    .out(_U1125_out)
);
assign _U1126_in = in[3];
assign _U1126_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1126 (
    .in(_U1126_in),
    .clk(_U1126_clk),
    .out(_U1126_out)
);
assign _U1127_in = in[4];
assign _U1127_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1127 (
    .in(_U1127_in),
    .clk(_U1127_clk),
    .out(_U1127_out)
);
assign out[4] = _U1127_out;
assign out[3] = _U1126_out;
assign out[2] = _U1125_out;
assign out[1] = _U1124_out;
assign out[0] = _U1123_out;
endmodule

module array_delay_U1115 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1116_in;
wire _U1116_clk;
wire [15:0] _U1116_out;
wire [15:0] _U1117_in;
wire _U1117_clk;
wire [15:0] _U1117_out;
wire [15:0] _U1118_in;
wire _U1118_clk;
wire [15:0] _U1118_out;
wire [15:0] _U1119_in;
wire _U1119_clk;
wire [15:0] _U1119_out;
wire [15:0] _U1120_in;
wire _U1120_clk;
wire [15:0] _U1120_out;
assign _U1116_in = in[0];
assign _U1116_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1116 (
    .in(_U1116_in),
    .clk(_U1116_clk),
    .out(_U1116_out)
);
assign _U1117_in = in[1];
assign _U1117_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1117 (
    .in(_U1117_in),
    .clk(_U1117_clk),
    .out(_U1117_out)
);
assign _U1118_in = in[2];
assign _U1118_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1118 (
    .in(_U1118_in),
    .clk(_U1118_clk),
    .out(_U1118_out)
);
assign _U1119_in = in[3];
assign _U1119_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1119 (
    .in(_U1119_in),
    .clk(_U1119_clk),
    .out(_U1119_out)
);
assign _U1120_in = in[4];
assign _U1120_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1120 (
    .in(_U1120_in),
    .clk(_U1120_clk),
    .out(_U1120_out)
);
assign out[4] = _U1120_out;
assign out[3] = _U1119_out;
assign out[2] = _U1118_out;
assign out[1] = _U1117_out;
assign out[0] = _U1116_out;
endmodule

module array_delay_U1108 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1109_in;
wire _U1109_clk;
wire [15:0] _U1109_out;
wire [15:0] _U1110_in;
wire _U1110_clk;
wire [15:0] _U1110_out;
wire [15:0] _U1111_in;
wire _U1111_clk;
wire [15:0] _U1111_out;
wire [15:0] _U1112_in;
wire _U1112_clk;
wire [15:0] _U1112_out;
wire [15:0] _U1113_in;
wire _U1113_clk;
wire [15:0] _U1113_out;
assign _U1109_in = in[0];
assign _U1109_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1109 (
    .in(_U1109_in),
    .clk(_U1109_clk),
    .out(_U1109_out)
);
assign _U1110_in = in[1];
assign _U1110_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1110 (
    .in(_U1110_in),
    .clk(_U1110_clk),
    .out(_U1110_out)
);
assign _U1111_in = in[2];
assign _U1111_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1111 (
    .in(_U1111_in),
    .clk(_U1111_clk),
    .out(_U1111_out)
);
assign _U1112_in = in[3];
assign _U1112_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1112 (
    .in(_U1112_in),
    .clk(_U1112_clk),
    .out(_U1112_out)
);
assign _U1113_in = in[4];
assign _U1113_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1113 (
    .in(_U1113_in),
    .clk(_U1113_clk),
    .out(_U1113_out)
);
assign out[4] = _U1113_out;
assign out[3] = _U1112_out;
assign out[2] = _U1111_out;
assign out[1] = _U1110_out;
assign out[0] = _U1109_out;
endmodule

module array_delay_U1101 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1102_in;
wire _U1102_clk;
wire [15:0] _U1102_out;
wire [15:0] _U1103_in;
wire _U1103_clk;
wire [15:0] _U1103_out;
wire [15:0] _U1104_in;
wire _U1104_clk;
wire [15:0] _U1104_out;
wire [15:0] _U1105_in;
wire _U1105_clk;
wire [15:0] _U1105_out;
wire [15:0] _U1106_in;
wire _U1106_clk;
wire [15:0] _U1106_out;
assign _U1102_in = in[0];
assign _U1102_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1102 (
    .in(_U1102_in),
    .clk(_U1102_clk),
    .out(_U1102_out)
);
assign _U1103_in = in[1];
assign _U1103_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1103 (
    .in(_U1103_in),
    .clk(_U1103_clk),
    .out(_U1103_out)
);
assign _U1104_in = in[2];
assign _U1104_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1104 (
    .in(_U1104_in),
    .clk(_U1104_clk),
    .out(_U1104_out)
);
assign _U1105_in = in[3];
assign _U1105_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1105 (
    .in(_U1105_in),
    .clk(_U1105_clk),
    .out(_U1105_out)
);
assign _U1106_in = in[4];
assign _U1106_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1106 (
    .in(_U1106_in),
    .clk(_U1106_clk),
    .out(_U1106_out)
);
assign out[4] = _U1106_out;
assign out[3] = _U1105_out;
assign out[2] = _U1104_out;
assign out[1] = _U1103_out;
assign out[0] = _U1102_out;
endmodule

module array_delay_U1094 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1095_in;
wire _U1095_clk;
wire [15:0] _U1095_out;
wire [15:0] _U1096_in;
wire _U1096_clk;
wire [15:0] _U1096_out;
wire [15:0] _U1097_in;
wire _U1097_clk;
wire [15:0] _U1097_out;
wire [15:0] _U1098_in;
wire _U1098_clk;
wire [15:0] _U1098_out;
wire [15:0] _U1099_in;
wire _U1099_clk;
wire [15:0] _U1099_out;
assign _U1095_in = in[0];
assign _U1095_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1095 (
    .in(_U1095_in),
    .clk(_U1095_clk),
    .out(_U1095_out)
);
assign _U1096_in = in[1];
assign _U1096_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1096 (
    .in(_U1096_in),
    .clk(_U1096_clk),
    .out(_U1096_out)
);
assign _U1097_in = in[2];
assign _U1097_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1097 (
    .in(_U1097_in),
    .clk(_U1097_clk),
    .out(_U1097_out)
);
assign _U1098_in = in[3];
assign _U1098_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1098 (
    .in(_U1098_in),
    .clk(_U1098_clk),
    .out(_U1098_out)
);
assign _U1099_in = in[4];
assign _U1099_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1099 (
    .in(_U1099_in),
    .clk(_U1099_clk),
    .out(_U1099_out)
);
assign out[4] = _U1099_out;
assign out[3] = _U1098_out;
assign out[2] = _U1097_out;
assign out[1] = _U1096_out;
assign out[0] = _U1095_out;
endmodule

module array_delay_U1087 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1088_in;
wire _U1088_clk;
wire [15:0] _U1088_out;
wire [15:0] _U1089_in;
wire _U1089_clk;
wire [15:0] _U1089_out;
wire [15:0] _U1090_in;
wire _U1090_clk;
wire [15:0] _U1090_out;
wire [15:0] _U1091_in;
wire _U1091_clk;
wire [15:0] _U1091_out;
wire [15:0] _U1092_in;
wire _U1092_clk;
wire [15:0] _U1092_out;
assign _U1088_in = in[0];
assign _U1088_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1088 (
    .in(_U1088_in),
    .clk(_U1088_clk),
    .out(_U1088_out)
);
assign _U1089_in = in[1];
assign _U1089_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1089 (
    .in(_U1089_in),
    .clk(_U1089_clk),
    .out(_U1089_out)
);
assign _U1090_in = in[2];
assign _U1090_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1090 (
    .in(_U1090_in),
    .clk(_U1090_clk),
    .out(_U1090_out)
);
assign _U1091_in = in[3];
assign _U1091_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1091 (
    .in(_U1091_in),
    .clk(_U1091_clk),
    .out(_U1091_out)
);
assign _U1092_in = in[4];
assign _U1092_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1092 (
    .in(_U1092_in),
    .clk(_U1092_clk),
    .out(_U1092_out)
);
assign out[4] = _U1092_out;
assign out[3] = _U1091_out;
assign out[2] = _U1090_out;
assign out[1] = _U1089_out;
assign out[0] = _U1088_out;
endmodule

module array_delay_U1080 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1081_in;
wire _U1081_clk;
wire [15:0] _U1081_out;
wire [15:0] _U1082_in;
wire _U1082_clk;
wire [15:0] _U1082_out;
wire [15:0] _U1083_in;
wire _U1083_clk;
wire [15:0] _U1083_out;
wire [15:0] _U1084_in;
wire _U1084_clk;
wire [15:0] _U1084_out;
wire [15:0] _U1085_in;
wire _U1085_clk;
wire [15:0] _U1085_out;
assign _U1081_in = in[0];
assign _U1081_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1081 (
    .in(_U1081_in),
    .clk(_U1081_clk),
    .out(_U1081_out)
);
assign _U1082_in = in[1];
assign _U1082_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1082 (
    .in(_U1082_in),
    .clk(_U1082_clk),
    .out(_U1082_out)
);
assign _U1083_in = in[2];
assign _U1083_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1083 (
    .in(_U1083_in),
    .clk(_U1083_clk),
    .out(_U1083_out)
);
assign _U1084_in = in[3];
assign _U1084_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1084 (
    .in(_U1084_in),
    .clk(_U1084_clk),
    .out(_U1084_out)
);
assign _U1085_in = in[4];
assign _U1085_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1085 (
    .in(_U1085_in),
    .clk(_U1085_clk),
    .out(_U1085_out)
);
assign out[4] = _U1085_out;
assign out[3] = _U1084_out;
assign out[2] = _U1083_out;
assign out[1] = _U1082_out;
assign out[0] = _U1081_out;
endmodule

module array_delay_U1073 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1074_in;
wire _U1074_clk;
wire [15:0] _U1074_out;
wire [15:0] _U1075_in;
wire _U1075_clk;
wire [15:0] _U1075_out;
wire [15:0] _U1076_in;
wire _U1076_clk;
wire [15:0] _U1076_out;
wire [15:0] _U1077_in;
wire _U1077_clk;
wire [15:0] _U1077_out;
wire [15:0] _U1078_in;
wire _U1078_clk;
wire [15:0] _U1078_out;
assign _U1074_in = in[0];
assign _U1074_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1074 (
    .in(_U1074_in),
    .clk(_U1074_clk),
    .out(_U1074_out)
);
assign _U1075_in = in[1];
assign _U1075_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1075 (
    .in(_U1075_in),
    .clk(_U1075_clk),
    .out(_U1075_out)
);
assign _U1076_in = in[2];
assign _U1076_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1076 (
    .in(_U1076_in),
    .clk(_U1076_clk),
    .out(_U1076_out)
);
assign _U1077_in = in[3];
assign _U1077_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1077 (
    .in(_U1077_in),
    .clk(_U1077_clk),
    .out(_U1077_out)
);
assign _U1078_in = in[4];
assign _U1078_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1078 (
    .in(_U1078_in),
    .clk(_U1078_clk),
    .out(_U1078_out)
);
assign out[4] = _U1078_out;
assign out[3] = _U1077_out;
assign out[2] = _U1076_out;
assign out[1] = _U1075_out;
assign out[0] = _U1074_out;
endmodule

module array_delay_U1066 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1067_in;
wire _U1067_clk;
wire [15:0] _U1067_out;
wire [15:0] _U1068_in;
wire _U1068_clk;
wire [15:0] _U1068_out;
wire [15:0] _U1069_in;
wire _U1069_clk;
wire [15:0] _U1069_out;
wire [15:0] _U1070_in;
wire _U1070_clk;
wire [15:0] _U1070_out;
wire [15:0] _U1071_in;
wire _U1071_clk;
wire [15:0] _U1071_out;
assign _U1067_in = in[0];
assign _U1067_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1067 (
    .in(_U1067_in),
    .clk(_U1067_clk),
    .out(_U1067_out)
);
assign _U1068_in = in[1];
assign _U1068_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1068 (
    .in(_U1068_in),
    .clk(_U1068_clk),
    .out(_U1068_out)
);
assign _U1069_in = in[2];
assign _U1069_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1069 (
    .in(_U1069_in),
    .clk(_U1069_clk),
    .out(_U1069_out)
);
assign _U1070_in = in[3];
assign _U1070_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1070 (
    .in(_U1070_in),
    .clk(_U1070_clk),
    .out(_U1070_out)
);
assign _U1071_in = in[4];
assign _U1071_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1071 (
    .in(_U1071_in),
    .clk(_U1071_clk),
    .out(_U1071_out)
);
assign out[4] = _U1071_out;
assign out[3] = _U1070_out;
assign out[2] = _U1069_out;
assign out[1] = _U1068_out;
assign out[0] = _U1067_out;
endmodule

module array_delay_U1059 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1060_in;
wire _U1060_clk;
wire [15:0] _U1060_out;
wire [15:0] _U1061_in;
wire _U1061_clk;
wire [15:0] _U1061_out;
wire [15:0] _U1062_in;
wire _U1062_clk;
wire [15:0] _U1062_out;
wire [15:0] _U1063_in;
wire _U1063_clk;
wire [15:0] _U1063_out;
wire [15:0] _U1064_in;
wire _U1064_clk;
wire [15:0] _U1064_out;
assign _U1060_in = in[0];
assign _U1060_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1060 (
    .in(_U1060_in),
    .clk(_U1060_clk),
    .out(_U1060_out)
);
assign _U1061_in = in[1];
assign _U1061_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1061 (
    .in(_U1061_in),
    .clk(_U1061_clk),
    .out(_U1061_out)
);
assign _U1062_in = in[2];
assign _U1062_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1062 (
    .in(_U1062_in),
    .clk(_U1062_clk),
    .out(_U1062_out)
);
assign _U1063_in = in[3];
assign _U1063_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1063 (
    .in(_U1063_in),
    .clk(_U1063_clk),
    .out(_U1063_out)
);
assign _U1064_in = in[4];
assign _U1064_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1064 (
    .in(_U1064_in),
    .clk(_U1064_clk),
    .out(_U1064_out)
);
assign out[4] = _U1064_out;
assign out[3] = _U1063_out;
assign out[2] = _U1062_out;
assign out[1] = _U1061_out;
assign out[0] = _U1060_out;
endmodule

module array_delay_U1052 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1053_in;
wire _U1053_clk;
wire [15:0] _U1053_out;
wire [15:0] _U1054_in;
wire _U1054_clk;
wire [15:0] _U1054_out;
wire [15:0] _U1055_in;
wire _U1055_clk;
wire [15:0] _U1055_out;
wire [15:0] _U1056_in;
wire _U1056_clk;
wire [15:0] _U1056_out;
wire [15:0] _U1057_in;
wire _U1057_clk;
wire [15:0] _U1057_out;
assign _U1053_in = in[0];
assign _U1053_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1053 (
    .in(_U1053_in),
    .clk(_U1053_clk),
    .out(_U1053_out)
);
assign _U1054_in = in[1];
assign _U1054_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1054 (
    .in(_U1054_in),
    .clk(_U1054_clk),
    .out(_U1054_out)
);
assign _U1055_in = in[2];
assign _U1055_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1055 (
    .in(_U1055_in),
    .clk(_U1055_clk),
    .out(_U1055_out)
);
assign _U1056_in = in[3];
assign _U1056_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1056 (
    .in(_U1056_in),
    .clk(_U1056_clk),
    .out(_U1056_out)
);
assign _U1057_in = in[4];
assign _U1057_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1057 (
    .in(_U1057_in),
    .clk(_U1057_clk),
    .out(_U1057_out)
);
assign out[4] = _U1057_out;
assign out[3] = _U1056_out;
assign out[2] = _U1055_out;
assign out[1] = _U1054_out;
assign out[0] = _U1053_out;
endmodule

module array_delay_U1045 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1046_in;
wire _U1046_clk;
wire [15:0] _U1046_out;
wire [15:0] _U1047_in;
wire _U1047_clk;
wire [15:0] _U1047_out;
wire [15:0] _U1048_in;
wire _U1048_clk;
wire [15:0] _U1048_out;
wire [15:0] _U1049_in;
wire _U1049_clk;
wire [15:0] _U1049_out;
wire [15:0] _U1050_in;
wire _U1050_clk;
wire [15:0] _U1050_out;
assign _U1046_in = in[0];
assign _U1046_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1046 (
    .in(_U1046_in),
    .clk(_U1046_clk),
    .out(_U1046_out)
);
assign _U1047_in = in[1];
assign _U1047_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1047 (
    .in(_U1047_in),
    .clk(_U1047_clk),
    .out(_U1047_out)
);
assign _U1048_in = in[2];
assign _U1048_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1048 (
    .in(_U1048_in),
    .clk(_U1048_clk),
    .out(_U1048_out)
);
assign _U1049_in = in[3];
assign _U1049_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1049 (
    .in(_U1049_in),
    .clk(_U1049_clk),
    .out(_U1049_out)
);
assign _U1050_in = in[4];
assign _U1050_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1050 (
    .in(_U1050_in),
    .clk(_U1050_clk),
    .out(_U1050_out)
);
assign out[4] = _U1050_out;
assign out[3] = _U1049_out;
assign out[2] = _U1048_out;
assign out[1] = _U1047_out;
assign out[0] = _U1046_out;
endmodule

module array_delay_U1038 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1039_in;
wire _U1039_clk;
wire [15:0] _U1039_out;
wire [15:0] _U1040_in;
wire _U1040_clk;
wire [15:0] _U1040_out;
wire [15:0] _U1041_in;
wire _U1041_clk;
wire [15:0] _U1041_out;
wire [15:0] _U1042_in;
wire _U1042_clk;
wire [15:0] _U1042_out;
wire [15:0] _U1043_in;
wire _U1043_clk;
wire [15:0] _U1043_out;
assign _U1039_in = in[0];
assign _U1039_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1039 (
    .in(_U1039_in),
    .clk(_U1039_clk),
    .out(_U1039_out)
);
assign _U1040_in = in[1];
assign _U1040_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1040 (
    .in(_U1040_in),
    .clk(_U1040_clk),
    .out(_U1040_out)
);
assign _U1041_in = in[2];
assign _U1041_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1041 (
    .in(_U1041_in),
    .clk(_U1041_clk),
    .out(_U1041_out)
);
assign _U1042_in = in[3];
assign _U1042_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1042 (
    .in(_U1042_in),
    .clk(_U1042_clk),
    .out(_U1042_out)
);
assign _U1043_in = in[4];
assign _U1043_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1043 (
    .in(_U1043_in),
    .clk(_U1043_clk),
    .out(_U1043_out)
);
assign out[4] = _U1043_out;
assign out[3] = _U1042_out;
assign out[2] = _U1041_out;
assign out[1] = _U1040_out;
assign out[0] = _U1039_out;
endmodule

module array_delay_U1012 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1013_in;
wire _U1013_clk;
wire [15:0] _U1013_out;
wire [15:0] _U1014_in;
wire _U1014_clk;
wire [15:0] _U1014_out;
wire [15:0] _U1015_in;
wire _U1015_clk;
wire [15:0] _U1015_out;
wire [15:0] _U1016_in;
wire _U1016_clk;
wire [15:0] _U1016_out;
wire [15:0] _U1017_in;
wire _U1017_clk;
wire [15:0] _U1017_out;
assign _U1013_in = in[0];
assign _U1013_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1013 (
    .in(_U1013_in),
    .clk(_U1013_clk),
    .out(_U1013_out)
);
assign _U1014_in = in[1];
assign _U1014_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1014 (
    .in(_U1014_in),
    .clk(_U1014_clk),
    .out(_U1014_out)
);
assign _U1015_in = in[2];
assign _U1015_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1015 (
    .in(_U1015_in),
    .clk(_U1015_clk),
    .out(_U1015_out)
);
assign _U1016_in = in[3];
assign _U1016_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1016 (
    .in(_U1016_in),
    .clk(_U1016_clk),
    .out(_U1016_out)
);
assign _U1017_in = in[4];
assign _U1017_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1017 (
    .in(_U1017_in),
    .clk(_U1017_clk),
    .out(_U1017_out)
);
assign out[4] = _U1017_out;
assign out[3] = _U1016_out;
assign out[2] = _U1015_out;
assign out[1] = _U1014_out;
assign out[0] = _U1013_out;
endmodule

module array_delay_U1005 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U1006_in;
wire _U1006_clk;
wire [15:0] _U1006_out;
wire [15:0] _U1007_in;
wire _U1007_clk;
wire [15:0] _U1007_out;
wire [15:0] _U1008_in;
wire _U1008_clk;
wire [15:0] _U1008_out;
wire [15:0] _U1009_in;
wire _U1009_clk;
wire [15:0] _U1009_out;
wire [15:0] _U1010_in;
wire _U1010_clk;
wire [15:0] _U1010_out;
assign _U1006_in = in[0];
assign _U1006_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1006 (
    .in(_U1006_in),
    .clk(_U1006_clk),
    .out(_U1006_out)
);
assign _U1007_in = in[1];
assign _U1007_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1007 (
    .in(_U1007_in),
    .clk(_U1007_clk),
    .out(_U1007_out)
);
assign _U1008_in = in[2];
assign _U1008_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1008 (
    .in(_U1008_in),
    .clk(_U1008_clk),
    .out(_U1008_out)
);
assign _U1009_in = in[3];
assign _U1009_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1009 (
    .in(_U1009_in),
    .clk(_U1009_clk),
    .out(_U1009_out)
);
assign _U1010_in = in[4];
assign _U1010_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1010 (
    .in(_U1010_in),
    .clk(_U1010_clk),
    .out(_U1010_out)
);
assign out[4] = _U1010_out;
assign out[3] = _U1009_out;
assign out[2] = _U1008_out;
assign out[1] = _U1007_out;
assign out[0] = _U1006_out;
endmodule

module aff__U969 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U968 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U969 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U93 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U92 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U93 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U781 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U780 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U781 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U70 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U69 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U70 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U593 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U592 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U593 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U47 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U46 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U47 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U405 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U404 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U405 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U382 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U381 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U382 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U359 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U358 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U359 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U336 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U335 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U336 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U313 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U312 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U313 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U290 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U289 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U290 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U267 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U266 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U267 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U244 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U243 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U244 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U24 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U23 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U24 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U2238 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U2237 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U2238 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U221 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U220 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U221 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U2191 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U2190 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U2191 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U2144 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U2143 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U2144 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U2097 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U2096 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U2097 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U2050 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U2049 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U2050 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U2003 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U2002 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U2003 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1956 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U1955 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1956 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1909 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h3e91);
endmodule

module affine_controller__U1908 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1909 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U185 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h00d8 * d[1])))) + (16'(16'h0048 * d[2])))) + (16'(16'h0009 * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h0002);
endmodule

module affine_controller__U184 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U185 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h0007;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h0007;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1721 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U1720 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1721 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U162 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U161 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U162 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1533 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U1532 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1533 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U139 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U138 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U139 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1345 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U1344 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1345 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U116 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U115 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U116 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1157 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h03ea);
endmodule

module affine_controller__U1156 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1157 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001f * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0001);
endmodule

module affine_controller__U0 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module _U996_pt__U997 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U990_pt__U991 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U981_pt__U982 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U978_pt__U979 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U969_pt__U970 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U966_pt__U967 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U963_pt__U964 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U95_pt__U96 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U951_pt__U952 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U946_pt__U947 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U941_pt__U942 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U934_pt__U935 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U927_pt__U928 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U924_pt__U925 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U918_pt__U919 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U912_pt__U913 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U910_pt__U911 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U908_pt__U909 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U904_pt__U905 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U901_pt__U902 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U8_pt__U9 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_4_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
wire [15:0] _U8_in;
assign _U8_in = in0_hw_input_stencil[0];
_U8_pt__U9 _U8 (
    .in(_U8_in),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil_4 (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read[0];
hcompute_hw_input_global_wrapper_stencil_4_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U898_pt__U899 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U888_pt__U889 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U881_pt__U882 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U87_pt__U88 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U873_pt__U874 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U870_pt__U871 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U854_pt__U855 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U838_pt__U839 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U835_pt__U836 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U818_pt__U819 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U810_pt__U811 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U80_pt__U81 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U807_pt__U808 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U797_pt__U798 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U795_pt__U796 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U792_pt__U793 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U783_pt__U784 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U780_pt__U781 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U776_pt__U777 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U760_pt__U761 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U757_pt__U758 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U752_pt__U753 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U749_pt__U750 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U73_pt__U74 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U735_pt__U736 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U732_pt__U733 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U730_pt__U731 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U726_pt__U727 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U719_pt__U720 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U711_pt__U712 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U704_pt__U705 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U6_pt__U7 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_3_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
wire [15:0] _U6_in;
assign _U6_in = in0_hw_input_stencil[0];
_U6_pt__U7 _U6 (
    .in(_U6_in),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil_3 (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read[0];
hcompute_hw_input_global_wrapper_stencil_3_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U698_pt__U699 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U692_pt__U693 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U684_pt__U685 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U67_pt__U68 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U672_pt__U673 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U663_pt__U664 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U661_pt__U662 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U658_pt__U659 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U653_pt__U654 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U647_pt__U648 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U644_pt__U645 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U640_pt__U641 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U637_pt__U638 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_11_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U637_in;
wire [15:0] _U637_out;
wire [15:0] _U639_in;
wire _U639_clk;
wire [15:0] _U639_out;
wire [15:0] _U640_in;
wire [15:0] _U640_out;
wire [15:0] _U642_in;
wire _U642_clk;
wire [15:0] _U642_out;
wire [15:0] _U643_in;
wire _U643_clk;
wire [15:0] _U643_out;
wire [15:0] _U644_in;
wire [15:0] _U644_out;
wire [15:0] _U646_in;
wire _U646_clk;
wire [15:0] _U646_out;
wire [15:0] _U647_in;
wire [15:0] _U647_out;
wire [15:0] _U649_in;
wire _U649_clk;
wire [15:0] _U649_out;
wire [15:0] _U650_in;
wire _U650_clk;
wire [15:0] _U650_out;
wire [15:0] _U651_in;
wire _U651_clk;
wire [15:0] _U651_out;
wire [15:0] _U652_in;
wire _U652_clk;
wire [15:0] _U652_out;
wire [15:0] _U653_in;
wire [15:0] _U653_out;
wire [15:0] _U655_in;
wire _U655_clk;
wire [15:0] _U655_out;
wire [15:0] _U656_in;
wire _U656_clk;
wire [15:0] _U656_out;
wire [15:0] _U657_in;
wire _U657_clk;
wire [15:0] _U657_out;
wire [15:0] _U658_in;
wire [15:0] _U658_out;
wire [15:0] _U660_in;
wire _U660_clk;
wire [15:0] _U660_out;
wire [15:0] _U661_in;
wire [15:0] _U661_out;
wire [15:0] _U663_in;
wire [15:0] _U663_out;
wire [15:0] _U665_in;
wire _U665_clk;
wire [15:0] _U665_out;
wire [15:0] _U666_in;
wire _U666_clk;
wire [15:0] _U666_out;
wire [15:0] _U667_in;
wire _U667_clk;
wire [15:0] _U667_out;
wire [15:0] _U668_in;
wire _U668_clk;
wire [15:0] _U668_out;
wire [15:0] _U669_in;
wire _U669_clk;
wire [15:0] _U669_out;
wire [15:0] _U670_in;
wire _U670_clk;
wire [15:0] _U670_out;
wire [15:0] _U671_in;
wire _U671_clk;
wire [15:0] _U671_out;
wire [15:0] _U672_in;
wire [15:0] _U672_out;
wire [15:0] _U674_in;
wire _U674_clk;
wire [15:0] _U674_out;
wire [15:0] _U675_in;
wire _U675_clk;
wire [15:0] _U675_out;
wire [15:0] _U676_in;
wire _U676_clk;
wire [15:0] _U676_out;
wire [15:0] _U677_in;
wire _U677_clk;
wire [15:0] _U677_out;
wire [15:0] _U678_in;
wire _U678_clk;
wire [15:0] _U678_out;
wire [15:0] _U679_in;
wire _U679_clk;
wire [15:0] _U679_out;
wire [15:0] _U680_in;
wire _U680_clk;
wire [15:0] _U680_out;
wire [15:0] _U681_in;
wire _U681_clk;
wire [15:0] _U681_out;
wire [15:0] _U682_in;
wire _U682_clk;
wire [15:0] _U682_out;
wire [15:0] _U683_in;
wire _U683_clk;
wire [15:0] _U683_out;
wire [15:0] _U684_in;
wire [15:0] _U684_out;
wire [15:0] _U686_in;
wire _U686_clk;
wire [15:0] _U686_out;
wire [15:0] _U687_in;
wire _U687_clk;
wire [15:0] _U687_out;
wire [15:0] _U688_in;
wire _U688_clk;
wire [15:0] _U688_out;
wire [15:0] _U689_in;
wire _U689_clk;
wire [15:0] _U689_out;
wire [15:0] _U690_in;
wire _U690_clk;
wire [15:0] _U690_out;
wire [15:0] _U691_in;
wire _U691_clk;
wire [15:0] _U691_out;
wire [15:0] _U692_in;
wire [15:0] _U692_out;
wire [15:0] _U694_in;
wire _U694_clk;
wire [15:0] _U694_out;
wire [15:0] _U695_in;
wire _U695_clk;
wire [15:0] _U695_out;
wire [15:0] _U696_in;
wire _U696_clk;
wire [15:0] _U696_out;
wire [15:0] _U697_in;
wire _U697_clk;
wire [15:0] _U697_out;
wire [15:0] _U698_in;
wire [15:0] _U698_out;
wire [15:0] _U700_in;
wire _U700_clk;
wire [15:0] _U700_out;
wire [15:0] _U701_in;
wire _U701_clk;
wire [15:0] _U701_out;
wire [15:0] _U702_in;
wire _U702_clk;
wire [15:0] _U702_out;
wire [15:0] _U703_in;
wire _U703_clk;
wire [15:0] _U703_out;
wire [15:0] _U704_in;
wire [15:0] _U704_out;
wire [15:0] _U706_in;
wire _U706_clk;
wire [15:0] _U706_out;
wire [15:0] _U707_in;
wire _U707_clk;
wire [15:0] _U707_out;
wire [15:0] _U708_in;
wire _U708_clk;
wire [15:0] _U708_out;
wire [15:0] _U709_in;
wire _U709_clk;
wire [15:0] _U709_out;
wire [15:0] _U710_in;
wire _U710_clk;
wire [15:0] _U710_out;
wire [15:0] _U711_in;
wire [15:0] _U711_out;
wire [15:0] _U713_in;
wire _U713_clk;
wire [15:0] _U713_out;
wire [15:0] _U714_in;
wire _U714_clk;
wire [15:0] _U714_out;
wire [15:0] _U715_in;
wire _U715_clk;
wire [15:0] _U715_out;
wire [15:0] _U716_in;
wire _U716_clk;
wire [15:0] _U716_out;
wire [15:0] _U717_in;
wire _U717_clk;
wire [15:0] _U717_out;
wire [15:0] _U718_in;
wire _U718_clk;
wire [15:0] _U718_out;
wire [15:0] _U719_in;
wire [15:0] _U719_out;
wire [15:0] _U721_in;
wire _U721_clk;
wire [15:0] _U721_out;
wire [15:0] _U722_in;
wire _U722_clk;
wire [15:0] _U722_out;
wire [15:0] _U723_in;
wire _U723_clk;
wire [15:0] _U723_out;
wire [15:0] _U724_in;
wire _U724_clk;
wire [15:0] _U724_out;
wire [15:0] _U725_in;
wire _U725_clk;
wire [15:0] _U725_out;
wire [15:0] _U726_in;
wire [15:0] _U726_out;
wire [15:0] _U728_in;
wire _U728_clk;
wire [15:0] _U728_out;
wire [15:0] _U729_in;
wire _U729_clk;
wire [15:0] _U729_out;
wire [15:0] _U730_in;
wire [15:0] _U730_out;
wire [15:0] _U732_in;
wire [15:0] _U732_out;
wire [15:0] _U734_in;
wire _U734_clk;
wire [15:0] _U734_out;
wire [15:0] _U735_in;
wire [15:0] _U735_out;
wire [15:0] _U737_in;
wire _U737_clk;
wire [15:0] _U737_out;
wire [15:0] _U738_in;
wire _U738_clk;
wire [15:0] _U738_out;
wire [15:0] _U739_in;
wire _U739_clk;
wire [15:0] _U739_out;
wire [15:0] _U740_in;
wire _U740_clk;
wire [15:0] _U740_out;
wire [15:0] _U741_in;
wire _U741_clk;
wire [15:0] _U741_out;
wire [15:0] _U742_in;
wire _U742_clk;
wire [15:0] _U742_out;
wire [15:0] _U743_in;
wire _U743_clk;
wire [15:0] _U743_out;
wire [15:0] _U744_in;
wire _U744_clk;
wire [15:0] _U744_out;
wire [15:0] _U745_in;
wire _U745_clk;
wire [15:0] _U745_out;
wire [15:0] _U746_in;
wire _U746_clk;
wire [15:0] _U746_out;
wire [15:0] _U747_in;
wire _U747_clk;
wire [15:0] _U747_out;
wire [15:0] _U748_in;
wire _U748_clk;
wire [15:0] _U748_out;
wire [15:0] _U749_in;
wire [15:0] _U749_out;
wire [15:0] _U751_in;
wire _U751_clk;
wire [15:0] _U751_out;
wire [15:0] _U752_in;
wire [15:0] _U752_out;
wire [15:0] _U754_in;
wire _U754_clk;
wire [15:0] _U754_out;
wire [15:0] _U755_in;
wire _U755_clk;
wire [15:0] _U755_out;
wire [15:0] _U756_in;
wire _U756_clk;
wire [15:0] _U756_out;
wire [15:0] _U757_in;
wire [15:0] _U757_out;
wire [15:0] _U759_in;
wire _U759_clk;
wire [15:0] _U759_out;
wire [15:0] _U760_in;
wire [15:0] _U760_out;
wire [15:0] _U762_in;
wire _U762_clk;
wire [15:0] _U762_out;
wire [15:0] _U763_in;
wire _U763_clk;
wire [15:0] _U763_out;
wire [15:0] _U764_in;
wire _U764_clk;
wire [15:0] _U764_out;
wire [15:0] _U765_in;
wire _U765_clk;
wire [15:0] _U765_out;
wire [15:0] _U766_in;
wire _U766_clk;
wire [15:0] _U766_out;
wire [15:0] _U767_in;
wire _U767_clk;
wire [15:0] _U767_out;
wire [15:0] _U768_in;
wire _U768_clk;
wire [15:0] _U768_out;
wire [15:0] _U769_in;
wire _U769_clk;
wire [15:0] _U769_out;
wire [15:0] _U770_in;
wire _U770_clk;
wire [15:0] _U770_out;
wire [15:0] _U771_in;
wire _U771_clk;
wire [15:0] _U771_out;
wire [15:0] _U772_in;
wire _U772_clk;
wire [15:0] _U772_out;
wire [15:0] _U773_in;
wire _U773_clk;
wire [15:0] _U773_out;
wire [15:0] _U774_in;
wire _U774_clk;
wire [15:0] _U774_out;
wire [15:0] _U775_in;
wire _U775_clk;
wire [15:0] _U775_out;
wire [15:0] _U776_in;
wire [15:0] _U776_out;
wire [15:0] _U778_in;
wire _U778_clk;
wire [15:0] _U778_out;
wire [15:0] _U779_in;
wire _U779_clk;
wire [15:0] _U779_out;
wire [15:0] _U780_in;
wire [15:0] _U780_out;
wire [15:0] _U782_in;
wire _U782_clk;
wire [15:0] _U782_out;
wire [15:0] _U783_in;
wire [15:0] _U783_out;
wire [15:0] _U785_in;
wire _U785_clk;
wire [15:0] _U785_out;
wire [15:0] _U786_in;
wire _U786_clk;
wire [15:0] _U786_out;
wire [15:0] _U787_in;
wire _U787_clk;
wire [15:0] _U787_out;
wire [15:0] _U788_in;
wire _U788_clk;
wire [15:0] _U788_out;
wire [15:0] _U789_in;
wire _U789_clk;
wire [15:0] _U789_out;
wire [15:0] _U790_in;
wire _U790_clk;
wire [15:0] _U790_out;
wire [15:0] _U791_in;
wire _U791_clk;
wire [15:0] _U791_out;
wire [15:0] _U792_in;
wire [15:0] _U792_out;
wire [15:0] _U794_in;
wire _U794_clk;
wire [15:0] _U794_out;
wire [15:0] _U795_in;
wire [15:0] _U797_in;
wire [15:0] _U797_out;
wire [15:0] _U799_in;
wire _U799_clk;
wire [15:0] _U799_out;
wire [15:0] _U800_in;
wire _U800_clk;
wire [15:0] _U800_out;
wire [15:0] _U801_in;
wire _U801_clk;
wire [15:0] _U801_out;
wire [15:0] _U802_in;
wire _U802_clk;
wire [15:0] _U802_out;
wire [15:0] _U803_in;
wire _U803_clk;
wire [15:0] _U803_out;
wire [15:0] _U804_in;
wire _U804_clk;
wire [15:0] _U804_out;
wire [15:0] _U805_in;
wire _U805_clk;
wire [15:0] _U805_out;
wire [15:0] _U806_in;
wire _U806_clk;
wire [15:0] _U806_out;
wire [15:0] _U807_in;
wire [15:0] _U807_out;
wire [15:0] _U809_in;
wire _U809_clk;
wire [15:0] _U809_out;
wire [15:0] _U810_in;
wire [15:0] _U810_out;
wire [15:0] _U812_in;
wire _U812_clk;
wire [15:0] _U812_out;
wire [15:0] _U813_in;
wire _U813_clk;
wire [15:0] _U813_out;
wire [15:0] _U814_in;
wire _U814_clk;
wire [15:0] _U814_out;
wire [15:0] _U815_in;
wire _U815_clk;
wire [15:0] _U815_out;
wire [15:0] _U816_in;
wire _U816_clk;
wire [15:0] _U816_out;
wire [15:0] _U817_in;
wire _U817_clk;
wire [15:0] _U817_out;
wire [15:0] _U818_in;
wire [15:0] _U818_out;
wire [15:0] _U820_in;
wire _U820_clk;
wire [15:0] _U820_out;
wire [15:0] _U821_in;
wire _U821_clk;
wire [15:0] _U821_out;
wire [15:0] _U822_in;
wire _U822_clk;
wire [15:0] _U822_out;
wire [15:0] _U823_in;
wire _U823_clk;
wire [15:0] _U823_out;
wire [15:0] _U824_in;
wire _U824_clk;
wire [15:0] _U824_out;
wire [15:0] _U825_in;
wire _U825_clk;
wire [15:0] _U825_out;
wire [15:0] _U826_in;
wire _U826_clk;
wire [15:0] _U826_out;
wire [15:0] _U827_in;
wire _U827_clk;
wire [15:0] _U827_out;
wire [15:0] _U828_in;
wire _U828_clk;
wire [15:0] _U828_out;
wire [15:0] _U829_in;
wire _U829_clk;
wire [15:0] _U829_out;
wire [15:0] _U830_in;
wire _U830_clk;
wire [15:0] _U830_out;
wire [15:0] _U831_in;
wire _U831_clk;
wire [15:0] _U831_out;
wire [15:0] _U832_in;
wire _U832_clk;
wire [15:0] _U832_out;
wire [15:0] _U833_in;
wire _U833_clk;
wire [15:0] _U833_out;
wire [15:0] _U834_in;
wire _U834_clk;
wire [15:0] _U834_out;
wire [15:0] _U835_in;
wire [15:0] _U835_out;
wire [15:0] _U837_in;
wire _U837_clk;
wire [15:0] _U837_out;
assign _U637_in = _U639_out;
_U637_pt__U638 _U637 (
    .in(_U637_in),
    .out(_U637_out)
);
assign _U639_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U639_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U639 (
    .in(_U639_in),
    .clk(_U639_clk),
    .out(_U639_out)
);
assign _U640_in = _U643_out;
_U640_pt__U641 _U640 (
    .in(_U640_in),
    .out(_U640_out)
);
assign _U642_in = in1_hw_input_global_wrapper_stencil[2];
assign _U642_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U642 (
    .in(_U642_in),
    .clk(_U642_clk),
    .out(_U642_out)
);
assign _U643_in = _U642_out;
assign _U643_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U643 (
    .in(_U643_in),
    .clk(_U643_clk),
    .out(_U643_out)
);
assign _U644_in = _U646_out;
_U644_pt__U645 _U644 (
    .in(_U644_in),
    .out(_U644_out)
);
assign _U646_in = 16'(_U698_out + _U749_out);
assign _U646_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U646 (
    .in(_U646_in),
    .clk(_U646_clk),
    .out(_U646_out)
);
assign _U647_in = _U652_out;
_U647_pt__U648 _U647 (
    .in(_U647_in),
    .out(_U647_out)
);
assign _U649_in = in1_hw_input_global_wrapper_stencil[4];
assign _U649_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U649 (
    .in(_U649_in),
    .clk(_U649_clk),
    .out(_U649_out)
);
assign _U650_in = _U649_out;
assign _U650_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U650 (
    .in(_U650_in),
    .clk(_U650_clk),
    .out(_U650_out)
);
assign _U651_in = _U650_out;
assign _U651_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U651 (
    .in(_U651_in),
    .clk(_U651_clk),
    .out(_U651_out)
);
assign _U652_in = _U651_out;
assign _U652_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U652 (
    .in(_U652_in),
    .clk(_U652_clk),
    .out(_U652_out)
);
assign _U653_in = _U657_out;
_U653_pt__U654 _U653 (
    .in(_U653_in),
    .out(_U653_out)
);
assign _U655_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U655_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U655 (
    .in(_U655_in),
    .clk(_U655_clk),
    .out(_U655_out)
);
assign _U656_in = _U655_out;
assign _U656_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U656 (
    .in(_U656_in),
    .clk(_U656_clk),
    .out(_U656_out)
);
assign _U657_in = _U656_out;
assign _U657_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U657 (
    .in(_U657_in),
    .clk(_U657_clk),
    .out(_U657_out)
);
assign _U658_in = _U660_out;
_U658_pt__U659 _U658 (
    .in(_U658_in),
    .out(_U658_out)
);
assign _U660_in = in1_hw_input_global_wrapper_stencil[1];
assign _U660_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U660 (
    .in(_U660_in),
    .clk(_U660_clk),
    .out(_U660_out)
);
assign _U661_in = in2_hw_kernel_global_wrapper_stencil[0];
_U661_pt__U662 _U661 (
    .in(_U661_in),
    .out(_U661_out)
);
assign _U663_in = _U671_out;
_U663_pt__U664 _U663 (
    .in(_U663_in),
    .out(_U663_out)
);
assign _U665_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U665_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U665 (
    .in(_U665_in),
    .clk(_U665_clk),
    .out(_U665_out)
);
assign _U666_in = _U665_out;
assign _U666_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U666 (
    .in(_U666_in),
    .clk(_U666_clk),
    .out(_U666_out)
);
assign _U667_in = _U666_out;
assign _U667_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U667 (
    .in(_U667_in),
    .clk(_U667_clk),
    .out(_U667_out)
);
assign _U668_in = _U667_out;
assign _U668_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U668 (
    .in(_U668_in),
    .clk(_U668_clk),
    .out(_U668_out)
);
assign _U669_in = _U668_out;
assign _U669_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U669 (
    .in(_U669_in),
    .clk(_U669_clk),
    .out(_U669_out)
);
assign _U670_in = _U669_out;
assign _U670_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U670 (
    .in(_U670_in),
    .clk(_U670_clk),
    .out(_U670_out)
);
assign _U671_in = _U670_out;
assign _U671_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U671 (
    .in(_U671_in),
    .clk(_U671_clk),
    .out(_U671_out)
);
assign _U672_in = _U683_out;
_U672_pt__U673 _U672 (
    .in(_U672_in),
    .out(_U672_out)
);
assign _U674_in = 16'(_U726_out * _U640_out);
assign _U674_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U674 (
    .in(_U674_in),
    .clk(_U674_clk),
    .out(_U674_out)
);
assign _U675_in = _U674_out;
assign _U675_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U675 (
    .in(_U675_in),
    .clk(_U675_clk),
    .out(_U675_out)
);
assign _U676_in = _U675_out;
assign _U676_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U676 (
    .in(_U676_in),
    .clk(_U676_clk),
    .out(_U676_out)
);
assign _U677_in = _U676_out;
assign _U677_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U677 (
    .in(_U677_in),
    .clk(_U677_clk),
    .out(_U677_out)
);
assign _U678_in = _U677_out;
assign _U678_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U678 (
    .in(_U678_in),
    .clk(_U678_clk),
    .out(_U678_out)
);
assign _U679_in = _U678_out;
assign _U679_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U679 (
    .in(_U679_in),
    .clk(_U679_clk),
    .out(_U679_out)
);
assign _U680_in = _U679_out;
assign _U680_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U680 (
    .in(_U680_in),
    .clk(_U680_clk),
    .out(_U680_out)
);
assign _U681_in = _U680_out;
assign _U681_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U681 (
    .in(_U681_in),
    .clk(_U681_clk),
    .out(_U681_out)
);
assign _U682_in = _U681_out;
assign _U682_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U682 (
    .in(_U682_in),
    .clk(_U682_clk),
    .out(_U682_out)
);
assign _U683_in = _U682_out;
assign _U683_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U683 (
    .in(_U683_in),
    .clk(_U683_clk),
    .out(_U683_out)
);
assign _U684_in = _U691_out;
_U684_pt__U685 _U684 (
    .in(_U684_in),
    .out(_U684_out)
);
assign _U686_in = in1_hw_input_global_wrapper_stencil[6];
assign _U686_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U686 (
    .in(_U686_in),
    .clk(_U686_clk),
    .out(_U686_out)
);
assign _U687_in = _U686_out;
assign _U687_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U687 (
    .in(_U687_in),
    .clk(_U687_clk),
    .out(_U687_out)
);
assign _U688_in = _U687_out;
assign _U688_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U688 (
    .in(_U688_in),
    .clk(_U688_clk),
    .out(_U688_out)
);
assign _U689_in = _U688_out;
assign _U689_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U689 (
    .in(_U689_in),
    .clk(_U689_clk),
    .out(_U689_out)
);
assign _U690_in = _U689_out;
assign _U690_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U690 (
    .in(_U690_in),
    .clk(_U690_clk),
    .out(_U690_out)
);
assign _U691_in = _U690_out;
assign _U691_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U691 (
    .in(_U691_in),
    .clk(_U691_clk),
    .out(_U691_out)
);
assign _U692_in = _U697_out;
_U692_pt__U693 _U692 (
    .in(_U692_in),
    .out(_U692_out)
);
assign _U694_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U694_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U694 (
    .in(_U694_in),
    .clk(_U694_clk),
    .out(_U694_out)
);
assign _U695_in = _U694_out;
assign _U695_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U695 (
    .in(_U695_in),
    .clk(_U695_clk),
    .out(_U695_out)
);
assign _U696_in = _U695_out;
assign _U696_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U696 (
    .in(_U696_in),
    .clk(_U696_clk),
    .out(_U696_out)
);
assign _U697_in = _U696_out;
assign _U697_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U697 (
    .in(_U697_in),
    .clk(_U697_clk),
    .out(_U697_out)
);
assign _U698_in = _U703_out;
_U698_pt__U699 _U698 (
    .in(_U698_in),
    .out(_U698_out)
);
assign _U700_in = 16'(_U704_out * _U719_out);
assign _U700_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U700 (
    .in(_U700_in),
    .clk(_U700_clk),
    .out(_U700_out)
);
assign _U701_in = _U700_out;
assign _U701_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U701 (
    .in(_U701_in),
    .clk(_U701_clk),
    .out(_U701_out)
);
assign _U702_in = _U701_out;
assign _U702_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U702 (
    .in(_U702_in),
    .clk(_U702_clk),
    .out(_U702_out)
);
assign _U703_in = _U702_out;
assign _U703_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U703 (
    .in(_U703_in),
    .clk(_U703_clk),
    .out(_U703_out)
);
assign _U704_in = _U710_out;
_U704_pt__U705 _U704 (
    .in(_U704_in),
    .out(_U704_out)
);
assign _U706_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U706_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U706 (
    .in(_U706_in),
    .clk(_U706_clk),
    .out(_U706_out)
);
assign _U707_in = _U706_out;
assign _U707_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U707 (
    .in(_U707_in),
    .clk(_U707_clk),
    .out(_U707_out)
);
assign _U708_in = _U707_out;
assign _U708_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U708 (
    .in(_U708_in),
    .clk(_U708_clk),
    .out(_U708_out)
);
assign _U709_in = _U708_out;
assign _U709_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U709 (
    .in(_U709_in),
    .clk(_U709_clk),
    .out(_U709_out)
);
assign _U710_in = _U709_out;
assign _U710_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U710 (
    .in(_U710_in),
    .clk(_U710_clk),
    .out(_U710_out)
);
assign _U711_in = _U718_out;
_U711_pt__U712 _U711 (
    .in(_U711_in),
    .out(_U711_out)
);
assign _U713_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U713_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U713 (
    .in(_U713_in),
    .clk(_U713_clk),
    .out(_U713_out)
);
assign _U714_in = _U713_out;
assign _U714_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U714 (
    .in(_U714_in),
    .clk(_U714_clk),
    .out(_U714_out)
);
assign _U715_in = _U714_out;
assign _U715_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U715 (
    .in(_U715_in),
    .clk(_U715_clk),
    .out(_U715_out)
);
assign _U716_in = _U715_out;
assign _U716_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U716 (
    .in(_U716_in),
    .clk(_U716_clk),
    .out(_U716_out)
);
assign _U717_in = _U716_out;
assign _U717_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U717 (
    .in(_U717_in),
    .clk(_U717_clk),
    .out(_U717_out)
);
assign _U718_in = _U717_out;
assign _U718_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U718 (
    .in(_U718_in),
    .clk(_U718_clk),
    .out(_U718_out)
);
assign _U719_in = _U725_out;
_U719_pt__U720 _U719 (
    .in(_U719_in),
    .out(_U719_out)
);
assign _U721_in = in1_hw_input_global_wrapper_stencil[5];
assign _U721_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U721 (
    .in(_U721_in),
    .clk(_U721_clk),
    .out(_U721_out)
);
assign _U722_in = _U721_out;
assign _U722_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U722 (
    .in(_U722_in),
    .clk(_U722_clk),
    .out(_U722_out)
);
assign _U723_in = _U722_out;
assign _U723_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U723 (
    .in(_U723_in),
    .clk(_U723_clk),
    .out(_U723_out)
);
assign _U724_in = _U723_out;
assign _U724_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U724 (
    .in(_U724_in),
    .clk(_U724_clk),
    .out(_U724_out)
);
assign _U725_in = _U724_out;
assign _U725_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U725 (
    .in(_U725_in),
    .clk(_U725_clk),
    .out(_U725_out)
);
assign _U726_in = _U729_out;
_U726_pt__U727 _U726 (
    .in(_U726_in),
    .out(_U726_out)
);
assign _U728_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U728_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U728 (
    .in(_U728_in),
    .clk(_U728_clk),
    .out(_U728_out)
);
assign _U729_in = _U728_out;
assign _U729_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U729 (
    .in(_U729_in),
    .clk(_U729_clk),
    .out(_U729_out)
);
assign _U730_in = in1_hw_input_global_wrapper_stencil[0];
_U730_pt__U731 _U730 (
    .in(_U730_in),
    .out(_U730_out)
);
assign _U732_in = _U734_out;
_U732_pt__U733 _U732 (
    .in(_U732_in),
    .out(_U732_out)
);
assign _U734_in = 16'(_U797_out + _U792_out);
assign _U734_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U734 (
    .in(_U734_in),
    .clk(_U734_clk),
    .out(_U734_out)
);
assign _U735_in = _U748_out;
_U735_pt__U736 _U735 (
    .in(_U735_in),
    .out(_U735_out)
);
assign _U737_in = 16'(_U637_out * _U658_out);
assign _U737_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U737 (
    .in(_U737_in),
    .clk(_U737_clk),
    .out(_U737_out)
);
assign _U738_in = _U737_out;
assign _U738_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U738 (
    .in(_U738_in),
    .clk(_U738_clk),
    .out(_U738_out)
);
assign _U739_in = _U738_out;
assign _U739_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U739 (
    .in(_U739_in),
    .clk(_U739_clk),
    .out(_U739_out)
);
assign _U740_in = _U739_out;
assign _U740_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U740 (
    .in(_U740_in),
    .clk(_U740_clk),
    .out(_U740_out)
);
assign _U741_in = _U740_out;
assign _U741_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U741 (
    .in(_U741_in),
    .clk(_U741_clk),
    .out(_U741_out)
);
assign _U742_in = _U741_out;
assign _U742_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U742 (
    .in(_U742_in),
    .clk(_U742_clk),
    .out(_U742_out)
);
assign _U743_in = _U742_out;
assign _U743_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U743 (
    .in(_U743_in),
    .clk(_U743_clk),
    .out(_U743_out)
);
assign _U744_in = _U743_out;
assign _U744_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U744 (
    .in(_U744_in),
    .clk(_U744_clk),
    .out(_U744_out)
);
assign _U745_in = _U744_out;
assign _U745_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U745 (
    .in(_U745_in),
    .clk(_U745_clk),
    .out(_U745_out)
);
assign _U746_in = _U745_out;
assign _U746_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U746 (
    .in(_U746_in),
    .clk(_U746_clk),
    .out(_U746_out)
);
assign _U747_in = _U746_out;
assign _U747_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U747 (
    .in(_U747_in),
    .clk(_U747_clk),
    .out(_U747_out)
);
assign _U748_in = _U747_out;
assign _U748_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U748 (
    .in(_U748_in),
    .clk(_U748_clk),
    .out(_U748_out)
);
assign _U749_in = _U751_out;
_U749_pt__U750 _U749 (
    .in(_U749_in),
    .out(_U749_out)
);
assign _U751_in = 16'(_U776_out + _U757_out);
assign _U751_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U751 (
    .in(_U751_in),
    .clk(_U751_clk),
    .out(_U751_out)
);
assign _U752_in = _U756_out;
_U752_pt__U753 _U752 (
    .in(_U752_in),
    .out(_U752_out)
);
assign _U754_in = in1_hw_input_global_wrapper_stencil[3];
assign _U754_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U754 (
    .in(_U754_in),
    .clk(_U754_clk),
    .out(_U754_out)
);
assign _U755_in = _U754_out;
assign _U755_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U755 (
    .in(_U755_in),
    .clk(_U755_clk),
    .out(_U755_out)
);
assign _U756_in = _U755_out;
assign _U756_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U756 (
    .in(_U756_in),
    .clk(_U756_clk),
    .out(_U756_out)
);
assign _U757_in = _U759_out;
_U757_pt__U758 _U757 (
    .in(_U757_in),
    .out(_U757_out)
);
assign _U759_in = 16'(_U663_out * _U783_out);
assign _U759_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U759 (
    .in(_U759_in),
    .clk(_U759_clk),
    .out(_U759_out)
);
assign _U760_in = _U775_out;
_U760_pt__U761 _U760 (
    .in(_U760_in),
    .out(_U760_out)
);
assign _U762_in = in0_conv_stencil[0];
assign _U762_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U762 (
    .in(_U762_in),
    .clk(_U762_clk),
    .out(_U762_out)
);
assign _U763_in = _U762_out;
assign _U763_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U763 (
    .in(_U763_in),
    .clk(_U763_clk),
    .out(_U763_out)
);
assign _U764_in = _U763_out;
assign _U764_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U764 (
    .in(_U764_in),
    .clk(_U764_clk),
    .out(_U764_out)
);
assign _U765_in = _U764_out;
assign _U765_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U765 (
    .in(_U765_in),
    .clk(_U765_clk),
    .out(_U765_out)
);
assign _U766_in = _U765_out;
assign _U766_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U766 (
    .in(_U766_in),
    .clk(_U766_clk),
    .out(_U766_out)
);
assign _U767_in = _U766_out;
assign _U767_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U767 (
    .in(_U767_in),
    .clk(_U767_clk),
    .out(_U767_out)
);
assign _U768_in = _U767_out;
assign _U768_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U768 (
    .in(_U768_in),
    .clk(_U768_clk),
    .out(_U768_out)
);
assign _U769_in = _U768_out;
assign _U769_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U769 (
    .in(_U769_in),
    .clk(_U769_clk),
    .out(_U769_out)
);
assign _U770_in = _U769_out;
assign _U770_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U770 (
    .in(_U770_in),
    .clk(_U770_clk),
    .out(_U770_out)
);
assign _U771_in = _U770_out;
assign _U771_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U771 (
    .in(_U771_in),
    .clk(_U771_clk),
    .out(_U771_out)
);
assign _U772_in = _U771_out;
assign _U772_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U772 (
    .in(_U772_in),
    .clk(_U772_clk),
    .out(_U772_out)
);
assign _U773_in = _U772_out;
assign _U773_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U773 (
    .in(_U773_in),
    .clk(_U773_clk),
    .out(_U773_out)
);
assign _U774_in = _U773_out;
assign _U774_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U774 (
    .in(_U774_in),
    .clk(_U774_clk),
    .out(_U774_out)
);
assign _U775_in = _U774_out;
assign _U775_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U775 (
    .in(_U775_in),
    .clk(_U775_clk),
    .out(_U775_out)
);
assign _U776_in = _U779_out;
_U776_pt__U777 _U776 (
    .in(_U776_in),
    .out(_U776_out)
);
assign _U778_in = 16'(_U711_out * _U684_out);
assign _U778_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U778 (
    .in(_U778_in),
    .clk(_U778_clk),
    .out(_U778_out)
);
assign _U779_in = _U778_out;
assign _U779_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U779 (
    .in(_U779_in),
    .clk(_U779_clk),
    .out(_U779_out)
);
assign _U780_in = _U782_out;
_U780_pt__U781 _U780 (
    .in(_U780_in),
    .out(_U780_out)
);
assign _U782_in = 16'(_U735_out + _U807_out);
assign _U782_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U782 (
    .in(_U782_in),
    .clk(_U782_clk),
    .out(_U782_out)
);
assign _U783_in = _U791_out;
_U783_pt__U784 _U783 (
    .in(_U783_in),
    .out(_U783_out)
);
assign _U785_in = in1_hw_input_global_wrapper_stencil[7];
assign _U785_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U785 (
    .in(_U785_in),
    .clk(_U785_clk),
    .out(_U785_out)
);
assign _U786_in = _U785_out;
assign _U786_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U786 (
    .in(_U786_in),
    .clk(_U786_clk),
    .out(_U786_out)
);
assign _U787_in = _U786_out;
assign _U787_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U787 (
    .in(_U787_in),
    .clk(_U787_clk),
    .out(_U787_out)
);
assign _U788_in = _U787_out;
assign _U788_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U788 (
    .in(_U788_in),
    .clk(_U788_clk),
    .out(_U788_out)
);
assign _U789_in = _U788_out;
assign _U789_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U789 (
    .in(_U789_in),
    .clk(_U789_clk),
    .out(_U789_out)
);
assign _U790_in = _U789_out;
assign _U790_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U790 (
    .in(_U790_in),
    .clk(_U790_clk),
    .out(_U790_out)
);
assign _U791_in = _U790_out;
assign _U791_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U791 (
    .in(_U791_in),
    .clk(_U791_clk),
    .out(_U791_out)
);
assign _U792_in = _U794_out;
_U792_pt__U793 _U792 (
    .in(_U792_in),
    .out(_U792_out)
);
assign _U794_in = 16'(_U810_out + _U644_out);
assign _U794_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U794 (
    .in(_U794_in),
    .clk(_U794_clk),
    .out(_U794_out)
);
assign _U795_in = 16'(_U818_out + _U835_out);
_U795_pt__U796 _U795 (
    .in(_U795_in),
    .out(out_conv_stencil)
);
assign _U797_in = _U806_out;
_U797_pt__U798 _U797 (
    .in(_U797_in),
    .out(_U797_out)
);
assign _U799_in = 16'(_U653_out * _U752_out);
assign _U799_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U799 (
    .in(_U799_in),
    .clk(_U799_clk),
    .out(_U799_out)
);
assign _U800_in = _U799_out;
assign _U800_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U800 (
    .in(_U800_in),
    .clk(_U800_clk),
    .out(_U800_out)
);
assign _U801_in = _U800_out;
assign _U801_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U801 (
    .in(_U801_in),
    .clk(_U801_clk),
    .out(_U801_out)
);
assign _U802_in = _U801_out;
assign _U802_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U802 (
    .in(_U802_in),
    .clk(_U802_clk),
    .out(_U802_out)
);
assign _U803_in = _U802_out;
assign _U803_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U803 (
    .in(_U803_in),
    .clk(_U803_clk),
    .out(_U803_out)
);
assign _U804_in = _U803_out;
assign _U804_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U804 (
    .in(_U804_in),
    .clk(_U804_clk),
    .out(_U804_out)
);
assign _U805_in = _U804_out;
assign _U805_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U805 (
    .in(_U805_in),
    .clk(_U805_clk),
    .out(_U805_out)
);
assign _U806_in = _U805_out;
assign _U806_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U806 (
    .in(_U806_in),
    .clk(_U806_clk),
    .out(_U806_out)
);
assign _U807_in = _U809_out;
_U807_pt__U808 _U807 (
    .in(_U807_in),
    .out(_U807_out)
);
assign _U809_in = 16'(_U672_out + _U732_out);
assign _U809_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U809 (
    .in(_U809_in),
    .clk(_U809_clk),
    .out(_U809_out)
);
assign _U810_in = _U817_out;
_U810_pt__U811 _U810 (
    .in(_U810_in),
    .out(_U810_out)
);
assign _U812_in = 16'(_U692_out * _U647_out);
assign _U812_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U812 (
    .in(_U812_in),
    .clk(_U812_clk),
    .out(_U812_out)
);
assign _U813_in = _U812_out;
assign _U813_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U813 (
    .in(_U813_in),
    .clk(_U813_clk),
    .out(_U813_out)
);
assign _U814_in = _U813_out;
assign _U814_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U814 (
    .in(_U814_in),
    .clk(_U814_clk),
    .out(_U814_out)
);
assign _U815_in = _U814_out;
assign _U815_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U815 (
    .in(_U815_in),
    .clk(_U815_clk),
    .out(_U815_out)
);
assign _U816_in = _U815_out;
assign _U816_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U816 (
    .in(_U816_in),
    .clk(_U816_clk),
    .out(_U816_out)
);
assign _U817_in = _U816_out;
assign _U817_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U817 (
    .in(_U817_in),
    .clk(_U817_clk),
    .out(_U817_out)
);
assign _U818_in = _U834_out;
_U818_pt__U819 _U818 (
    .in(_U818_in),
    .out(_U818_out)
);
assign _U820_in = 16'(_U661_out * _U730_out);
assign _U820_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U820 (
    .in(_U820_in),
    .clk(_U820_clk),
    .out(_U820_out)
);
assign _U821_in = _U820_out;
assign _U821_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U821 (
    .in(_U821_in),
    .clk(_U821_clk),
    .out(_U821_out)
);
assign _U822_in = _U821_out;
assign _U822_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U822 (
    .in(_U822_in),
    .clk(_U822_clk),
    .out(_U822_out)
);
assign _U823_in = _U822_out;
assign _U823_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U823 (
    .in(_U823_in),
    .clk(_U823_clk),
    .out(_U823_out)
);
assign _U824_in = _U823_out;
assign _U824_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U824 (
    .in(_U824_in),
    .clk(_U824_clk),
    .out(_U824_out)
);
assign _U825_in = _U824_out;
assign _U825_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U825 (
    .in(_U825_in),
    .clk(_U825_clk),
    .out(_U825_out)
);
assign _U826_in = _U825_out;
assign _U826_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U826 (
    .in(_U826_in),
    .clk(_U826_clk),
    .out(_U826_out)
);
assign _U827_in = _U826_out;
assign _U827_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U827 (
    .in(_U827_in),
    .clk(_U827_clk),
    .out(_U827_out)
);
assign _U828_in = _U827_out;
assign _U828_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U828 (
    .in(_U828_in),
    .clk(_U828_clk),
    .out(_U828_out)
);
assign _U829_in = _U828_out;
assign _U829_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U829 (
    .in(_U829_in),
    .clk(_U829_clk),
    .out(_U829_out)
);
assign _U830_in = _U829_out;
assign _U830_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U830 (
    .in(_U830_in),
    .clk(_U830_clk),
    .out(_U830_out)
);
assign _U831_in = _U830_out;
assign _U831_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U831 (
    .in(_U831_in),
    .clk(_U831_clk),
    .out(_U831_out)
);
assign _U832_in = _U831_out;
assign _U832_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U832 (
    .in(_U832_in),
    .clk(_U832_clk),
    .out(_U832_out)
);
assign _U833_in = _U832_out;
assign _U833_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U833 (
    .in(_U833_in),
    .clk(_U833_clk),
    .out(_U833_out)
);
assign _U834_in = _U833_out;
assign _U834_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U834 (
    .in(_U834_in),
    .clk(_U834_clk),
    .out(_U834_out)
);
assign _U835_in = _U837_out;
_U835_pt__U836 _U835 (
    .in(_U835_in),
    .out(_U835_out)
);
assign _U837_in = 16'(_U760_out + _U780_out);
assign _U837_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U837 (
    .in(_U837_in),
    .clk(_U837_clk),
    .out(_U837_out)
);
endmodule

module cu_op_hcompute_conv_stencil_11 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_11_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_11_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_11_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[0];
hcompute_conv_stencil_11_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_11_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U630_pt__U631 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U623_pt__U624 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U61_pt__U62 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U615_pt__U616 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U607_pt__U608 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U603_pt__U604 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U599_pt__U600 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U596_pt__U597 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U593_pt__U594 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U587_pt__U588 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U581_pt__U582 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U579_pt__U580 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U577_pt__U578 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U572_pt__U573 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U56_pt__U57 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U567_pt__U568 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U558_pt__U559 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U549_pt__U550 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U533_pt__U534 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U528_pt__U529 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U524_pt__U525 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U521_pt__U522 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U51_pt__U52 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U512_pt__U513 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U509_pt__U510 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U4_pt__U5 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_2_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
wire [15:0] _U4_in;
assign _U4_in = in0_hw_input_stencil[0];
_U4_pt__U5 _U4 (
    .in(_U4_in),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil_2 (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read[0];
hcompute_hw_input_global_wrapper_stencil_2_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U498_pt__U499 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U495_pt__U496 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U492_pt__U493 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U489_pt__U490 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U487_pt__U488 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U47_pt__U48 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U478_pt__U479 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U475_pt__U476 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U472_pt__U473 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U460_pt__U461 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U446_pt__U447 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U43_pt__U44 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U436_pt__U437 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_10_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U436_in;
wire [15:0] _U436_out;
wire [15:0] _U438_in;
wire _U438_clk;
wire [15:0] _U438_out;
wire [15:0] _U439_in;
wire _U439_clk;
wire [15:0] _U439_out;
wire [15:0] _U440_in;
wire _U440_clk;
wire [15:0] _U440_out;
wire [15:0] _U441_in;
wire _U441_clk;
wire [15:0] _U441_out;
wire [15:0] _U442_in;
wire _U442_clk;
wire [15:0] _U442_out;
wire [15:0] _U443_in;
wire _U443_clk;
wire [15:0] _U443_out;
wire [15:0] _U444_in;
wire _U444_clk;
wire [15:0] _U444_out;
wire [15:0] _U445_in;
wire _U445_clk;
wire [15:0] _U445_out;
wire [15:0] _U446_in;
wire [15:0] _U446_out;
wire [15:0] _U448_in;
wire _U448_clk;
wire [15:0] _U448_out;
wire [15:0] _U449_in;
wire _U449_clk;
wire [15:0] _U449_out;
wire [15:0] _U450_in;
wire _U450_clk;
wire [15:0] _U450_out;
wire [15:0] _U451_in;
wire _U451_clk;
wire [15:0] _U451_out;
wire [15:0] _U452_in;
wire _U452_clk;
wire [15:0] _U452_out;
wire [15:0] _U453_in;
wire _U453_clk;
wire [15:0] _U453_out;
wire [15:0] _U454_in;
wire _U454_clk;
wire [15:0] _U454_out;
wire [15:0] _U455_in;
wire _U455_clk;
wire [15:0] _U455_out;
wire [15:0] _U456_in;
wire _U456_clk;
wire [15:0] _U456_out;
wire [15:0] _U457_in;
wire _U457_clk;
wire [15:0] _U457_out;
wire [15:0] _U458_in;
wire _U458_clk;
wire [15:0] _U458_out;
wire [15:0] _U459_in;
wire _U459_clk;
wire [15:0] _U459_out;
wire [15:0] _U460_in;
wire [15:0] _U460_out;
wire [15:0] _U462_in;
wire _U462_clk;
wire [15:0] _U462_out;
wire [15:0] _U463_in;
wire _U463_clk;
wire [15:0] _U463_out;
wire [15:0] _U464_in;
wire _U464_clk;
wire [15:0] _U464_out;
wire [15:0] _U465_in;
wire _U465_clk;
wire [15:0] _U465_out;
wire [15:0] _U466_in;
wire _U466_clk;
wire [15:0] _U466_out;
wire [15:0] _U467_in;
wire _U467_clk;
wire [15:0] _U467_out;
wire [15:0] _U468_in;
wire _U468_clk;
wire [15:0] _U468_out;
wire [15:0] _U469_in;
wire _U469_clk;
wire [15:0] _U469_out;
wire [15:0] _U470_in;
wire _U470_clk;
wire [15:0] _U470_out;
wire [15:0] _U471_in;
wire _U471_clk;
wire [15:0] _U471_out;
wire [15:0] _U472_in;
wire [15:0] _U472_out;
wire [15:0] _U474_in;
wire _U474_clk;
wire [15:0] _U474_out;
wire [15:0] _U475_in;
wire [15:0] _U475_out;
wire [15:0] _U477_in;
wire _U477_clk;
wire [15:0] _U477_out;
wire [15:0] _U478_in;
wire [15:0] _U478_out;
wire [15:0] _U480_in;
wire _U480_clk;
wire [15:0] _U480_out;
wire [15:0] _U481_in;
wire _U481_clk;
wire [15:0] _U481_out;
wire [15:0] _U482_in;
wire _U482_clk;
wire [15:0] _U482_out;
wire [15:0] _U483_in;
wire _U483_clk;
wire [15:0] _U483_out;
wire [15:0] _U484_in;
wire _U484_clk;
wire [15:0] _U484_out;
wire [15:0] _U485_in;
wire _U485_clk;
wire [15:0] _U485_out;
wire [15:0] _U486_in;
wire _U486_clk;
wire [15:0] _U486_out;
wire [15:0] _U487_in;
wire [15:0] _U489_in;
wire [15:0] _U489_out;
wire [15:0] _U491_in;
wire _U491_clk;
wire [15:0] _U491_out;
wire [15:0] _U492_in;
wire [15:0] _U492_out;
wire [15:0] _U494_in;
wire _U494_clk;
wire [15:0] _U494_out;
wire [15:0] _U495_in;
wire [15:0] _U495_out;
wire [15:0] _U497_in;
wire _U497_clk;
wire [15:0] _U497_out;
wire [15:0] _U498_in;
wire [15:0] _U498_out;
wire [15:0] _U500_in;
wire _U500_clk;
wire [15:0] _U500_out;
wire [15:0] _U501_in;
wire _U501_clk;
wire [15:0] _U501_out;
wire [15:0] _U502_in;
wire _U502_clk;
wire [15:0] _U502_out;
wire [15:0] _U503_in;
wire _U503_clk;
wire [15:0] _U503_out;
wire [15:0] _U504_in;
wire _U504_clk;
wire [15:0] _U504_out;
wire [15:0] _U505_in;
wire _U505_clk;
wire [15:0] _U505_out;
wire [15:0] _U506_in;
wire _U506_clk;
wire [15:0] _U506_out;
wire [15:0] _U507_in;
wire _U507_clk;
wire [15:0] _U507_out;
wire [15:0] _U508_in;
wire _U508_clk;
wire [15:0] _U508_out;
wire [15:0] _U509_in;
wire [15:0] _U509_out;
wire [15:0] _U511_in;
wire _U511_clk;
wire [15:0] _U511_out;
wire [15:0] _U512_in;
wire [15:0] _U512_out;
wire [15:0] _U514_in;
wire _U514_clk;
wire [15:0] _U514_out;
wire [15:0] _U515_in;
wire _U515_clk;
wire [15:0] _U515_out;
wire [15:0] _U516_in;
wire _U516_clk;
wire [15:0] _U516_out;
wire [15:0] _U517_in;
wire _U517_clk;
wire [15:0] _U517_out;
wire [15:0] _U518_in;
wire _U518_clk;
wire [15:0] _U518_out;
wire [15:0] _U519_in;
wire _U519_clk;
wire [15:0] _U519_out;
wire [15:0] _U520_in;
wire _U520_clk;
wire [15:0] _U520_out;
wire [15:0] _U521_in;
wire [15:0] _U521_out;
wire [15:0] _U523_in;
wire _U523_clk;
wire [15:0] _U523_out;
wire [15:0] _U524_in;
wire [15:0] _U524_out;
wire [15:0] _U526_in;
wire _U526_clk;
wire [15:0] _U526_out;
wire [15:0] _U527_in;
wire _U527_clk;
wire [15:0] _U527_out;
wire [15:0] _U528_in;
wire [15:0] _U528_out;
wire [15:0] _U530_in;
wire _U530_clk;
wire [15:0] _U530_out;
wire [15:0] _U531_in;
wire _U531_clk;
wire [15:0] _U531_out;
wire [15:0] _U532_in;
wire _U532_clk;
wire [15:0] _U532_out;
wire [15:0] _U533_in;
wire [15:0] _U533_out;
wire [15:0] _U535_in;
wire _U535_clk;
wire [15:0] _U535_out;
wire [15:0] _U536_in;
wire _U536_clk;
wire [15:0] _U536_out;
wire [15:0] _U537_in;
wire _U537_clk;
wire [15:0] _U537_out;
wire [15:0] _U538_in;
wire _U538_clk;
wire [15:0] _U538_out;
wire [15:0] _U539_in;
wire _U539_clk;
wire [15:0] _U539_out;
wire [15:0] _U540_in;
wire _U540_clk;
wire [15:0] _U540_out;
wire [15:0] _U541_in;
wire _U541_clk;
wire [15:0] _U541_out;
wire [15:0] _U542_in;
wire _U542_clk;
wire [15:0] _U542_out;
wire [15:0] _U543_in;
wire _U543_clk;
wire [15:0] _U543_out;
wire [15:0] _U544_in;
wire _U544_clk;
wire [15:0] _U544_out;
wire [15:0] _U545_in;
wire _U545_clk;
wire [15:0] _U545_out;
wire [15:0] _U546_in;
wire _U546_clk;
wire [15:0] _U546_out;
wire [15:0] _U547_in;
wire _U547_clk;
wire [15:0] _U547_out;
wire [15:0] _U548_in;
wire _U548_clk;
wire [15:0] _U548_out;
wire [15:0] _U549_in;
wire [15:0] _U549_out;
wire [15:0] _U551_in;
wire _U551_clk;
wire [15:0] _U551_out;
wire [15:0] _U552_in;
wire _U552_clk;
wire [15:0] _U552_out;
wire [15:0] _U553_in;
wire _U553_clk;
wire [15:0] _U553_out;
wire [15:0] _U554_in;
wire _U554_clk;
wire [15:0] _U554_out;
wire [15:0] _U555_in;
wire _U555_clk;
wire [15:0] _U555_out;
wire [15:0] _U556_in;
wire _U556_clk;
wire [15:0] _U556_out;
wire [15:0] _U557_in;
wire _U557_clk;
wire [15:0] _U557_out;
wire [15:0] _U558_in;
wire [15:0] _U558_out;
wire [15:0] _U560_in;
wire _U560_clk;
wire [15:0] _U560_out;
wire [15:0] _U561_in;
wire _U561_clk;
wire [15:0] _U561_out;
wire [15:0] _U562_in;
wire _U562_clk;
wire [15:0] _U562_out;
wire [15:0] _U563_in;
wire _U563_clk;
wire [15:0] _U563_out;
wire [15:0] _U564_in;
wire _U564_clk;
wire [15:0] _U564_out;
wire [15:0] _U565_in;
wire _U565_clk;
wire [15:0] _U565_out;
wire [15:0] _U566_in;
wire _U566_clk;
wire [15:0] _U566_out;
wire [15:0] _U567_in;
wire [15:0] _U567_out;
wire [15:0] _U569_in;
wire _U569_clk;
wire [15:0] _U569_out;
wire [15:0] _U570_in;
wire _U570_clk;
wire [15:0] _U570_out;
wire [15:0] _U571_in;
wire _U571_clk;
wire [15:0] _U571_out;
wire [15:0] _U572_in;
wire [15:0] _U572_out;
wire [15:0] _U574_in;
wire _U574_clk;
wire [15:0] _U574_out;
wire [15:0] _U575_in;
wire _U575_clk;
wire [15:0] _U575_out;
wire [15:0] _U576_in;
wire _U576_clk;
wire [15:0] _U576_out;
wire [15:0] _U577_in;
wire [15:0] _U577_out;
wire [15:0] _U579_in;
wire [15:0] _U579_out;
wire [15:0] _U581_in;
wire [15:0] _U581_out;
wire [15:0] _U583_in;
wire _U583_clk;
wire [15:0] _U583_out;
wire [15:0] _U584_in;
wire _U584_clk;
wire [15:0] _U584_out;
wire [15:0] _U585_in;
wire _U585_clk;
wire [15:0] _U585_out;
wire [15:0] _U586_in;
wire _U586_clk;
wire [15:0] _U586_out;
wire [15:0] _U587_in;
wire [15:0] _U587_out;
wire [15:0] _U589_in;
wire _U589_clk;
wire [15:0] _U589_out;
wire [15:0] _U590_in;
wire _U590_clk;
wire [15:0] _U590_out;
wire [15:0] _U591_in;
wire _U591_clk;
wire [15:0] _U591_out;
wire [15:0] _U592_in;
wire _U592_clk;
wire [15:0] _U592_out;
wire [15:0] _U593_in;
wire [15:0] _U593_out;
wire [15:0] _U595_in;
wire _U595_clk;
wire [15:0] _U595_out;
wire [15:0] _U596_in;
wire [15:0] _U596_out;
wire [15:0] _U598_in;
wire _U598_clk;
wire [15:0] _U598_out;
wire [15:0] _U599_in;
wire [15:0] _U599_out;
wire [15:0] _U601_in;
wire _U601_clk;
wire [15:0] _U601_out;
wire [15:0] _U602_in;
wire _U602_clk;
wire [15:0] _U602_out;
wire [15:0] _U603_in;
wire [15:0] _U603_out;
wire [15:0] _U605_in;
wire _U605_clk;
wire [15:0] _U605_out;
wire [15:0] _U606_in;
wire _U606_clk;
wire [15:0] _U606_out;
wire [15:0] _U607_in;
wire [15:0] _U607_out;
wire [15:0] _U609_in;
wire _U609_clk;
wire [15:0] _U609_out;
wire [15:0] _U610_in;
wire _U610_clk;
wire [15:0] _U610_out;
wire [15:0] _U611_in;
wire _U611_clk;
wire [15:0] _U611_out;
wire [15:0] _U612_in;
wire _U612_clk;
wire [15:0] _U612_out;
wire [15:0] _U613_in;
wire _U613_clk;
wire [15:0] _U613_out;
wire [15:0] _U614_in;
wire _U614_clk;
wire [15:0] _U614_out;
wire [15:0] _U615_in;
wire [15:0] _U615_out;
wire [15:0] _U617_in;
wire _U617_clk;
wire [15:0] _U617_out;
wire [15:0] _U618_in;
wire _U618_clk;
wire [15:0] _U618_out;
wire [15:0] _U619_in;
wire _U619_clk;
wire [15:0] _U619_out;
wire [15:0] _U620_in;
wire _U620_clk;
wire [15:0] _U620_out;
wire [15:0] _U621_in;
wire _U621_clk;
wire [15:0] _U621_out;
wire [15:0] _U622_in;
wire _U622_clk;
wire [15:0] _U622_out;
wire [15:0] _U623_in;
wire [15:0] _U623_out;
wire [15:0] _U625_in;
wire _U625_clk;
wire [15:0] _U625_out;
wire [15:0] _U626_in;
wire _U626_clk;
wire [15:0] _U626_out;
wire [15:0] _U627_in;
wire _U627_clk;
wire [15:0] _U627_out;
wire [15:0] _U628_in;
wire _U628_clk;
wire [15:0] _U628_out;
wire [15:0] _U629_in;
wire _U629_clk;
wire [15:0] _U629_out;
wire [15:0] _U630_in;
wire [15:0] _U630_out;
wire [15:0] _U632_in;
wire _U632_clk;
wire [15:0] _U632_out;
wire [15:0] _U633_in;
wire _U633_clk;
wire [15:0] _U633_out;
wire [15:0] _U634_in;
wire _U634_clk;
wire [15:0] _U634_out;
wire [15:0] _U635_in;
wire _U635_clk;
wire [15:0] _U635_out;
wire [15:0] _U636_in;
wire _U636_clk;
wire [15:0] _U636_out;
assign _U436_in = _U445_out;
_U436_pt__U437 _U436 (
    .in(_U436_in),
    .out(_U436_out)
);
assign _U438_in = 16'(_U549_out * _U558_out);
assign _U438_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U438 (
    .in(_U438_in),
    .clk(_U438_clk),
    .out(_U438_out)
);
assign _U439_in = _U438_out;
assign _U439_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U439 (
    .in(_U439_in),
    .clk(_U439_clk),
    .out(_U439_out)
);
assign _U440_in = _U439_out;
assign _U440_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U440 (
    .in(_U440_in),
    .clk(_U440_clk),
    .out(_U440_out)
);
assign _U441_in = _U440_out;
assign _U441_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U441 (
    .in(_U441_in),
    .clk(_U441_clk),
    .out(_U441_out)
);
assign _U442_in = _U441_out;
assign _U442_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U442 (
    .in(_U442_in),
    .clk(_U442_clk),
    .out(_U442_out)
);
assign _U443_in = _U442_out;
assign _U443_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U443 (
    .in(_U443_in),
    .clk(_U443_clk),
    .out(_U443_out)
);
assign _U444_in = _U443_out;
assign _U444_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U444 (
    .in(_U444_in),
    .clk(_U444_clk),
    .out(_U444_out)
);
assign _U445_in = _U444_out;
assign _U445_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U445 (
    .in(_U445_in),
    .clk(_U445_clk),
    .out(_U445_out)
);
assign _U446_in = _U459_out;
_U446_pt__U447 _U446 (
    .in(_U446_in),
    .out(_U446_out)
);
assign _U448_in = 16'(_U577_out * _U579_out);
assign _U448_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U448 (
    .in(_U448_in),
    .clk(_U448_clk),
    .out(_U448_out)
);
assign _U449_in = _U448_out;
assign _U449_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U449 (
    .in(_U449_in),
    .clk(_U449_clk),
    .out(_U449_out)
);
assign _U450_in = _U449_out;
assign _U450_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U450 (
    .in(_U450_in),
    .clk(_U450_clk),
    .out(_U450_out)
);
assign _U451_in = _U450_out;
assign _U451_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U451 (
    .in(_U451_in),
    .clk(_U451_clk),
    .out(_U451_out)
);
assign _U452_in = _U451_out;
assign _U452_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U452 (
    .in(_U452_in),
    .clk(_U452_clk),
    .out(_U452_out)
);
assign _U453_in = _U452_out;
assign _U453_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U453 (
    .in(_U453_in),
    .clk(_U453_clk),
    .out(_U453_out)
);
assign _U454_in = _U453_out;
assign _U454_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U454 (
    .in(_U454_in),
    .clk(_U454_clk),
    .out(_U454_out)
);
assign _U455_in = _U454_out;
assign _U455_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U455 (
    .in(_U455_in),
    .clk(_U455_clk),
    .out(_U455_out)
);
assign _U456_in = _U455_out;
assign _U456_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U456 (
    .in(_U456_in),
    .clk(_U456_clk),
    .out(_U456_out)
);
assign _U457_in = _U456_out;
assign _U457_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U457 (
    .in(_U457_in),
    .clk(_U457_clk),
    .out(_U457_out)
);
assign _U458_in = _U457_out;
assign _U458_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U458 (
    .in(_U458_in),
    .clk(_U458_clk),
    .out(_U458_out)
);
assign _U459_in = _U458_out;
assign _U459_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U459 (
    .in(_U459_in),
    .clk(_U459_clk),
    .out(_U459_out)
);
assign _U460_in = _U471_out;
_U460_pt__U461 _U460 (
    .in(_U460_in),
    .out(_U460_out)
);
assign _U462_in = 16'(_U567_out * _U572_out);
assign _U462_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U462 (
    .in(_U462_in),
    .clk(_U462_clk),
    .out(_U462_out)
);
assign _U463_in = _U462_out;
assign _U463_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U463 (
    .in(_U463_in),
    .clk(_U463_clk),
    .out(_U463_out)
);
assign _U464_in = _U463_out;
assign _U464_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U464 (
    .in(_U464_in),
    .clk(_U464_clk),
    .out(_U464_out)
);
assign _U465_in = _U464_out;
assign _U465_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U465 (
    .in(_U465_in),
    .clk(_U465_clk),
    .out(_U465_out)
);
assign _U466_in = _U465_out;
assign _U466_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U466 (
    .in(_U466_in),
    .clk(_U466_clk),
    .out(_U466_out)
);
assign _U467_in = _U466_out;
assign _U467_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U467 (
    .in(_U467_in),
    .clk(_U467_clk),
    .out(_U467_out)
);
assign _U468_in = _U467_out;
assign _U468_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U468 (
    .in(_U468_in),
    .clk(_U468_clk),
    .out(_U468_out)
);
assign _U469_in = _U468_out;
assign _U469_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U469 (
    .in(_U469_in),
    .clk(_U469_clk),
    .out(_U469_out)
);
assign _U470_in = _U469_out;
assign _U470_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U470 (
    .in(_U470_in),
    .clk(_U470_clk),
    .out(_U470_out)
);
assign _U471_in = _U470_out;
assign _U471_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U471 (
    .in(_U471_in),
    .clk(_U471_clk),
    .out(_U471_out)
);
assign _U472_in = _U474_out;
_U472_pt__U473 _U472 (
    .in(_U472_in),
    .out(_U472_out)
);
assign _U474_in = 16'(_U533_out + _U492_out);
assign _U474_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U474 (
    .in(_U474_in),
    .clk(_U474_clk),
    .out(_U474_out)
);
assign _U475_in = _U477_out;
_U475_pt__U476 _U475 (
    .in(_U475_in),
    .out(_U475_out)
);
assign _U477_in = 16'(_U478_out + _U495_out);
assign _U477_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U477 (
    .in(_U477_in),
    .clk(_U477_clk),
    .out(_U477_out)
);
assign _U478_in = _U486_out;
_U478_pt__U479 _U478 (
    .in(_U478_in),
    .out(_U478_out)
);
assign _U480_in = 16'(_U581_out * _U587_out);
assign _U480_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U480 (
    .in(_U480_in),
    .clk(_U480_clk),
    .out(_U480_out)
);
assign _U481_in = _U480_out;
assign _U481_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U481 (
    .in(_U481_in),
    .clk(_U481_clk),
    .out(_U481_out)
);
assign _U482_in = _U481_out;
assign _U482_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U482 (
    .in(_U482_in),
    .clk(_U482_clk),
    .out(_U482_out)
);
assign _U483_in = _U482_out;
assign _U483_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U483 (
    .in(_U483_in),
    .clk(_U483_clk),
    .out(_U483_out)
);
assign _U484_in = _U483_out;
assign _U484_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U484 (
    .in(_U484_in),
    .clk(_U484_clk),
    .out(_U484_out)
);
assign _U485_in = _U484_out;
assign _U485_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U485 (
    .in(_U485_in),
    .clk(_U485_clk),
    .out(_U485_out)
);
assign _U486_in = _U485_out;
assign _U486_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U486 (
    .in(_U486_in),
    .clk(_U486_clk),
    .out(_U486_out)
);
assign _U487_in = 16'(_U436_out + _U472_out);
_U487_pt__U488 _U487 (
    .in(_U487_in),
    .out(out_conv_stencil)
);
assign _U489_in = _U491_out;
_U489_pt__U490 _U489 (
    .in(_U489_in),
    .out(_U489_out)
);
assign _U491_in = 16'(_U446_out + _U475_out);
assign _U491_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U491 (
    .in(_U491_in),
    .clk(_U491_clk),
    .out(_U491_out)
);
assign _U492_in = _U494_out;
_U492_pt__U493 _U492 (
    .in(_U492_in),
    .out(_U492_out)
);
assign _U494_in = 16'(_U460_out + _U489_out);
assign _U494_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U494 (
    .in(_U494_in),
    .clk(_U494_clk),
    .out(_U494_out)
);
assign _U495_in = _U497_out;
_U495_pt__U496 _U495 (
    .in(_U495_in),
    .out(_U495_out)
);
assign _U497_in = 16'(_U498_out + _U509_out);
assign _U497_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U497 (
    .in(_U497_in),
    .clk(_U497_clk),
    .out(_U497_out)
);
assign _U498_in = _U508_out;
_U498_pt__U499 _U498 (
    .in(_U498_in),
    .out(_U498_out)
);
assign _U500_in = 16'(_U593_out * _U596_out);
assign _U500_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U500 (
    .in(_U500_in),
    .clk(_U500_clk),
    .out(_U500_out)
);
assign _U501_in = _U500_out;
assign _U501_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U501 (
    .in(_U501_in),
    .clk(_U501_clk),
    .out(_U501_out)
);
assign _U502_in = _U501_out;
assign _U502_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U502 (
    .in(_U502_in),
    .clk(_U502_clk),
    .out(_U502_out)
);
assign _U503_in = _U502_out;
assign _U503_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U503 (
    .in(_U503_in),
    .clk(_U503_clk),
    .out(_U503_out)
);
assign _U504_in = _U503_out;
assign _U504_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U504 (
    .in(_U504_in),
    .clk(_U504_clk),
    .out(_U504_out)
);
assign _U505_in = _U504_out;
assign _U505_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U505 (
    .in(_U505_in),
    .clk(_U505_clk),
    .out(_U505_out)
);
assign _U506_in = _U505_out;
assign _U506_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U506 (
    .in(_U506_in),
    .clk(_U506_clk),
    .out(_U506_out)
);
assign _U507_in = _U506_out;
assign _U507_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U507 (
    .in(_U507_in),
    .clk(_U507_clk),
    .out(_U507_out)
);
assign _U508_in = _U507_out;
assign _U508_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U508 (
    .in(_U508_in),
    .clk(_U508_clk),
    .out(_U508_out)
);
assign _U509_in = _U511_out;
_U509_pt__U510 _U509 (
    .in(_U509_in),
    .out(_U509_out)
);
assign _U511_in = 16'(_U512_out + _U521_out);
assign _U511_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U511 (
    .in(_U511_in),
    .clk(_U511_clk),
    .out(_U511_out)
);
assign _U512_in = _U520_out;
_U512_pt__U513 _U512 (
    .in(_U512_in),
    .out(_U512_out)
);
assign _U514_in = 16'(_U599_out * _U603_out);
assign _U514_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U514 (
    .in(_U514_in),
    .clk(_U514_clk),
    .out(_U514_out)
);
assign _U515_in = _U514_out;
assign _U515_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U515 (
    .in(_U515_in),
    .clk(_U515_clk),
    .out(_U515_out)
);
assign _U516_in = _U515_out;
assign _U516_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U516 (
    .in(_U516_in),
    .clk(_U516_clk),
    .out(_U516_out)
);
assign _U517_in = _U516_out;
assign _U517_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U517 (
    .in(_U517_in),
    .clk(_U517_clk),
    .out(_U517_out)
);
assign _U518_in = _U517_out;
assign _U518_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U518 (
    .in(_U518_in),
    .clk(_U518_clk),
    .out(_U518_out)
);
assign _U519_in = _U518_out;
assign _U519_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U519 (
    .in(_U519_in),
    .clk(_U519_clk),
    .out(_U519_out)
);
assign _U520_in = _U519_out;
assign _U520_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U520 (
    .in(_U520_in),
    .clk(_U520_clk),
    .out(_U520_out)
);
assign _U521_in = _U523_out;
_U521_pt__U522 _U521 (
    .in(_U521_in),
    .out(_U521_out)
);
assign _U523_in = 16'(_U524_out + _U528_out);
assign _U523_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U523 (
    .in(_U523_in),
    .clk(_U523_clk),
    .out(_U523_out)
);
assign _U524_in = _U527_out;
_U524_pt__U525 _U524 (
    .in(_U524_in),
    .out(_U524_out)
);
assign _U526_in = 16'(_U607_out * _U615_out);
assign _U526_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U526 (
    .in(_U526_in),
    .clk(_U526_clk),
    .out(_U526_out)
);
assign _U527_in = _U526_out;
assign _U527_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U527 (
    .in(_U527_in),
    .clk(_U527_clk),
    .out(_U527_out)
);
assign _U528_in = _U532_out;
_U528_pt__U529 _U528 (
    .in(_U528_in),
    .out(_U528_out)
);
assign _U530_in = 16'(_U623_out * _U630_out);
assign _U530_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U530 (
    .in(_U530_in),
    .clk(_U530_clk),
    .out(_U530_out)
);
assign _U531_in = _U530_out;
assign _U531_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U531 (
    .in(_U531_in),
    .clk(_U531_clk),
    .out(_U531_out)
);
assign _U532_in = _U531_out;
assign _U532_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U532 (
    .in(_U532_in),
    .clk(_U532_clk),
    .out(_U532_out)
);
assign _U533_in = _U548_out;
_U533_pt__U534 _U533 (
    .in(_U533_in),
    .out(_U533_out)
);
assign _U535_in = in0_conv_stencil[0];
assign _U535_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U535 (
    .in(_U535_in),
    .clk(_U535_clk),
    .out(_U535_out)
);
assign _U536_in = _U535_out;
assign _U536_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U536 (
    .in(_U536_in),
    .clk(_U536_clk),
    .out(_U536_out)
);
assign _U537_in = _U536_out;
assign _U537_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U537 (
    .in(_U537_in),
    .clk(_U537_clk),
    .out(_U537_out)
);
assign _U538_in = _U537_out;
assign _U538_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U538 (
    .in(_U538_in),
    .clk(_U538_clk),
    .out(_U538_out)
);
assign _U539_in = _U538_out;
assign _U539_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U539 (
    .in(_U539_in),
    .clk(_U539_clk),
    .out(_U539_out)
);
assign _U540_in = _U539_out;
assign _U540_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U540 (
    .in(_U540_in),
    .clk(_U540_clk),
    .out(_U540_out)
);
assign _U541_in = _U540_out;
assign _U541_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U541 (
    .in(_U541_in),
    .clk(_U541_clk),
    .out(_U541_out)
);
assign _U542_in = _U541_out;
assign _U542_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U542 (
    .in(_U542_in),
    .clk(_U542_clk),
    .out(_U542_out)
);
assign _U543_in = _U542_out;
assign _U543_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U543 (
    .in(_U543_in),
    .clk(_U543_clk),
    .out(_U543_out)
);
assign _U544_in = _U543_out;
assign _U544_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U544 (
    .in(_U544_in),
    .clk(_U544_clk),
    .out(_U544_out)
);
assign _U545_in = _U544_out;
assign _U545_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U545 (
    .in(_U545_in),
    .clk(_U545_clk),
    .out(_U545_out)
);
assign _U546_in = _U545_out;
assign _U546_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U546 (
    .in(_U546_in),
    .clk(_U546_clk),
    .out(_U546_out)
);
assign _U547_in = _U546_out;
assign _U547_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U547 (
    .in(_U547_in),
    .clk(_U547_clk),
    .out(_U547_out)
);
assign _U548_in = _U547_out;
assign _U548_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U548 (
    .in(_U548_in),
    .clk(_U548_clk),
    .out(_U548_out)
);
assign _U549_in = _U557_out;
_U549_pt__U550 _U549 (
    .in(_U549_in),
    .out(_U549_out)
);
assign _U551_in = in2_hw_kernel_global_wrapper_stencil[0];
assign _U551_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U551 (
    .in(_U551_in),
    .clk(_U551_clk),
    .out(_U551_out)
);
assign _U552_in = _U551_out;
assign _U552_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U552 (
    .in(_U552_in),
    .clk(_U552_clk),
    .out(_U552_out)
);
assign _U553_in = _U552_out;
assign _U553_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U553 (
    .in(_U553_in),
    .clk(_U553_clk),
    .out(_U553_out)
);
assign _U554_in = _U553_out;
assign _U554_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U554 (
    .in(_U554_in),
    .clk(_U554_clk),
    .out(_U554_out)
);
assign _U555_in = _U554_out;
assign _U555_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U555 (
    .in(_U555_in),
    .clk(_U555_clk),
    .out(_U555_out)
);
assign _U556_in = _U555_out;
assign _U556_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U556 (
    .in(_U556_in),
    .clk(_U556_clk),
    .out(_U556_out)
);
assign _U557_in = _U556_out;
assign _U557_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U557 (
    .in(_U557_in),
    .clk(_U557_clk),
    .out(_U557_out)
);
assign _U558_in = _U566_out;
_U558_pt__U559 _U558 (
    .in(_U558_in),
    .out(_U558_out)
);
assign _U560_in = in1_hw_input_global_wrapper_stencil[0];
assign _U560_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U560 (
    .in(_U560_in),
    .clk(_U560_clk),
    .out(_U560_out)
);
assign _U561_in = _U560_out;
assign _U561_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U561 (
    .in(_U561_in),
    .clk(_U561_clk),
    .out(_U561_out)
);
assign _U562_in = _U561_out;
assign _U562_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U562 (
    .in(_U562_in),
    .clk(_U562_clk),
    .out(_U562_out)
);
assign _U563_in = _U562_out;
assign _U563_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U563 (
    .in(_U563_in),
    .clk(_U563_clk),
    .out(_U563_out)
);
assign _U564_in = _U563_out;
assign _U564_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U564 (
    .in(_U564_in),
    .clk(_U564_clk),
    .out(_U564_out)
);
assign _U565_in = _U564_out;
assign _U565_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U565 (
    .in(_U565_in),
    .clk(_U565_clk),
    .out(_U565_out)
);
assign _U566_in = _U565_out;
assign _U566_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U566 (
    .in(_U566_in),
    .clk(_U566_clk),
    .out(_U566_out)
);
assign _U567_in = _U571_out;
_U567_pt__U568 _U567 (
    .in(_U567_in),
    .out(_U567_out)
);
assign _U569_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U569_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U569 (
    .in(_U569_in),
    .clk(_U569_clk),
    .out(_U569_out)
);
assign _U570_in = _U569_out;
assign _U570_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U570 (
    .in(_U570_in),
    .clk(_U570_clk),
    .out(_U570_out)
);
assign _U571_in = _U570_out;
assign _U571_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U571 (
    .in(_U571_in),
    .clk(_U571_clk),
    .out(_U571_out)
);
assign _U572_in = _U576_out;
_U572_pt__U573 _U572 (
    .in(_U572_in),
    .out(_U572_out)
);
assign _U574_in = in1_hw_input_global_wrapper_stencil[1];
assign _U574_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U574 (
    .in(_U574_in),
    .clk(_U574_clk),
    .out(_U574_out)
);
assign _U575_in = _U574_out;
assign _U575_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U575 (
    .in(_U575_in),
    .clk(_U575_clk),
    .out(_U575_out)
);
assign _U576_in = _U575_out;
assign _U576_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U576 (
    .in(_U576_in),
    .clk(_U576_clk),
    .out(_U576_out)
);
assign _U577_in = in2_hw_kernel_global_wrapper_stencil[2];
_U577_pt__U578 _U577 (
    .in(_U577_in),
    .out(_U577_out)
);
assign _U579_in = in1_hw_input_global_wrapper_stencil[2];
_U579_pt__U580 _U579 (
    .in(_U579_in),
    .out(_U579_out)
);
assign _U581_in = _U586_out;
_U581_pt__U582 _U581 (
    .in(_U581_in),
    .out(_U581_out)
);
assign _U583_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U583_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U583 (
    .in(_U583_in),
    .clk(_U583_clk),
    .out(_U583_out)
);
assign _U584_in = _U583_out;
assign _U584_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U584 (
    .in(_U584_in),
    .clk(_U584_clk),
    .out(_U584_out)
);
assign _U585_in = _U584_out;
assign _U585_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U585 (
    .in(_U585_in),
    .clk(_U585_clk),
    .out(_U585_out)
);
assign _U586_in = _U585_out;
assign _U586_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U586 (
    .in(_U586_in),
    .clk(_U586_clk),
    .out(_U586_out)
);
assign _U587_in = _U592_out;
_U587_pt__U588 _U587 (
    .in(_U587_in),
    .out(_U587_out)
);
assign _U589_in = in1_hw_input_global_wrapper_stencil[3];
assign _U589_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U589 (
    .in(_U589_in),
    .clk(_U589_clk),
    .out(_U589_out)
);
assign _U590_in = _U589_out;
assign _U590_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U590 (
    .in(_U590_in),
    .clk(_U590_clk),
    .out(_U590_out)
);
assign _U591_in = _U590_out;
assign _U591_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U591 (
    .in(_U591_in),
    .clk(_U591_clk),
    .out(_U591_out)
);
assign _U592_in = _U591_out;
assign _U592_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U592 (
    .in(_U592_in),
    .clk(_U592_clk),
    .out(_U592_out)
);
assign _U593_in = _U595_out;
_U593_pt__U594 _U593 (
    .in(_U593_in),
    .out(_U593_out)
);
assign _U595_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U595_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U595 (
    .in(_U595_in),
    .clk(_U595_clk),
    .out(_U595_out)
);
assign _U596_in = _U598_out;
_U596_pt__U597 _U596 (
    .in(_U596_in),
    .out(_U596_out)
);
assign _U598_in = in1_hw_input_global_wrapper_stencil[4];
assign _U598_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U598 (
    .in(_U598_in),
    .clk(_U598_clk),
    .out(_U598_out)
);
assign _U599_in = _U602_out;
_U599_pt__U600 _U599 (
    .in(_U599_in),
    .out(_U599_out)
);
assign _U601_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U601_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U601 (
    .in(_U601_in),
    .clk(_U601_clk),
    .out(_U601_out)
);
assign _U602_in = _U601_out;
assign _U602_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U602 (
    .in(_U602_in),
    .clk(_U602_clk),
    .out(_U602_out)
);
assign _U603_in = _U606_out;
_U603_pt__U604 _U603 (
    .in(_U603_in),
    .out(_U603_out)
);
assign _U605_in = in1_hw_input_global_wrapper_stencil[5];
assign _U605_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U605 (
    .in(_U605_in),
    .clk(_U605_clk),
    .out(_U605_out)
);
assign _U606_in = _U605_out;
assign _U606_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U606 (
    .in(_U606_in),
    .clk(_U606_clk),
    .out(_U606_out)
);
assign _U607_in = _U614_out;
_U607_pt__U608 _U607 (
    .in(_U607_in),
    .out(_U607_out)
);
assign _U609_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U609_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U609 (
    .in(_U609_in),
    .clk(_U609_clk),
    .out(_U609_out)
);
assign _U610_in = _U609_out;
assign _U610_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U610 (
    .in(_U610_in),
    .clk(_U610_clk),
    .out(_U610_out)
);
assign _U611_in = _U610_out;
assign _U611_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U611 (
    .in(_U611_in),
    .clk(_U611_clk),
    .out(_U611_out)
);
assign _U612_in = _U611_out;
assign _U612_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U612 (
    .in(_U612_in),
    .clk(_U612_clk),
    .out(_U612_out)
);
assign _U613_in = _U612_out;
assign _U613_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U613 (
    .in(_U613_in),
    .clk(_U613_clk),
    .out(_U613_out)
);
assign _U614_in = _U613_out;
assign _U614_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U614 (
    .in(_U614_in),
    .clk(_U614_clk),
    .out(_U614_out)
);
assign _U615_in = _U622_out;
_U615_pt__U616 _U615 (
    .in(_U615_in),
    .out(_U615_out)
);
assign _U617_in = in1_hw_input_global_wrapper_stencil[6];
assign _U617_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U617 (
    .in(_U617_in),
    .clk(_U617_clk),
    .out(_U617_out)
);
assign _U618_in = _U617_out;
assign _U618_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U618 (
    .in(_U618_in),
    .clk(_U618_clk),
    .out(_U618_out)
);
assign _U619_in = _U618_out;
assign _U619_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U619 (
    .in(_U619_in),
    .clk(_U619_clk),
    .out(_U619_out)
);
assign _U620_in = _U619_out;
assign _U620_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U620 (
    .in(_U620_in),
    .clk(_U620_clk),
    .out(_U620_out)
);
assign _U621_in = _U620_out;
assign _U621_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U621 (
    .in(_U621_in),
    .clk(_U621_clk),
    .out(_U621_out)
);
assign _U622_in = _U621_out;
assign _U622_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U622 (
    .in(_U622_in),
    .clk(_U622_clk),
    .out(_U622_out)
);
assign _U623_in = _U629_out;
_U623_pt__U624 _U623 (
    .in(_U623_in),
    .out(_U623_out)
);
assign _U625_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U625_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U625 (
    .in(_U625_in),
    .clk(_U625_clk),
    .out(_U625_out)
);
assign _U626_in = _U625_out;
assign _U626_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U626 (
    .in(_U626_in),
    .clk(_U626_clk),
    .out(_U626_out)
);
assign _U627_in = _U626_out;
assign _U627_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U627 (
    .in(_U627_in),
    .clk(_U627_clk),
    .out(_U627_out)
);
assign _U628_in = _U627_out;
assign _U628_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U628 (
    .in(_U628_in),
    .clk(_U628_clk),
    .out(_U628_out)
);
assign _U629_in = _U628_out;
assign _U629_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U629 (
    .in(_U629_in),
    .clk(_U629_clk),
    .out(_U629_out)
);
assign _U630_in = _U636_out;
_U630_pt__U631 _U630 (
    .in(_U630_in),
    .out(_U630_out)
);
assign _U632_in = in1_hw_input_global_wrapper_stencil[7];
assign _U632_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U632 (
    .in(_U632_in),
    .clk(_U632_clk),
    .out(_U632_out)
);
assign _U633_in = _U632_out;
assign _U633_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U633 (
    .in(_U633_in),
    .clk(_U633_clk),
    .out(_U633_out)
);
assign _U634_in = _U633_out;
assign _U634_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U634 (
    .in(_U634_in),
    .clk(_U634_clk),
    .out(_U634_out)
);
assign _U635_in = _U634_out;
assign _U635_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U635 (
    .in(_U635_in),
    .clk(_U635_clk),
    .out(_U635_out)
);
assign _U636_in = _U635_out;
assign _U636_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U636 (
    .in(_U636_in),
    .clk(_U636_clk),
    .out(_U636_out)
);
endmodule

module cu_op_hcompute_conv_stencil_10 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_10_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_10_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_10_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[0];
hcompute_conv_stencil_10_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_10_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U431_pt__U432 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U426_pt__U427 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U424_pt__U425 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U422_pt__U423 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U418_pt__U419 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U414_pt__U415 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U40_pt__U41 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U407_pt__U408 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U400_pt__U401 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U394_pt__U395 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U388_pt__U389 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U385_pt__U386 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U382_pt__U383 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U37_pt__U38 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U373_pt__U374 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U364_pt__U365 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U356_pt__U357 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U34_pt__U35 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U348_pt__U349 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U332_pt__U333 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U32_pt__U33 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_7_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U32_in;
assign _U32_in = 16'h0000;
_U32_pt__U33 _U32 (
    .in(_U32_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_7 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_7_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_7_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_7_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U322_pt__U323 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U319_pt__U320 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U316_pt__U317 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U30_pt__U31 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_6_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U30_in;
assign _U30_in = 16'h0000;
_U30_pt__U31 _U30 (
    .in(_U30_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_6 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_6_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_6_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_6_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U302_pt__U303 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U2_pt__U3 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_1_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
wire [15:0] _U2_in;
assign _U2_in = in0_hw_input_stencil[0];
_U2_pt__U3 _U2 (
    .in(_U2_in),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil_1 (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read[0];
hcompute_hw_input_global_wrapper_stencil_1_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U299_pt__U300 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U296_pt__U297 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U293_pt__U294 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U290_pt__U291 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U28_pt__U29 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_5_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U28_in;
assign _U28_in = 16'h0000;
_U28_pt__U29 _U28 (
    .in(_U28_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_5 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_5_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U282_pt__U283 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U276_pt__U277 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U26_pt__U27 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_4_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U26_in;
assign _U26_in = 16'h0000;
_U26_pt__U27 _U26 (
    .in(_U26_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_4 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_4_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U268_pt__U269 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U266_pt__U267 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U263_pt__U264 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U254_pt__U255 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U24_pt__U25 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_3_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U24_in;
assign _U24_in = 16'h0000;
_U24_pt__U25 _U24 (
    .in(_U24_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_3 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_3_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U247_pt__U248 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U235_pt__U236 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_9_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U235_in;
wire [15:0] _U235_out;
wire [15:0] _U237_in;
wire _U237_clk;
wire [15:0] _U237_out;
wire [15:0] _U238_in;
wire _U238_clk;
wire [15:0] _U238_out;
wire [15:0] _U239_in;
wire _U239_clk;
wire [15:0] _U239_out;
wire [15:0] _U240_in;
wire _U240_clk;
wire [15:0] _U240_out;
wire [15:0] _U241_in;
wire _U241_clk;
wire [15:0] _U241_out;
wire [15:0] _U242_in;
wire _U242_clk;
wire [15:0] _U242_out;
wire [15:0] _U243_in;
wire _U243_clk;
wire [15:0] _U243_out;
wire [15:0] _U244_in;
wire _U244_clk;
wire [15:0] _U244_out;
wire [15:0] _U245_in;
wire _U245_clk;
wire [15:0] _U245_out;
wire [15:0] _U246_in;
wire _U246_clk;
wire [15:0] _U246_out;
wire [15:0] _U247_in;
wire [15:0] _U247_out;
wire [15:0] _U249_in;
wire _U249_clk;
wire [15:0] _U249_out;
wire [15:0] _U250_in;
wire _U250_clk;
wire [15:0] _U250_out;
wire [15:0] _U251_in;
wire _U251_clk;
wire [15:0] _U251_out;
wire [15:0] _U252_in;
wire _U252_clk;
wire [15:0] _U252_out;
wire [15:0] _U253_in;
wire _U253_clk;
wire [15:0] _U253_out;
wire [15:0] _U254_in;
wire [15:0] _U254_out;
wire [15:0] _U256_in;
wire _U256_clk;
wire [15:0] _U256_out;
wire [15:0] _U257_in;
wire _U257_clk;
wire [15:0] _U257_out;
wire [15:0] _U258_in;
wire _U258_clk;
wire [15:0] _U258_out;
wire [15:0] _U259_in;
wire _U259_clk;
wire [15:0] _U259_out;
wire [15:0] _U260_in;
wire _U260_clk;
wire [15:0] _U260_out;
wire [15:0] _U261_in;
wire _U261_clk;
wire [15:0] _U261_out;
wire [15:0] _U262_in;
wire _U262_clk;
wire [15:0] _U262_out;
wire [15:0] _U263_in;
wire [15:0] _U263_out;
wire [15:0] _U265_in;
wire _U265_clk;
wire [15:0] _U265_out;
wire [15:0] _U266_in;
wire [15:0] _U268_in;
wire [15:0] _U268_out;
wire [15:0] _U270_in;
wire _U270_clk;
wire [15:0] _U270_out;
wire [15:0] _U271_in;
wire _U271_clk;
wire [15:0] _U271_out;
wire [15:0] _U272_in;
wire _U272_clk;
wire [15:0] _U272_out;
wire [15:0] _U273_in;
wire _U273_clk;
wire [15:0] _U273_out;
wire [15:0] _U274_in;
wire _U274_clk;
wire [15:0] _U274_out;
wire [15:0] _U275_in;
wire _U275_clk;
wire [15:0] _U275_out;
wire [15:0] _U276_in;
wire [15:0] _U276_out;
wire [15:0] _U278_in;
wire _U278_clk;
wire [15:0] _U278_out;
wire [15:0] _U279_in;
wire _U279_clk;
wire [15:0] _U279_out;
wire [15:0] _U280_in;
wire _U280_clk;
wire [15:0] _U280_out;
wire [15:0] _U281_in;
wire _U281_clk;
wire [15:0] _U281_out;
wire [15:0] _U282_in;
wire [15:0] _U282_out;
wire [15:0] _U284_in;
wire _U284_clk;
wire [15:0] _U284_out;
wire [15:0] _U285_in;
wire _U285_clk;
wire [15:0] _U285_out;
wire [15:0] _U286_in;
wire _U286_clk;
wire [15:0] _U286_out;
wire [15:0] _U287_in;
wire _U287_clk;
wire [15:0] _U287_out;
wire [15:0] _U288_in;
wire _U288_clk;
wire [15:0] _U288_out;
wire [15:0] _U289_in;
wire _U289_clk;
wire [15:0] _U289_out;
wire [15:0] _U290_in;
wire [15:0] _U290_out;
wire [15:0] _U292_in;
wire _U292_clk;
wire [15:0] _U292_out;
wire [15:0] _U293_in;
wire [15:0] _U293_out;
wire [15:0] _U295_in;
wire _U295_clk;
wire [15:0] _U295_out;
wire [15:0] _U296_in;
wire [15:0] _U296_out;
wire [15:0] _U298_in;
wire _U298_clk;
wire [15:0] _U298_out;
wire [15:0] _U299_in;
wire [15:0] _U299_out;
wire [15:0] _U301_in;
wire _U301_clk;
wire [15:0] _U301_out;
wire [15:0] _U302_in;
wire [15:0] _U302_out;
wire [15:0] _U304_in;
wire _U304_clk;
wire [15:0] _U304_out;
wire [15:0] _U305_in;
wire _U305_clk;
wire [15:0] _U305_out;
wire [15:0] _U306_in;
wire _U306_clk;
wire [15:0] _U306_out;
wire [15:0] _U307_in;
wire _U307_clk;
wire [15:0] _U307_out;
wire [15:0] _U308_in;
wire _U308_clk;
wire [15:0] _U308_out;
wire [15:0] _U309_in;
wire _U309_clk;
wire [15:0] _U309_out;
wire [15:0] _U310_in;
wire _U310_clk;
wire [15:0] _U310_out;
wire [15:0] _U311_in;
wire _U311_clk;
wire [15:0] _U311_out;
wire [15:0] _U312_in;
wire _U312_clk;
wire [15:0] _U312_out;
wire [15:0] _U313_in;
wire _U313_clk;
wire [15:0] _U313_out;
wire [15:0] _U314_in;
wire _U314_clk;
wire [15:0] _U314_out;
wire [15:0] _U315_in;
wire _U315_clk;
wire [15:0] _U315_out;
wire [15:0] _U316_in;
wire [15:0] _U316_out;
wire [15:0] _U318_in;
wire _U318_clk;
wire [15:0] _U318_out;
wire [15:0] _U319_in;
wire [15:0] _U319_out;
wire [15:0] _U321_in;
wire _U321_clk;
wire [15:0] _U321_out;
wire [15:0] _U322_in;
wire [15:0] _U322_out;
wire [15:0] _U324_in;
wire _U324_clk;
wire [15:0] _U324_out;
wire [15:0] _U325_in;
wire _U325_clk;
wire [15:0] _U325_out;
wire [15:0] _U326_in;
wire _U326_clk;
wire [15:0] _U326_out;
wire [15:0] _U327_in;
wire _U327_clk;
wire [15:0] _U327_out;
wire [15:0] _U328_in;
wire _U328_clk;
wire [15:0] _U328_out;
wire [15:0] _U329_in;
wire _U329_clk;
wire [15:0] _U329_out;
wire [15:0] _U330_in;
wire _U330_clk;
wire [15:0] _U330_out;
wire [15:0] _U331_in;
wire _U331_clk;
wire [15:0] _U331_out;
wire [15:0] _U332_in;
wire [15:0] _U332_out;
wire [15:0] _U334_in;
wire _U334_clk;
wire [15:0] _U334_out;
wire [15:0] _U335_in;
wire _U335_clk;
wire [15:0] _U335_out;
wire [15:0] _U336_in;
wire _U336_clk;
wire [15:0] _U336_out;
wire [15:0] _U337_in;
wire _U337_clk;
wire [15:0] _U337_out;
wire [15:0] _U338_in;
wire _U338_clk;
wire [15:0] _U338_out;
wire [15:0] _U339_in;
wire _U339_clk;
wire [15:0] _U339_out;
wire [15:0] _U340_in;
wire _U340_clk;
wire [15:0] _U340_out;
wire [15:0] _U341_in;
wire _U341_clk;
wire [15:0] _U341_out;
wire [15:0] _U342_in;
wire _U342_clk;
wire [15:0] _U342_out;
wire [15:0] _U343_in;
wire _U343_clk;
wire [15:0] _U343_out;
wire [15:0] _U344_in;
wire _U344_clk;
wire [15:0] _U344_out;
wire [15:0] _U345_in;
wire _U345_clk;
wire [15:0] _U345_out;
wire [15:0] _U346_in;
wire _U346_clk;
wire [15:0] _U346_out;
wire [15:0] _U347_in;
wire _U347_clk;
wire [15:0] _U347_out;
wire [15:0] _U348_in;
wire [15:0] _U348_out;
wire [15:0] _U350_in;
wire _U350_clk;
wire [15:0] _U350_out;
wire [15:0] _U351_in;
wire _U351_clk;
wire [15:0] _U351_out;
wire [15:0] _U352_in;
wire _U352_clk;
wire [15:0] _U352_out;
wire [15:0] _U353_in;
wire _U353_clk;
wire [15:0] _U353_out;
wire [15:0] _U354_in;
wire _U354_clk;
wire [15:0] _U354_out;
wire [15:0] _U355_in;
wire _U355_clk;
wire [15:0] _U355_out;
wire [15:0] _U356_in;
wire [15:0] _U356_out;
wire [15:0] _U358_in;
wire _U358_clk;
wire [15:0] _U358_out;
wire [15:0] _U359_in;
wire _U359_clk;
wire [15:0] _U359_out;
wire [15:0] _U360_in;
wire _U360_clk;
wire [15:0] _U360_out;
wire [15:0] _U361_in;
wire _U361_clk;
wire [15:0] _U361_out;
wire [15:0] _U362_in;
wire _U362_clk;
wire [15:0] _U362_out;
wire [15:0] _U363_in;
wire _U363_clk;
wire [15:0] _U363_out;
wire [15:0] _U364_in;
wire [15:0] _U364_out;
wire [15:0] _U366_in;
wire _U366_clk;
wire [15:0] _U366_out;
wire [15:0] _U367_in;
wire _U367_clk;
wire [15:0] _U367_out;
wire [15:0] _U368_in;
wire _U368_clk;
wire [15:0] _U368_out;
wire [15:0] _U369_in;
wire _U369_clk;
wire [15:0] _U369_out;
wire [15:0] _U370_in;
wire _U370_clk;
wire [15:0] _U370_out;
wire [15:0] _U371_in;
wire _U371_clk;
wire [15:0] _U371_out;
wire [15:0] _U372_in;
wire _U372_clk;
wire [15:0] _U372_out;
wire [15:0] _U373_in;
wire [15:0] _U373_out;
wire [15:0] _U375_in;
wire _U375_clk;
wire [15:0] _U375_out;
wire [15:0] _U376_in;
wire _U376_clk;
wire [15:0] _U376_out;
wire [15:0] _U377_in;
wire _U377_clk;
wire [15:0] _U377_out;
wire [15:0] _U378_in;
wire _U378_clk;
wire [15:0] _U378_out;
wire [15:0] _U379_in;
wire _U379_clk;
wire [15:0] _U379_out;
wire [15:0] _U380_in;
wire _U380_clk;
wire [15:0] _U380_out;
wire [15:0] _U381_in;
wire _U381_clk;
wire [15:0] _U381_out;
wire [15:0] _U382_in;
wire [15:0] _U382_out;
wire [15:0] _U384_in;
wire _U384_clk;
wire [15:0] _U384_out;
wire [15:0] _U385_in;
wire [15:0] _U385_out;
wire [15:0] _U387_in;
wire _U387_clk;
wire [15:0] _U387_out;
wire [15:0] _U388_in;
wire [15:0] _U388_out;
wire [15:0] _U390_in;
wire _U390_clk;
wire [15:0] _U390_out;
wire [15:0] _U391_in;
wire _U391_clk;
wire [15:0] _U391_out;
wire [15:0] _U392_in;
wire _U392_clk;
wire [15:0] _U392_out;
wire [15:0] _U393_in;
wire _U393_clk;
wire [15:0] _U393_out;
wire [15:0] _U394_in;
wire [15:0] _U394_out;
wire [15:0] _U396_in;
wire _U396_clk;
wire [15:0] _U396_out;
wire [15:0] _U397_in;
wire _U397_clk;
wire [15:0] _U397_out;
wire [15:0] _U398_in;
wire _U398_clk;
wire [15:0] _U398_out;
wire [15:0] _U399_in;
wire _U399_clk;
wire [15:0] _U399_out;
wire [15:0] _U400_in;
wire [15:0] _U400_out;
wire [15:0] _U402_in;
wire _U402_clk;
wire [15:0] _U402_out;
wire [15:0] _U403_in;
wire _U403_clk;
wire [15:0] _U403_out;
wire [15:0] _U404_in;
wire _U404_clk;
wire [15:0] _U404_out;
wire [15:0] _U405_in;
wire _U405_clk;
wire [15:0] _U405_out;
wire [15:0] _U406_in;
wire _U406_clk;
wire [15:0] _U406_out;
wire [15:0] _U407_in;
wire [15:0] _U407_out;
wire [15:0] _U409_in;
wire _U409_clk;
wire [15:0] _U409_out;
wire [15:0] _U410_in;
wire _U410_clk;
wire [15:0] _U410_out;
wire [15:0] _U411_in;
wire _U411_clk;
wire [15:0] _U411_out;
wire [15:0] _U412_in;
wire _U412_clk;
wire [15:0] _U412_out;
wire [15:0] _U413_in;
wire _U413_clk;
wire [15:0] _U413_out;
wire [15:0] _U414_in;
wire [15:0] _U414_out;
wire [15:0] _U416_in;
wire _U416_clk;
wire [15:0] _U416_out;
wire [15:0] _U417_in;
wire _U417_clk;
wire [15:0] _U417_out;
wire [15:0] _U418_in;
wire [15:0] _U418_out;
wire [15:0] _U420_in;
wire _U420_clk;
wire [15:0] _U420_out;
wire [15:0] _U421_in;
wire _U421_clk;
wire [15:0] _U421_out;
wire [15:0] _U422_in;
wire [15:0] _U422_out;
wire [15:0] _U424_in;
wire [15:0] _U424_out;
wire [15:0] _U426_in;
wire [15:0] _U426_out;
wire [15:0] _U428_in;
wire _U428_clk;
wire [15:0] _U428_out;
wire [15:0] _U429_in;
wire _U429_clk;
wire [15:0] _U429_out;
wire [15:0] _U430_in;
wire _U430_clk;
wire [15:0] _U430_out;
wire [15:0] _U431_in;
wire [15:0] _U431_out;
wire [15:0] _U433_in;
wire _U433_clk;
wire [15:0] _U433_out;
wire [15:0] _U434_in;
wire _U434_clk;
wire [15:0] _U434_out;
wire [15:0] _U435_in;
wire _U435_clk;
wire [15:0] _U435_out;
assign _U235_in = _U246_out;
_U235_pt__U236 _U235 (
    .in(_U235_in),
    .out(_U235_out)
);
assign _U237_in = 16'(_U382_out * _U385_out);
assign _U237_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U237 (
    .in(_U237_in),
    .clk(_U237_clk),
    .out(_U237_out)
);
assign _U238_in = _U237_out;
assign _U238_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U238 (
    .in(_U238_in),
    .clk(_U238_clk),
    .out(_U238_out)
);
assign _U239_in = _U238_out;
assign _U239_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U239 (
    .in(_U239_in),
    .clk(_U239_clk),
    .out(_U239_out)
);
assign _U240_in = _U239_out;
assign _U240_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U240 (
    .in(_U240_in),
    .clk(_U240_clk),
    .out(_U240_out)
);
assign _U241_in = _U240_out;
assign _U241_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U241 (
    .in(_U241_in),
    .clk(_U241_clk),
    .out(_U241_out)
);
assign _U242_in = _U241_out;
assign _U242_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U242 (
    .in(_U242_in),
    .clk(_U242_clk),
    .out(_U242_out)
);
assign _U243_in = _U242_out;
assign _U243_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U243 (
    .in(_U243_in),
    .clk(_U243_clk),
    .out(_U243_out)
);
assign _U244_in = _U243_out;
assign _U244_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U244 (
    .in(_U244_in),
    .clk(_U244_clk),
    .out(_U244_out)
);
assign _U245_in = _U244_out;
assign _U245_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U245 (
    .in(_U245_in),
    .clk(_U245_clk),
    .out(_U245_out)
);
assign _U246_in = _U245_out;
assign _U246_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U246 (
    .in(_U246_in),
    .clk(_U246_clk),
    .out(_U246_out)
);
assign _U247_in = _U253_out;
_U247_pt__U248 _U247 (
    .in(_U247_in),
    .out(_U247_out)
);
assign _U249_in = 16'(_U364_out * _U373_out);
assign _U249_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U249 (
    .in(_U249_in),
    .clk(_U249_clk),
    .out(_U249_out)
);
assign _U250_in = _U249_out;
assign _U250_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U250 (
    .in(_U250_in),
    .clk(_U250_clk),
    .out(_U250_out)
);
assign _U251_in = _U250_out;
assign _U251_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U251 (
    .in(_U251_in),
    .clk(_U251_clk),
    .out(_U251_out)
);
assign _U252_in = _U251_out;
assign _U252_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U252 (
    .in(_U252_in),
    .clk(_U252_clk),
    .out(_U252_out)
);
assign _U253_in = _U252_out;
assign _U253_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U253 (
    .in(_U253_in),
    .clk(_U253_clk),
    .out(_U253_out)
);
assign _U254_in = _U262_out;
_U254_pt__U255 _U254 (
    .in(_U254_in),
    .out(_U254_out)
);
assign _U256_in = 16'(_U348_out * _U356_out);
assign _U256_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U256 (
    .in(_U256_in),
    .clk(_U256_clk),
    .out(_U256_out)
);
assign _U257_in = _U256_out;
assign _U257_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U257 (
    .in(_U257_in),
    .clk(_U257_clk),
    .out(_U257_out)
);
assign _U258_in = _U257_out;
assign _U258_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U258 (
    .in(_U258_in),
    .clk(_U258_clk),
    .out(_U258_out)
);
assign _U259_in = _U258_out;
assign _U259_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U259 (
    .in(_U259_in),
    .clk(_U259_clk),
    .out(_U259_out)
);
assign _U260_in = _U259_out;
assign _U260_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U260 (
    .in(_U260_in),
    .clk(_U260_clk),
    .out(_U260_out)
);
assign _U261_in = _U260_out;
assign _U261_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U261 (
    .in(_U261_in),
    .clk(_U261_clk),
    .out(_U261_out)
);
assign _U262_in = _U261_out;
assign _U262_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U262 (
    .in(_U262_in),
    .clk(_U262_clk),
    .out(_U262_out)
);
assign _U263_in = _U265_out;
_U263_pt__U264 _U263 (
    .in(_U263_in),
    .out(_U263_out)
);
assign _U265_in = 16'(_U235_out + _U296_out);
assign _U265_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U265 (
    .in(_U265_in),
    .clk(_U265_clk),
    .out(_U265_out)
);
assign _U266_in = 16'(_U302_out + _U316_out);
_U266_pt__U267 _U266 (
    .in(_U266_in),
    .out(out_conv_stencil)
);
assign _U268_in = _U275_out;
_U268_pt__U269 _U268 (
    .in(_U268_in),
    .out(_U268_out)
);
assign _U270_in = 16'(_U414_out * _U418_out);
assign _U270_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U270 (
    .in(_U270_in),
    .clk(_U270_clk),
    .out(_U270_out)
);
assign _U271_in = _U270_out;
assign _U271_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U271 (
    .in(_U271_in),
    .clk(_U271_clk),
    .out(_U271_out)
);
assign _U272_in = _U271_out;
assign _U272_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U272 (
    .in(_U272_in),
    .clk(_U272_clk),
    .out(_U272_out)
);
assign _U273_in = _U272_out;
assign _U273_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U273 (
    .in(_U273_in),
    .clk(_U273_clk),
    .out(_U273_out)
);
assign _U274_in = _U273_out;
assign _U274_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U274 (
    .in(_U274_in),
    .clk(_U274_clk),
    .out(_U274_out)
);
assign _U275_in = _U274_out;
assign _U275_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U275 (
    .in(_U275_in),
    .clk(_U275_clk),
    .out(_U275_out)
);
assign _U276_in = _U281_out;
_U276_pt__U277 _U276 (
    .in(_U276_in),
    .out(_U276_out)
);
assign _U278_in = 16'(_U400_out * _U407_out);
assign _U278_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U278 (
    .in(_U278_in),
    .clk(_U278_clk),
    .out(_U278_out)
);
assign _U279_in = _U278_out;
assign _U279_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U279 (
    .in(_U279_in),
    .clk(_U279_clk),
    .out(_U279_out)
);
assign _U280_in = _U279_out;
assign _U280_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U280 (
    .in(_U280_in),
    .clk(_U280_clk),
    .out(_U280_out)
);
assign _U281_in = _U280_out;
assign _U281_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U281 (
    .in(_U281_in),
    .clk(_U281_clk),
    .out(_U281_out)
);
assign _U282_in = _U289_out;
_U282_pt__U283 _U282 (
    .in(_U282_in),
    .out(_U282_out)
);
assign _U284_in = 16'(_U388_out * _U394_out);
assign _U284_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U284 (
    .in(_U284_in),
    .clk(_U284_clk),
    .out(_U284_out)
);
assign _U285_in = _U284_out;
assign _U285_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U285 (
    .in(_U285_in),
    .clk(_U285_clk),
    .out(_U285_out)
);
assign _U286_in = _U285_out;
assign _U286_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U286 (
    .in(_U286_in),
    .clk(_U286_clk),
    .out(_U286_out)
);
assign _U287_in = _U286_out;
assign _U287_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U287 (
    .in(_U287_in),
    .clk(_U287_clk),
    .out(_U287_out)
);
assign _U288_in = _U287_out;
assign _U288_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U288 (
    .in(_U288_in),
    .clk(_U288_clk),
    .out(_U288_out)
);
assign _U289_in = _U288_out;
assign _U289_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U289 (
    .in(_U289_in),
    .clk(_U289_clk),
    .out(_U289_out)
);
assign _U290_in = _U292_out;
_U290_pt__U291 _U290 (
    .in(_U290_in),
    .out(_U290_out)
);
assign _U292_in = 16'(_U247_out + _U263_out);
assign _U292_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U292 (
    .in(_U292_in),
    .clk(_U292_clk),
    .out(_U292_out)
);
assign _U293_in = _U295_out;
_U293_pt__U294 _U293 (
    .in(_U293_in),
    .out(_U293_out)
);
assign _U295_in = 16'(_U254_out + _U290_out);
assign _U295_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U295 (
    .in(_U295_in),
    .clk(_U295_clk),
    .out(_U295_out)
);
assign _U296_in = _U298_out;
_U296_pt__U297 _U296 (
    .in(_U296_in),
    .out(_U296_out)
);
assign _U298_in = 16'(_U282_out + _U319_out);
assign _U298_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U298 (
    .in(_U298_in),
    .clk(_U298_clk),
    .out(_U298_out)
);
assign _U299_in = _U301_out;
_U299_pt__U300 _U299 (
    .in(_U299_in),
    .out(_U299_out)
);
assign _U301_in = 16'(_U268_out + _U322_out);
assign _U301_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U301 (
    .in(_U301_in),
    .clk(_U301_clk),
    .out(_U301_out)
);
assign _U302_in = _U315_out;
_U302_pt__U303 _U302 (
    .in(_U302_in),
    .out(_U302_out)
);
assign _U304_in = 16'(_U426_out * _U431_out);
assign _U304_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U304 (
    .in(_U304_in),
    .clk(_U304_clk),
    .out(_U304_out)
);
assign _U305_in = _U304_out;
assign _U305_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U305 (
    .in(_U305_in),
    .clk(_U305_clk),
    .out(_U305_out)
);
assign _U306_in = _U305_out;
assign _U306_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U306 (
    .in(_U306_in),
    .clk(_U306_clk),
    .out(_U306_out)
);
assign _U307_in = _U306_out;
assign _U307_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U307 (
    .in(_U307_in),
    .clk(_U307_clk),
    .out(_U307_out)
);
assign _U308_in = _U307_out;
assign _U308_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U308 (
    .in(_U308_in),
    .clk(_U308_clk),
    .out(_U308_out)
);
assign _U309_in = _U308_out;
assign _U309_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U309 (
    .in(_U309_in),
    .clk(_U309_clk),
    .out(_U309_out)
);
assign _U310_in = _U309_out;
assign _U310_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U310 (
    .in(_U310_in),
    .clk(_U310_clk),
    .out(_U310_out)
);
assign _U311_in = _U310_out;
assign _U311_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U311 (
    .in(_U311_in),
    .clk(_U311_clk),
    .out(_U311_out)
);
assign _U312_in = _U311_out;
assign _U312_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U312 (
    .in(_U312_in),
    .clk(_U312_clk),
    .out(_U312_out)
);
assign _U313_in = _U312_out;
assign _U313_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U313 (
    .in(_U313_in),
    .clk(_U313_clk),
    .out(_U313_out)
);
assign _U314_in = _U313_out;
assign _U314_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U314 (
    .in(_U314_in),
    .clk(_U314_clk),
    .out(_U314_out)
);
assign _U315_in = _U314_out;
assign _U315_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U315 (
    .in(_U315_in),
    .clk(_U315_clk),
    .out(_U315_out)
);
assign _U316_in = _U318_out;
_U316_pt__U317 _U316 (
    .in(_U316_in),
    .out(_U316_out)
);
assign _U318_in = 16'(_U332_out + _U293_out);
assign _U318_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U318 (
    .in(_U318_in),
    .clk(_U318_clk),
    .out(_U318_out)
);
assign _U319_in = _U321_out;
_U319_pt__U320 _U319 (
    .in(_U319_in),
    .out(_U319_out)
);
assign _U321_in = 16'(_U276_out + _U299_out);
assign _U321_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U321 (
    .in(_U321_in),
    .clk(_U321_clk),
    .out(_U321_out)
);
assign _U322_in = _U331_out;
_U322_pt__U323 _U322 (
    .in(_U322_in),
    .out(_U322_out)
);
assign _U324_in = 16'(_U422_out * _U424_out);
assign _U324_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U324 (
    .in(_U324_in),
    .clk(_U324_clk),
    .out(_U324_out)
);
assign _U325_in = _U324_out;
assign _U325_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U325 (
    .in(_U325_in),
    .clk(_U325_clk),
    .out(_U325_out)
);
assign _U326_in = _U325_out;
assign _U326_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U326 (
    .in(_U326_in),
    .clk(_U326_clk),
    .out(_U326_out)
);
assign _U327_in = _U326_out;
assign _U327_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U327 (
    .in(_U327_in),
    .clk(_U327_clk),
    .out(_U327_out)
);
assign _U328_in = _U327_out;
assign _U328_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U328 (
    .in(_U328_in),
    .clk(_U328_clk),
    .out(_U328_out)
);
assign _U329_in = _U328_out;
assign _U329_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U329 (
    .in(_U329_in),
    .clk(_U329_clk),
    .out(_U329_out)
);
assign _U330_in = _U329_out;
assign _U330_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U330 (
    .in(_U330_in),
    .clk(_U330_clk),
    .out(_U330_out)
);
assign _U331_in = _U330_out;
assign _U331_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U331 (
    .in(_U331_in),
    .clk(_U331_clk),
    .out(_U331_out)
);
assign _U332_in = _U347_out;
_U332_pt__U333 _U332 (
    .in(_U332_in),
    .out(_U332_out)
);
assign _U334_in = in0_conv_stencil[0];
assign _U334_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U334 (
    .in(_U334_in),
    .clk(_U334_clk),
    .out(_U334_out)
);
assign _U335_in = _U334_out;
assign _U335_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U335 (
    .in(_U335_in),
    .clk(_U335_clk),
    .out(_U335_out)
);
assign _U336_in = _U335_out;
assign _U336_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U336 (
    .in(_U336_in),
    .clk(_U336_clk),
    .out(_U336_out)
);
assign _U337_in = _U336_out;
assign _U337_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U337 (
    .in(_U337_in),
    .clk(_U337_clk),
    .out(_U337_out)
);
assign _U338_in = _U337_out;
assign _U338_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U338 (
    .in(_U338_in),
    .clk(_U338_clk),
    .out(_U338_out)
);
assign _U339_in = _U338_out;
assign _U339_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U339 (
    .in(_U339_in),
    .clk(_U339_clk),
    .out(_U339_out)
);
assign _U340_in = _U339_out;
assign _U340_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U340 (
    .in(_U340_in),
    .clk(_U340_clk),
    .out(_U340_out)
);
assign _U341_in = _U340_out;
assign _U341_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U341 (
    .in(_U341_in),
    .clk(_U341_clk),
    .out(_U341_out)
);
assign _U342_in = _U341_out;
assign _U342_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U342 (
    .in(_U342_in),
    .clk(_U342_clk),
    .out(_U342_out)
);
assign _U343_in = _U342_out;
assign _U343_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U343 (
    .in(_U343_in),
    .clk(_U343_clk),
    .out(_U343_out)
);
assign _U344_in = _U343_out;
assign _U344_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U344 (
    .in(_U344_in),
    .clk(_U344_clk),
    .out(_U344_out)
);
assign _U345_in = _U344_out;
assign _U345_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U345 (
    .in(_U345_in),
    .clk(_U345_clk),
    .out(_U345_out)
);
assign _U346_in = _U345_out;
assign _U346_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U346 (
    .in(_U346_in),
    .clk(_U346_clk),
    .out(_U346_out)
);
assign _U347_in = _U346_out;
assign _U347_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U347 (
    .in(_U347_in),
    .clk(_U347_clk),
    .out(_U347_out)
);
assign _U348_in = _U355_out;
_U348_pt__U349 _U348 (
    .in(_U348_in),
    .out(_U348_out)
);
assign _U350_in = in2_hw_kernel_global_wrapper_stencil[0];
assign _U350_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U350 (
    .in(_U350_in),
    .clk(_U350_clk),
    .out(_U350_out)
);
assign _U351_in = _U350_out;
assign _U351_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U351 (
    .in(_U351_in),
    .clk(_U351_clk),
    .out(_U351_out)
);
assign _U352_in = _U351_out;
assign _U352_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U352 (
    .in(_U352_in),
    .clk(_U352_clk),
    .out(_U352_out)
);
assign _U353_in = _U352_out;
assign _U353_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U353 (
    .in(_U353_in),
    .clk(_U353_clk),
    .out(_U353_out)
);
assign _U354_in = _U353_out;
assign _U354_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U354 (
    .in(_U354_in),
    .clk(_U354_clk),
    .out(_U354_out)
);
assign _U355_in = _U354_out;
assign _U355_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U355 (
    .in(_U355_in),
    .clk(_U355_clk),
    .out(_U355_out)
);
assign _U356_in = _U363_out;
_U356_pt__U357 _U356 (
    .in(_U356_in),
    .out(_U356_out)
);
assign _U358_in = in1_hw_input_global_wrapper_stencil[0];
assign _U358_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U358 (
    .in(_U358_in),
    .clk(_U358_clk),
    .out(_U358_out)
);
assign _U359_in = _U358_out;
assign _U359_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U359 (
    .in(_U359_in),
    .clk(_U359_clk),
    .out(_U359_out)
);
assign _U360_in = _U359_out;
assign _U360_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U360 (
    .in(_U360_in),
    .clk(_U360_clk),
    .out(_U360_out)
);
assign _U361_in = _U360_out;
assign _U361_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U361 (
    .in(_U361_in),
    .clk(_U361_clk),
    .out(_U361_out)
);
assign _U362_in = _U361_out;
assign _U362_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U362 (
    .in(_U362_in),
    .clk(_U362_clk),
    .out(_U362_out)
);
assign _U363_in = _U362_out;
assign _U363_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U363 (
    .in(_U363_in),
    .clk(_U363_clk),
    .out(_U363_out)
);
assign _U364_in = _U372_out;
_U364_pt__U365 _U364 (
    .in(_U364_in),
    .out(_U364_out)
);
assign _U366_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U366_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U366 (
    .in(_U366_in),
    .clk(_U366_clk),
    .out(_U366_out)
);
assign _U367_in = _U366_out;
assign _U367_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U367 (
    .in(_U367_in),
    .clk(_U367_clk),
    .out(_U367_out)
);
assign _U368_in = _U367_out;
assign _U368_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U368 (
    .in(_U368_in),
    .clk(_U368_clk),
    .out(_U368_out)
);
assign _U369_in = _U368_out;
assign _U369_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U369 (
    .in(_U369_in),
    .clk(_U369_clk),
    .out(_U369_out)
);
assign _U370_in = _U369_out;
assign _U370_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U370 (
    .in(_U370_in),
    .clk(_U370_clk),
    .out(_U370_out)
);
assign _U371_in = _U370_out;
assign _U371_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U371 (
    .in(_U371_in),
    .clk(_U371_clk),
    .out(_U371_out)
);
assign _U372_in = _U371_out;
assign _U372_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U372 (
    .in(_U372_in),
    .clk(_U372_clk),
    .out(_U372_out)
);
assign _U373_in = _U381_out;
_U373_pt__U374 _U373 (
    .in(_U373_in),
    .out(_U373_out)
);
assign _U375_in = in1_hw_input_global_wrapper_stencil[1];
assign _U375_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U375 (
    .in(_U375_in),
    .clk(_U375_clk),
    .out(_U375_out)
);
assign _U376_in = _U375_out;
assign _U376_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U376 (
    .in(_U376_in),
    .clk(_U376_clk),
    .out(_U376_out)
);
assign _U377_in = _U376_out;
assign _U377_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U377 (
    .in(_U377_in),
    .clk(_U377_clk),
    .out(_U377_out)
);
assign _U378_in = _U377_out;
assign _U378_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U378 (
    .in(_U378_in),
    .clk(_U378_clk),
    .out(_U378_out)
);
assign _U379_in = _U378_out;
assign _U379_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U379 (
    .in(_U379_in),
    .clk(_U379_clk),
    .out(_U379_out)
);
assign _U380_in = _U379_out;
assign _U380_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U380 (
    .in(_U380_in),
    .clk(_U380_clk),
    .out(_U380_out)
);
assign _U381_in = _U380_out;
assign _U381_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U381 (
    .in(_U381_in),
    .clk(_U381_clk),
    .out(_U381_out)
);
assign _U382_in = _U384_out;
_U382_pt__U383 _U382 (
    .in(_U382_in),
    .out(_U382_out)
);
assign _U384_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U384_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U384 (
    .in(_U384_in),
    .clk(_U384_clk),
    .out(_U384_out)
);
assign _U385_in = _U387_out;
_U385_pt__U386 _U385 (
    .in(_U385_in),
    .out(_U385_out)
);
assign _U387_in = in1_hw_input_global_wrapper_stencil[2];
assign _U387_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U387 (
    .in(_U387_in),
    .clk(_U387_clk),
    .out(_U387_out)
);
assign _U388_in = _U393_out;
_U388_pt__U389 _U388 (
    .in(_U388_in),
    .out(_U388_out)
);
assign _U390_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U390_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U390 (
    .in(_U390_in),
    .clk(_U390_clk),
    .out(_U390_out)
);
assign _U391_in = _U390_out;
assign _U391_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U391 (
    .in(_U391_in),
    .clk(_U391_clk),
    .out(_U391_out)
);
assign _U392_in = _U391_out;
assign _U392_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U392 (
    .in(_U392_in),
    .clk(_U392_clk),
    .out(_U392_out)
);
assign _U393_in = _U392_out;
assign _U393_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U393 (
    .in(_U393_in),
    .clk(_U393_clk),
    .out(_U393_out)
);
assign _U394_in = _U399_out;
_U394_pt__U395 _U394 (
    .in(_U394_in),
    .out(_U394_out)
);
assign _U396_in = in1_hw_input_global_wrapper_stencil[3];
assign _U396_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U396 (
    .in(_U396_in),
    .clk(_U396_clk),
    .out(_U396_out)
);
assign _U397_in = _U396_out;
assign _U397_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U397 (
    .in(_U397_in),
    .clk(_U397_clk),
    .out(_U397_out)
);
assign _U398_in = _U397_out;
assign _U398_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U398 (
    .in(_U398_in),
    .clk(_U398_clk),
    .out(_U398_out)
);
assign _U399_in = _U398_out;
assign _U399_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U399 (
    .in(_U399_in),
    .clk(_U399_clk),
    .out(_U399_out)
);
assign _U400_in = _U406_out;
_U400_pt__U401 _U400 (
    .in(_U400_in),
    .out(_U400_out)
);
assign _U402_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U402_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U402 (
    .in(_U402_in),
    .clk(_U402_clk),
    .out(_U402_out)
);
assign _U403_in = _U402_out;
assign _U403_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U403 (
    .in(_U403_in),
    .clk(_U403_clk),
    .out(_U403_out)
);
assign _U404_in = _U403_out;
assign _U404_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U404 (
    .in(_U404_in),
    .clk(_U404_clk),
    .out(_U404_out)
);
assign _U405_in = _U404_out;
assign _U405_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U405 (
    .in(_U405_in),
    .clk(_U405_clk),
    .out(_U405_out)
);
assign _U406_in = _U405_out;
assign _U406_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U406 (
    .in(_U406_in),
    .clk(_U406_clk),
    .out(_U406_out)
);
assign _U407_in = _U413_out;
_U407_pt__U408 _U407 (
    .in(_U407_in),
    .out(_U407_out)
);
assign _U409_in = in1_hw_input_global_wrapper_stencil[4];
assign _U409_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U409 (
    .in(_U409_in),
    .clk(_U409_clk),
    .out(_U409_out)
);
assign _U410_in = _U409_out;
assign _U410_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U410 (
    .in(_U410_in),
    .clk(_U410_clk),
    .out(_U410_out)
);
assign _U411_in = _U410_out;
assign _U411_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U411 (
    .in(_U411_in),
    .clk(_U411_clk),
    .out(_U411_out)
);
assign _U412_in = _U411_out;
assign _U412_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U412 (
    .in(_U412_in),
    .clk(_U412_clk),
    .out(_U412_out)
);
assign _U413_in = _U412_out;
assign _U413_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U413 (
    .in(_U413_in),
    .clk(_U413_clk),
    .out(_U413_out)
);
assign _U414_in = _U417_out;
_U414_pt__U415 _U414 (
    .in(_U414_in),
    .out(_U414_out)
);
assign _U416_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U416_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U416 (
    .in(_U416_in),
    .clk(_U416_clk),
    .out(_U416_out)
);
assign _U417_in = _U416_out;
assign _U417_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U417 (
    .in(_U417_in),
    .clk(_U417_clk),
    .out(_U417_out)
);
assign _U418_in = _U421_out;
_U418_pt__U419 _U418 (
    .in(_U418_in),
    .out(_U418_out)
);
assign _U420_in = in1_hw_input_global_wrapper_stencil[5];
assign _U420_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U420 (
    .in(_U420_in),
    .clk(_U420_clk),
    .out(_U420_out)
);
assign _U421_in = _U420_out;
assign _U421_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U421 (
    .in(_U421_in),
    .clk(_U421_clk),
    .out(_U421_out)
);
assign _U422_in = in2_hw_kernel_global_wrapper_stencil[6];
_U422_pt__U423 _U422 (
    .in(_U422_in),
    .out(_U422_out)
);
assign _U424_in = in1_hw_input_global_wrapper_stencil[6];
_U424_pt__U425 _U424 (
    .in(_U424_in),
    .out(_U424_out)
);
assign _U426_in = _U430_out;
_U426_pt__U427 _U426 (
    .in(_U426_in),
    .out(_U426_out)
);
assign _U428_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U428_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U428 (
    .in(_U428_in),
    .clk(_U428_clk),
    .out(_U428_out)
);
assign _U429_in = _U428_out;
assign _U429_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U429 (
    .in(_U429_in),
    .clk(_U429_clk),
    .out(_U429_out)
);
assign _U430_in = _U429_out;
assign _U430_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U430 (
    .in(_U430_in),
    .clk(_U430_clk),
    .out(_U430_out)
);
assign _U431_in = _U435_out;
_U431_pt__U432 _U431 (
    .in(_U431_in),
    .out(_U431_out)
);
assign _U433_in = in1_hw_input_global_wrapper_stencil[7];
assign _U433_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U433 (
    .in(_U433_in),
    .clk(_U433_clk),
    .out(_U433_out)
);
assign _U434_in = _U433_out;
assign _U434_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U434 (
    .in(_U434_in),
    .clk(_U434_clk),
    .out(_U434_out)
);
assign _U435_in = _U434_out;
assign _U435_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U435 (
    .in(_U435_in),
    .clk(_U435_clk),
    .out(_U435_out)
);
endmodule

module cu_op_hcompute_conv_stencil_9 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_9_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_9_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_9_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[0];
hcompute_conv_stencil_9_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_9_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U233_pt__U234 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U231_pt__U232 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U22_pt__U23 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_2_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U22_in;
assign _U22_in = 16'h0000;
_U22_pt__U23 _U22 (
    .in(_U22_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_2 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_2_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U215_pt__U216 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U212_pt__U213 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U20_pt__U21 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_1_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U20_in;
assign _U20_in = 16'h0000;
_U20_pt__U21 _U20 (
    .in(_U20_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_1 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_1_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U208_pt__U209 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U205_pt__U206 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U199_pt__U200 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U196_pt__U197 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U18_pt__U19 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U18_in;
assign _U18_in = 16'h0000;
_U18_pt__U19 _U18 (
    .in(_U18_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U188_pt__U189 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U185_pt__U186 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U175_pt__U176 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U172_pt__U173 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U16_pt__U17 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_kernel_global_wrapper_stencil_pipelined (
    output [15:0] out_hw_kernel_global_wrapper_stencil,
    input [15:0] in0_hw_kernel_stencil [0:0]
);
wire [15:0] _U16_in;
assign _U16_in = in0_hw_kernel_stencil[0];
_U16_pt__U17 _U16 (
    .in(_U16_in),
    .out(out_hw_kernel_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_kernel_global_wrapper_stencil (
    input clk,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_kernel_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_kernel_stencil [0:0];
assign inner_compute_in0_hw_kernel_stencil[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
hcompute_hw_kernel_global_wrapper_stencil_pipelined inner_compute (
    .out_hw_kernel_global_wrapper_stencil(inner_compute_out_hw_kernel_global_wrapper_stencil),
    .in0_hw_kernel_stencil(inner_compute_in0_hw_kernel_stencil)
);
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = inner_compute_out_hw_kernel_global_wrapper_stencil;
endmodule

module _U1656_pt__U1657 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_7_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
wire [15:0] _U1656_in;
assign _U1656_in = in0_conv_stencil[0];
_U1656_pt__U1657 _U1656 (
    .in(_U1656_in),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil_7 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_7_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_7_read[0];
hcompute_hw_output_stencil_7_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1654_pt__U1655 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_6_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
wire [15:0] _U1654_in;
assign _U1654_in = in0_conv_stencil[0];
_U1654_pt__U1655 _U1654 (
    .in(_U1654_in),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil_6 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_6_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_6_read[0];
hcompute_hw_output_stencil_6_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1652_pt__U1653 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_5_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
wire [15:0] _U1652_in;
assign _U1652_in = in0_conv_stencil[0];
_U1652_pt__U1653 _U1652 (
    .in(_U1652_in),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil_5 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_5_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_5_read[0];
hcompute_hw_output_stencil_5_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1650_pt__U1651 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_4_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
wire [15:0] _U1650_in;
assign _U1650_in = in0_conv_stencil[0];
_U1650_pt__U1651 _U1650 (
    .in(_U1650_in),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil_4 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_4_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_4_read[0];
hcompute_hw_output_stencil_4_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1648_pt__U1649 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_3_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
wire [15:0] _U1648_in;
assign _U1648_in = in0_conv_stencil[0];
_U1648_pt__U1649 _U1648 (
    .in(_U1648_in),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil_3 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_3_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_3_read[0];
hcompute_hw_output_stencil_3_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1646_pt__U1647 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_2_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
wire [15:0] _U1646_in;
assign _U1646_in = in0_conv_stencil[0];
_U1646_pt__U1647 _U1646 (
    .in(_U1646_in),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil_2 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_2_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_2_read[0];
hcompute_hw_output_stencil_2_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1644_pt__U1645 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_1_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
wire [15:0] _U1644_in;
assign _U1644_in = in0_conv_stencil[0];
_U1644_pt__U1645 _U1644 (
    .in(_U1644_in),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil_1 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_1_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_1_read[0];
hcompute_hw_output_stencil_1_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1642_pt__U1643 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
wire [15:0] _U1642_in;
assign _U1642_in = in0_conv_stencil[0];
_U1642_pt__U1643 _U1642 (
    .in(_U1642_in),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0],
    output [15:0] hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
hcompute_hw_output_stencil_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U1640_pt__U1641 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1624_pt__U1625 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1621_pt__U1622 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1617_pt__U1618 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1614_pt__U1615 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U160_pt__U161 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1608_pt__U1609 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1605_pt__U1606 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1597_pt__U1598 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1590_pt__U1591 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1584_pt__U1585 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U157_pt__U158 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1578_pt__U1579 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1573_pt__U1574 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1568_pt__U1569 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1564_pt__U1565 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1560_pt__U1561 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1557_pt__U1558 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1554_pt__U1555 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1552_pt__U1553 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1549_pt__U1550 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1539_pt__U1540 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1536_pt__U1537 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1524_pt__U1525 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1521_pt__U1522 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1518_pt__U1519 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1504_pt__U1505 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1502_pt__U1503 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U14_pt__U15 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_7_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
wire [15:0] _U14_in;
assign _U14_in = in0_hw_input_stencil[0];
_U14_pt__U15 _U14 (
    .in(_U14_in),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil_7 (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read[0];
hcompute_hw_input_global_wrapper_stencil_7_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U1499_pt__U1500 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1490_pt__U1491 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1481_pt__U1482 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1473_pt__U1474 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1465_pt__U1466 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1458_pt__U1459 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1441_pt__U1442 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_15_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U1441_in;
wire [15:0] _U1441_out;
wire [15:0] _U1443_in;
wire _U1443_clk;
wire [15:0] _U1443_out;
wire [15:0] _U1444_in;
wire _U1444_clk;
wire [15:0] _U1444_out;
wire [15:0] _U1445_in;
wire _U1445_clk;
wire [15:0] _U1445_out;
wire [15:0] _U1446_in;
wire _U1446_clk;
wire [15:0] _U1446_out;
wire [15:0] _U1447_in;
wire _U1447_clk;
wire [15:0] _U1447_out;
wire [15:0] _U1448_in;
wire _U1448_clk;
wire [15:0] _U1448_out;
wire [15:0] _U1449_in;
wire _U1449_clk;
wire [15:0] _U1449_out;
wire [15:0] _U1450_in;
wire _U1450_clk;
wire [15:0] _U1450_out;
wire [15:0] _U1451_in;
wire _U1451_clk;
wire [15:0] _U1451_out;
wire [15:0] _U1452_in;
wire _U1452_clk;
wire [15:0] _U1452_out;
wire [15:0] _U1453_in;
wire _U1453_clk;
wire [15:0] _U1453_out;
wire [15:0] _U1454_in;
wire _U1454_clk;
wire [15:0] _U1454_out;
wire [15:0] _U1455_in;
wire _U1455_clk;
wire [15:0] _U1455_out;
wire [15:0] _U1456_in;
wire _U1456_clk;
wire [15:0] _U1456_out;
wire [15:0] _U1457_in;
wire _U1457_clk;
wire [15:0] _U1457_out;
wire [15:0] _U1458_in;
wire [15:0] _U1458_out;
wire [15:0] _U1460_in;
wire _U1460_clk;
wire [15:0] _U1460_out;
wire [15:0] _U1461_in;
wire _U1461_clk;
wire [15:0] _U1461_out;
wire [15:0] _U1462_in;
wire _U1462_clk;
wire [15:0] _U1462_out;
wire [15:0] _U1463_in;
wire _U1463_clk;
wire [15:0] _U1463_out;
wire [15:0] _U1464_in;
wire _U1464_clk;
wire [15:0] _U1464_out;
wire [15:0] _U1465_in;
wire [15:0] _U1465_out;
wire [15:0] _U1467_in;
wire _U1467_clk;
wire [15:0] _U1467_out;
wire [15:0] _U1468_in;
wire _U1468_clk;
wire [15:0] _U1468_out;
wire [15:0] _U1469_in;
wire _U1469_clk;
wire [15:0] _U1469_out;
wire [15:0] _U1470_in;
wire _U1470_clk;
wire [15:0] _U1470_out;
wire [15:0] _U1471_in;
wire _U1471_clk;
wire [15:0] _U1471_out;
wire [15:0] _U1472_in;
wire _U1472_clk;
wire [15:0] _U1472_out;
wire [15:0] _U1473_in;
wire [15:0] _U1473_out;
wire [15:0] _U1475_in;
wire _U1475_clk;
wire [15:0] _U1475_out;
wire [15:0] _U1476_in;
wire _U1476_clk;
wire [15:0] _U1476_out;
wire [15:0] _U1477_in;
wire _U1477_clk;
wire [15:0] _U1477_out;
wire [15:0] _U1478_in;
wire _U1478_clk;
wire [15:0] _U1478_out;
wire [15:0] _U1479_in;
wire _U1479_clk;
wire [15:0] _U1479_out;
wire [15:0] _U1480_in;
wire _U1480_clk;
wire [15:0] _U1480_out;
wire [15:0] _U1481_in;
wire [15:0] _U1481_out;
wire [15:0] _U1483_in;
wire _U1483_clk;
wire [15:0] _U1483_out;
wire [15:0] _U1484_in;
wire _U1484_clk;
wire [15:0] _U1484_out;
wire [15:0] _U1485_in;
wire _U1485_clk;
wire [15:0] _U1485_out;
wire [15:0] _U1486_in;
wire _U1486_clk;
wire [15:0] _U1486_out;
wire [15:0] _U1487_in;
wire _U1487_clk;
wire [15:0] _U1487_out;
wire [15:0] _U1488_in;
wire _U1488_clk;
wire [15:0] _U1488_out;
wire [15:0] _U1489_in;
wire _U1489_clk;
wire [15:0] _U1489_out;
wire [15:0] _U1490_in;
wire [15:0] _U1490_out;
wire [15:0] _U1492_in;
wire _U1492_clk;
wire [15:0] _U1492_out;
wire [15:0] _U1493_in;
wire _U1493_clk;
wire [15:0] _U1493_out;
wire [15:0] _U1494_in;
wire _U1494_clk;
wire [15:0] _U1494_out;
wire [15:0] _U1495_in;
wire _U1495_clk;
wire [15:0] _U1495_out;
wire [15:0] _U1496_in;
wire _U1496_clk;
wire [15:0] _U1496_out;
wire [15:0] _U1497_in;
wire _U1497_clk;
wire [15:0] _U1497_out;
wire [15:0] _U1498_in;
wire _U1498_clk;
wire [15:0] _U1498_out;
wire [15:0] _U1499_in;
wire [15:0] _U1499_out;
wire [15:0] _U1501_in;
wire _U1501_clk;
wire [15:0] _U1501_out;
wire [15:0] _U1502_in;
wire [15:0] _U1504_in;
wire [15:0] _U1504_out;
wire [15:0] _U1506_in;
wire _U1506_clk;
wire [15:0] _U1506_out;
wire [15:0] _U1507_in;
wire _U1507_clk;
wire [15:0] _U1507_out;
wire [15:0] _U1508_in;
wire _U1508_clk;
wire [15:0] _U1508_out;
wire [15:0] _U1509_in;
wire _U1509_clk;
wire [15:0] _U1509_out;
wire [15:0] _U1510_in;
wire _U1510_clk;
wire [15:0] _U1510_out;
wire [15:0] _U1511_in;
wire _U1511_clk;
wire [15:0] _U1511_out;
wire [15:0] _U1512_in;
wire _U1512_clk;
wire [15:0] _U1512_out;
wire [15:0] _U1513_in;
wire _U1513_clk;
wire [15:0] _U1513_out;
wire [15:0] _U1514_in;
wire _U1514_clk;
wire [15:0] _U1514_out;
wire [15:0] _U1515_in;
wire _U1515_clk;
wire [15:0] _U1515_out;
wire [15:0] _U1516_in;
wire _U1516_clk;
wire [15:0] _U1516_out;
wire [15:0] _U1517_in;
wire _U1517_clk;
wire [15:0] _U1517_out;
wire [15:0] _U1518_in;
wire [15:0] _U1518_out;
wire [15:0] _U1520_in;
wire _U1520_clk;
wire [15:0] _U1520_out;
wire [15:0] _U1521_in;
wire [15:0] _U1521_out;
wire [15:0] _U1523_in;
wire _U1523_clk;
wire [15:0] _U1523_out;
wire [15:0] _U1524_in;
wire [15:0] _U1524_out;
wire [15:0] _U1526_in;
wire _U1526_clk;
wire [15:0] _U1526_out;
wire [15:0] _U1527_in;
wire _U1527_clk;
wire [15:0] _U1527_out;
wire [15:0] _U1528_in;
wire _U1528_clk;
wire [15:0] _U1528_out;
wire [15:0] _U1529_in;
wire _U1529_clk;
wire [15:0] _U1529_out;
wire [15:0] _U1530_in;
wire _U1530_clk;
wire [15:0] _U1530_out;
wire [15:0] _U1531_in;
wire _U1531_clk;
wire [15:0] _U1531_out;
wire [15:0] _U1532_in;
wire _U1532_clk;
wire [15:0] _U1532_out;
wire [15:0] _U1533_in;
wire _U1533_clk;
wire [15:0] _U1533_out;
wire [15:0] _U1534_in;
wire _U1534_clk;
wire [15:0] _U1534_out;
wire [15:0] _U1535_in;
wire _U1535_clk;
wire [15:0] _U1535_out;
wire [15:0] _U1536_in;
wire [15:0] _U1536_out;
wire [15:0] _U1538_in;
wire _U1538_clk;
wire [15:0] _U1538_out;
wire [15:0] _U1539_in;
wire [15:0] _U1539_out;
wire [15:0] _U1541_in;
wire _U1541_clk;
wire [15:0] _U1541_out;
wire [15:0] _U1542_in;
wire _U1542_clk;
wire [15:0] _U1542_out;
wire [15:0] _U1543_in;
wire _U1543_clk;
wire [15:0] _U1543_out;
wire [15:0] _U1544_in;
wire _U1544_clk;
wire [15:0] _U1544_out;
wire [15:0] _U1545_in;
wire _U1545_clk;
wire [15:0] _U1545_out;
wire [15:0] _U1546_in;
wire _U1546_clk;
wire [15:0] _U1546_out;
wire [15:0] _U1547_in;
wire _U1547_clk;
wire [15:0] _U1547_out;
wire [15:0] _U1548_in;
wire _U1548_clk;
wire [15:0] _U1548_out;
wire [15:0] _U1549_in;
wire [15:0] _U1549_out;
wire [15:0] _U1551_in;
wire _U1551_clk;
wire [15:0] _U1551_out;
wire [15:0] _U1552_in;
wire [15:0] _U1552_out;
wire [15:0] _U1554_in;
wire [15:0] _U1554_out;
wire [15:0] _U1556_in;
wire _U1556_clk;
wire [15:0] _U1556_out;
wire [15:0] _U1557_in;
wire [15:0] _U1557_out;
wire [15:0] _U1559_in;
wire _U1559_clk;
wire [15:0] _U1559_out;
wire [15:0] _U1560_in;
wire [15:0] _U1560_out;
wire [15:0] _U1562_in;
wire _U1562_clk;
wire [15:0] _U1562_out;
wire [15:0] _U1563_in;
wire _U1563_clk;
wire [15:0] _U1563_out;
wire [15:0] _U1564_in;
wire [15:0] _U1564_out;
wire [15:0] _U1566_in;
wire _U1566_clk;
wire [15:0] _U1566_out;
wire [15:0] _U1567_in;
wire _U1567_clk;
wire [15:0] _U1567_out;
wire [15:0] _U1568_in;
wire [15:0] _U1568_out;
wire [15:0] _U1570_in;
wire _U1570_clk;
wire [15:0] _U1570_out;
wire [15:0] _U1571_in;
wire _U1571_clk;
wire [15:0] _U1571_out;
wire [15:0] _U1572_in;
wire _U1572_clk;
wire [15:0] _U1572_out;
wire [15:0] _U1573_in;
wire [15:0] _U1573_out;
wire [15:0] _U1575_in;
wire _U1575_clk;
wire [15:0] _U1575_out;
wire [15:0] _U1576_in;
wire _U1576_clk;
wire [15:0] _U1576_out;
wire [15:0] _U1577_in;
wire _U1577_clk;
wire [15:0] _U1577_out;
wire [15:0] _U1578_in;
wire [15:0] _U1578_out;
wire [15:0] _U1580_in;
wire _U1580_clk;
wire [15:0] _U1580_out;
wire [15:0] _U1581_in;
wire _U1581_clk;
wire [15:0] _U1581_out;
wire [15:0] _U1582_in;
wire _U1582_clk;
wire [15:0] _U1582_out;
wire [15:0] _U1583_in;
wire _U1583_clk;
wire [15:0] _U1583_out;
wire [15:0] _U1584_in;
wire [15:0] _U1584_out;
wire [15:0] _U1586_in;
wire _U1586_clk;
wire [15:0] _U1586_out;
wire [15:0] _U1587_in;
wire _U1587_clk;
wire [15:0] _U1587_out;
wire [15:0] _U1588_in;
wire _U1588_clk;
wire [15:0] _U1588_out;
wire [15:0] _U1589_in;
wire _U1589_clk;
wire [15:0] _U1589_out;
wire [15:0] _U1590_in;
wire [15:0] _U1590_out;
wire [15:0] _U1592_in;
wire _U1592_clk;
wire [15:0] _U1592_out;
wire [15:0] _U1593_in;
wire _U1593_clk;
wire [15:0] _U1593_out;
wire [15:0] _U1594_in;
wire _U1594_clk;
wire [15:0] _U1594_out;
wire [15:0] _U1595_in;
wire _U1595_clk;
wire [15:0] _U1595_out;
wire [15:0] _U1596_in;
wire _U1596_clk;
wire [15:0] _U1596_out;
wire [15:0] _U1597_in;
wire [15:0] _U1597_out;
wire [15:0] _U1599_in;
wire _U1599_clk;
wire [15:0] _U1599_out;
wire [15:0] _U1600_in;
wire _U1600_clk;
wire [15:0] _U1600_out;
wire [15:0] _U1601_in;
wire _U1601_clk;
wire [15:0] _U1601_out;
wire [15:0] _U1602_in;
wire _U1602_clk;
wire [15:0] _U1602_out;
wire [15:0] _U1603_in;
wire _U1603_clk;
wire [15:0] _U1603_out;
wire [15:0] _U1604_in;
wire _U1604_clk;
wire [15:0] _U1604_out;
wire [15:0] _U1605_in;
wire [15:0] _U1605_out;
wire [15:0] _U1607_in;
wire _U1607_clk;
wire [15:0] _U1607_out;
wire [15:0] _U1608_in;
wire [15:0] _U1608_out;
wire [15:0] _U1610_in;
wire _U1610_clk;
wire [15:0] _U1610_out;
wire [15:0] _U1611_in;
wire _U1611_clk;
wire [15:0] _U1611_out;
wire [15:0] _U1612_in;
wire _U1612_clk;
wire [15:0] _U1612_out;
wire [15:0] _U1613_in;
wire _U1613_clk;
wire [15:0] _U1613_out;
wire [15:0] _U1614_in;
wire [15:0] _U1614_out;
wire [15:0] _U1616_in;
wire _U1616_clk;
wire [15:0] _U1616_out;
wire [15:0] _U1617_in;
wire [15:0] _U1617_out;
wire [15:0] _U1619_in;
wire _U1619_clk;
wire [15:0] _U1619_out;
wire [15:0] _U1620_in;
wire _U1620_clk;
wire [15:0] _U1620_out;
wire [15:0] _U1621_in;
wire [15:0] _U1621_out;
wire [15:0] _U1623_in;
wire _U1623_clk;
wire [15:0] _U1623_out;
wire [15:0] _U1624_in;
wire [15:0] _U1624_out;
wire [15:0] _U1626_in;
wire _U1626_clk;
wire [15:0] _U1626_out;
wire [15:0] _U1627_in;
wire _U1627_clk;
wire [15:0] _U1627_out;
wire [15:0] _U1628_in;
wire _U1628_clk;
wire [15:0] _U1628_out;
wire [15:0] _U1629_in;
wire _U1629_clk;
wire [15:0] _U1629_out;
wire [15:0] _U1630_in;
wire _U1630_clk;
wire [15:0] _U1630_out;
wire [15:0] _U1631_in;
wire _U1631_clk;
wire [15:0] _U1631_out;
wire [15:0] _U1632_in;
wire _U1632_clk;
wire [15:0] _U1632_out;
wire [15:0] _U1633_in;
wire _U1633_clk;
wire [15:0] _U1633_out;
wire [15:0] _U1634_in;
wire _U1634_clk;
wire [15:0] _U1634_out;
wire [15:0] _U1635_in;
wire _U1635_clk;
wire [15:0] _U1635_out;
wire [15:0] _U1636_in;
wire _U1636_clk;
wire [15:0] _U1636_out;
wire [15:0] _U1637_in;
wire _U1637_clk;
wire [15:0] _U1637_out;
wire [15:0] _U1638_in;
wire _U1638_clk;
wire [15:0] _U1638_out;
wire [15:0] _U1639_in;
wire _U1639_clk;
wire [15:0] _U1639_out;
wire [15:0] _U1640_in;
wire [15:0] _U1640_out;
assign _U1441_in = _U1457_out;
_U1441_pt__U1442 _U1441 (
    .in(_U1441_in),
    .out(_U1441_out)
);
assign _U1443_in = 16'(_U1640_out * _U1552_out);
assign _U1443_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1443 (
    .in(_U1443_in),
    .clk(_U1443_clk),
    .out(_U1443_out)
);
assign _U1444_in = _U1443_out;
assign _U1444_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1444 (
    .in(_U1444_in),
    .clk(_U1444_clk),
    .out(_U1444_out)
);
assign _U1445_in = _U1444_out;
assign _U1445_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1445 (
    .in(_U1445_in),
    .clk(_U1445_clk),
    .out(_U1445_out)
);
assign _U1446_in = _U1445_out;
assign _U1446_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1446 (
    .in(_U1446_in),
    .clk(_U1446_clk),
    .out(_U1446_out)
);
assign _U1447_in = _U1446_out;
assign _U1447_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1447 (
    .in(_U1447_in),
    .clk(_U1447_clk),
    .out(_U1447_out)
);
assign _U1448_in = _U1447_out;
assign _U1448_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1448 (
    .in(_U1448_in),
    .clk(_U1448_clk),
    .out(_U1448_out)
);
assign _U1449_in = _U1448_out;
assign _U1449_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1449 (
    .in(_U1449_in),
    .clk(_U1449_clk),
    .out(_U1449_out)
);
assign _U1450_in = _U1449_out;
assign _U1450_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1450 (
    .in(_U1450_in),
    .clk(_U1450_clk),
    .out(_U1450_out)
);
assign _U1451_in = _U1450_out;
assign _U1451_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1451 (
    .in(_U1451_in),
    .clk(_U1451_clk),
    .out(_U1451_out)
);
assign _U1452_in = _U1451_out;
assign _U1452_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1452 (
    .in(_U1452_in),
    .clk(_U1452_clk),
    .out(_U1452_out)
);
assign _U1453_in = _U1452_out;
assign _U1453_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1453 (
    .in(_U1453_in),
    .clk(_U1453_clk),
    .out(_U1453_out)
);
assign _U1454_in = _U1453_out;
assign _U1454_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1454 (
    .in(_U1454_in),
    .clk(_U1454_clk),
    .out(_U1454_out)
);
assign _U1455_in = _U1454_out;
assign _U1455_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1455 (
    .in(_U1455_in),
    .clk(_U1455_clk),
    .out(_U1455_out)
);
assign _U1456_in = _U1455_out;
assign _U1456_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1456 (
    .in(_U1456_in),
    .clk(_U1456_clk),
    .out(_U1456_out)
);
assign _U1457_in = _U1456_out;
assign _U1457_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1457 (
    .in(_U1457_in),
    .clk(_U1457_clk),
    .out(_U1457_out)
);
assign _U1458_in = _U1464_out;
_U1458_pt__U1459 _U1458 (
    .in(_U1458_in),
    .out(_U1458_out)
);
assign _U1460_in = in1_hw_input_global_wrapper_stencil[5];
assign _U1460_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1460 (
    .in(_U1460_in),
    .clk(_U1460_clk),
    .out(_U1460_out)
);
assign _U1461_in = _U1460_out;
assign _U1461_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1461 (
    .in(_U1461_in),
    .clk(_U1461_clk),
    .out(_U1461_out)
);
assign _U1462_in = _U1461_out;
assign _U1462_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1462 (
    .in(_U1462_in),
    .clk(_U1462_clk),
    .out(_U1462_out)
);
assign _U1463_in = _U1462_out;
assign _U1463_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1463 (
    .in(_U1463_in),
    .clk(_U1463_clk),
    .out(_U1463_out)
);
assign _U1464_in = _U1463_out;
assign _U1464_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1464 (
    .in(_U1464_in),
    .clk(_U1464_clk),
    .out(_U1464_out)
);
assign _U1465_in = _U1472_out;
_U1465_pt__U1466 _U1465 (
    .in(_U1465_in),
    .out(_U1465_out)
);
assign _U1467_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U1467_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1467 (
    .in(_U1467_in),
    .clk(_U1467_clk),
    .out(_U1467_out)
);
assign _U1468_in = _U1467_out;
assign _U1468_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1468 (
    .in(_U1468_in),
    .clk(_U1468_clk),
    .out(_U1468_out)
);
assign _U1469_in = _U1468_out;
assign _U1469_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1469 (
    .in(_U1469_in),
    .clk(_U1469_clk),
    .out(_U1469_out)
);
assign _U1470_in = _U1469_out;
assign _U1470_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1470 (
    .in(_U1470_in),
    .clk(_U1470_clk),
    .out(_U1470_out)
);
assign _U1471_in = _U1470_out;
assign _U1471_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1471 (
    .in(_U1471_in),
    .clk(_U1471_clk),
    .out(_U1471_out)
);
assign _U1472_in = _U1471_out;
assign _U1472_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1472 (
    .in(_U1472_in),
    .clk(_U1472_clk),
    .out(_U1472_out)
);
assign _U1473_in = _U1480_out;
_U1473_pt__U1474 _U1473 (
    .in(_U1473_in),
    .out(_U1473_out)
);
assign _U1475_in = in1_hw_input_global_wrapper_stencil[6];
assign _U1475_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1475 (
    .in(_U1475_in),
    .clk(_U1475_clk),
    .out(_U1475_out)
);
assign _U1476_in = _U1475_out;
assign _U1476_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1476 (
    .in(_U1476_in),
    .clk(_U1476_clk),
    .out(_U1476_out)
);
assign _U1477_in = _U1476_out;
assign _U1477_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1477 (
    .in(_U1477_in),
    .clk(_U1477_clk),
    .out(_U1477_out)
);
assign _U1478_in = _U1477_out;
assign _U1478_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1478 (
    .in(_U1478_in),
    .clk(_U1478_clk),
    .out(_U1478_out)
);
assign _U1479_in = _U1478_out;
assign _U1479_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1479 (
    .in(_U1479_in),
    .clk(_U1479_clk),
    .out(_U1479_out)
);
assign _U1480_in = _U1479_out;
assign _U1480_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1480 (
    .in(_U1480_in),
    .clk(_U1480_clk),
    .out(_U1480_out)
);
assign _U1481_in = _U1489_out;
_U1481_pt__U1482 _U1481 (
    .in(_U1481_in),
    .out(_U1481_out)
);
assign _U1483_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U1483_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1483 (
    .in(_U1483_in),
    .clk(_U1483_clk),
    .out(_U1483_out)
);
assign _U1484_in = _U1483_out;
assign _U1484_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1484 (
    .in(_U1484_in),
    .clk(_U1484_clk),
    .out(_U1484_out)
);
assign _U1485_in = _U1484_out;
assign _U1485_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1485 (
    .in(_U1485_in),
    .clk(_U1485_clk),
    .out(_U1485_out)
);
assign _U1486_in = _U1485_out;
assign _U1486_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1486 (
    .in(_U1486_in),
    .clk(_U1486_clk),
    .out(_U1486_out)
);
assign _U1487_in = _U1486_out;
assign _U1487_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1487 (
    .in(_U1487_in),
    .clk(_U1487_clk),
    .out(_U1487_out)
);
assign _U1488_in = _U1487_out;
assign _U1488_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1488 (
    .in(_U1488_in),
    .clk(_U1488_clk),
    .out(_U1488_out)
);
assign _U1489_in = _U1488_out;
assign _U1489_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1489 (
    .in(_U1489_in),
    .clk(_U1489_clk),
    .out(_U1489_out)
);
assign _U1490_in = _U1498_out;
_U1490_pt__U1491 _U1490 (
    .in(_U1490_in),
    .out(_U1490_out)
);
assign _U1492_in = in1_hw_input_global_wrapper_stencil[7];
assign _U1492_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1492 (
    .in(_U1492_in),
    .clk(_U1492_clk),
    .out(_U1492_out)
);
assign _U1493_in = _U1492_out;
assign _U1493_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1493 (
    .in(_U1493_in),
    .clk(_U1493_clk),
    .out(_U1493_out)
);
assign _U1494_in = _U1493_out;
assign _U1494_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1494 (
    .in(_U1494_in),
    .clk(_U1494_clk),
    .out(_U1494_out)
);
assign _U1495_in = _U1494_out;
assign _U1495_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1495 (
    .in(_U1495_in),
    .clk(_U1495_clk),
    .out(_U1495_out)
);
assign _U1496_in = _U1495_out;
assign _U1496_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1496 (
    .in(_U1496_in),
    .clk(_U1496_clk),
    .out(_U1496_out)
);
assign _U1497_in = _U1496_out;
assign _U1497_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1497 (
    .in(_U1497_in),
    .clk(_U1497_clk),
    .out(_U1497_out)
);
assign _U1498_in = _U1497_out;
assign _U1498_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1498 (
    .in(_U1498_in),
    .clk(_U1498_clk),
    .out(_U1498_out)
);
assign _U1499_in = _U1501_out;
_U1499_pt__U1500 _U1499 (
    .in(_U1499_in),
    .out(_U1499_out)
);
assign _U1501_in = 16'(_U1624_out + _U1521_out);
assign _U1501_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1501 (
    .in(_U1501_in),
    .clk(_U1501_clk),
    .out(_U1501_out)
);
assign _U1502_in = 16'(_U1441_out + _U1499_out);
_U1502_pt__U1503 _U1502 (
    .in(_U1502_in),
    .out(out_conv_stencil)
);
assign _U1504_in = _U1517_out;
_U1504_pt__U1505 _U1504 (
    .in(_U1504_in),
    .out(_U1504_out)
);
assign _U1506_in = 16'(_U1554_out * _U1557_out);
assign _U1506_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1506 (
    .in(_U1506_in),
    .clk(_U1506_clk),
    .out(_U1506_out)
);
assign _U1507_in = _U1506_out;
assign _U1507_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1507 (
    .in(_U1507_in),
    .clk(_U1507_clk),
    .out(_U1507_out)
);
assign _U1508_in = _U1507_out;
assign _U1508_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1508 (
    .in(_U1508_in),
    .clk(_U1508_clk),
    .out(_U1508_out)
);
assign _U1509_in = _U1508_out;
assign _U1509_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1509 (
    .in(_U1509_in),
    .clk(_U1509_clk),
    .out(_U1509_out)
);
assign _U1510_in = _U1509_out;
assign _U1510_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1510 (
    .in(_U1510_in),
    .clk(_U1510_clk),
    .out(_U1510_out)
);
assign _U1511_in = _U1510_out;
assign _U1511_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1511 (
    .in(_U1511_in),
    .clk(_U1511_clk),
    .out(_U1511_out)
);
assign _U1512_in = _U1511_out;
assign _U1512_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1512 (
    .in(_U1512_in),
    .clk(_U1512_clk),
    .out(_U1512_out)
);
assign _U1513_in = _U1512_out;
assign _U1513_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1513 (
    .in(_U1513_in),
    .clk(_U1513_clk),
    .out(_U1513_out)
);
assign _U1514_in = _U1513_out;
assign _U1514_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1514 (
    .in(_U1514_in),
    .clk(_U1514_clk),
    .out(_U1514_out)
);
assign _U1515_in = _U1514_out;
assign _U1515_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1515 (
    .in(_U1515_in),
    .clk(_U1515_clk),
    .out(_U1515_out)
);
assign _U1516_in = _U1515_out;
assign _U1516_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1516 (
    .in(_U1516_in),
    .clk(_U1516_clk),
    .out(_U1516_out)
);
assign _U1517_in = _U1516_out;
assign _U1517_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1517 (
    .in(_U1517_in),
    .clk(_U1517_clk),
    .out(_U1517_out)
);
assign _U1518_in = _U1520_out;
_U1518_pt__U1519 _U1518 (
    .in(_U1518_in),
    .out(_U1518_out)
);
assign _U1520_in = 16'(_U1524_out + _U1536_out);
assign _U1520_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1520 (
    .in(_U1520_in),
    .clk(_U1520_clk),
    .out(_U1520_out)
);
assign _U1521_in = _U1523_out;
_U1521_pt__U1522 _U1521 (
    .in(_U1521_in),
    .out(_U1521_out)
);
assign _U1523_in = 16'(_U1504_out + _U1518_out);
assign _U1523_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1523 (
    .in(_U1523_in),
    .clk(_U1523_clk),
    .out(_U1523_out)
);
assign _U1524_in = _U1535_out;
_U1524_pt__U1525 _U1524 (
    .in(_U1524_in),
    .out(_U1524_out)
);
assign _U1526_in = 16'(_U1560_out * _U1564_out);
assign _U1526_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1526 (
    .in(_U1526_in),
    .clk(_U1526_clk),
    .out(_U1526_out)
);
assign _U1527_in = _U1526_out;
assign _U1527_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1527 (
    .in(_U1527_in),
    .clk(_U1527_clk),
    .out(_U1527_out)
);
assign _U1528_in = _U1527_out;
assign _U1528_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1528 (
    .in(_U1528_in),
    .clk(_U1528_clk),
    .out(_U1528_out)
);
assign _U1529_in = _U1528_out;
assign _U1529_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1529 (
    .in(_U1529_in),
    .clk(_U1529_clk),
    .out(_U1529_out)
);
assign _U1530_in = _U1529_out;
assign _U1530_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1530 (
    .in(_U1530_in),
    .clk(_U1530_clk),
    .out(_U1530_out)
);
assign _U1531_in = _U1530_out;
assign _U1531_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1531 (
    .in(_U1531_in),
    .clk(_U1531_clk),
    .out(_U1531_out)
);
assign _U1532_in = _U1531_out;
assign _U1532_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1532 (
    .in(_U1532_in),
    .clk(_U1532_clk),
    .out(_U1532_out)
);
assign _U1533_in = _U1532_out;
assign _U1533_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1533 (
    .in(_U1533_in),
    .clk(_U1533_clk),
    .out(_U1533_out)
);
assign _U1534_in = _U1533_out;
assign _U1534_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1534 (
    .in(_U1534_in),
    .clk(_U1534_clk),
    .out(_U1534_out)
);
assign _U1535_in = _U1534_out;
assign _U1535_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1535 (
    .in(_U1535_in),
    .clk(_U1535_clk),
    .out(_U1535_out)
);
assign _U1536_in = _U1538_out;
_U1536_pt__U1537 _U1536 (
    .in(_U1536_in),
    .out(_U1536_out)
);
assign _U1538_in = 16'(_U1539_out + _U1549_out);
assign _U1538_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1538 (
    .in(_U1538_in),
    .clk(_U1538_clk),
    .out(_U1538_out)
);
assign _U1539_in = _U1548_out;
_U1539_pt__U1540 _U1539 (
    .in(_U1539_in),
    .out(_U1539_out)
);
assign _U1541_in = 16'(_U1568_out * _U1573_out);
assign _U1541_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1541 (
    .in(_U1541_in),
    .clk(_U1541_clk),
    .out(_U1541_out)
);
assign _U1542_in = _U1541_out;
assign _U1542_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1542 (
    .in(_U1542_in),
    .clk(_U1542_clk),
    .out(_U1542_out)
);
assign _U1543_in = _U1542_out;
assign _U1543_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1543 (
    .in(_U1543_in),
    .clk(_U1543_clk),
    .out(_U1543_out)
);
assign _U1544_in = _U1543_out;
assign _U1544_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1544 (
    .in(_U1544_in),
    .clk(_U1544_clk),
    .out(_U1544_out)
);
assign _U1545_in = _U1544_out;
assign _U1545_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1545 (
    .in(_U1545_in),
    .clk(_U1545_clk),
    .out(_U1545_out)
);
assign _U1546_in = _U1545_out;
assign _U1546_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1546 (
    .in(_U1546_in),
    .clk(_U1546_clk),
    .out(_U1546_out)
);
assign _U1547_in = _U1546_out;
assign _U1547_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1547 (
    .in(_U1547_in),
    .clk(_U1547_clk),
    .out(_U1547_out)
);
assign _U1548_in = _U1547_out;
assign _U1548_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1548 (
    .in(_U1548_in),
    .clk(_U1548_clk),
    .out(_U1548_out)
);
assign _U1549_in = _U1551_out;
_U1549_pt__U1550 _U1549 (
    .in(_U1549_in),
    .out(_U1549_out)
);
assign _U1551_in = 16'(_U1597_out + _U1605_out);
assign _U1551_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1551 (
    .in(_U1551_in),
    .clk(_U1551_clk),
    .out(_U1551_out)
);
assign _U1552_in = in1_hw_input_global_wrapper_stencil[0];
_U1552_pt__U1553 _U1552 (
    .in(_U1552_in),
    .out(_U1552_out)
);
assign _U1554_in = _U1556_out;
_U1554_pt__U1555 _U1554 (
    .in(_U1554_in),
    .out(_U1554_out)
);
assign _U1556_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U1556_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1556 (
    .in(_U1556_in),
    .clk(_U1556_clk),
    .out(_U1556_out)
);
assign _U1557_in = _U1559_out;
_U1557_pt__U1558 _U1557 (
    .in(_U1557_in),
    .out(_U1557_out)
);
assign _U1559_in = in1_hw_input_global_wrapper_stencil[1];
assign _U1559_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1559 (
    .in(_U1559_in),
    .clk(_U1559_clk),
    .out(_U1559_out)
);
assign _U1560_in = _U1563_out;
_U1560_pt__U1561 _U1560 (
    .in(_U1560_in),
    .out(_U1560_out)
);
assign _U1562_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U1562_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1562 (
    .in(_U1562_in),
    .clk(_U1562_clk),
    .out(_U1562_out)
);
assign _U1563_in = _U1562_out;
assign _U1563_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1563 (
    .in(_U1563_in),
    .clk(_U1563_clk),
    .out(_U1563_out)
);
assign _U1564_in = _U1567_out;
_U1564_pt__U1565 _U1564 (
    .in(_U1564_in),
    .out(_U1564_out)
);
assign _U1566_in = in1_hw_input_global_wrapper_stencil[2];
assign _U1566_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1566 (
    .in(_U1566_in),
    .clk(_U1566_clk),
    .out(_U1566_out)
);
assign _U1567_in = _U1566_out;
assign _U1567_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1567 (
    .in(_U1567_in),
    .clk(_U1567_clk),
    .out(_U1567_out)
);
assign _U1568_in = _U1572_out;
_U1568_pt__U1569 _U1568 (
    .in(_U1568_in),
    .out(_U1568_out)
);
assign _U1570_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U1570_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1570 (
    .in(_U1570_in),
    .clk(_U1570_clk),
    .out(_U1570_out)
);
assign _U1571_in = _U1570_out;
assign _U1571_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1571 (
    .in(_U1571_in),
    .clk(_U1571_clk),
    .out(_U1571_out)
);
assign _U1572_in = _U1571_out;
assign _U1572_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1572 (
    .in(_U1572_in),
    .clk(_U1572_clk),
    .out(_U1572_out)
);
assign _U1573_in = _U1577_out;
_U1573_pt__U1574 _U1573 (
    .in(_U1573_in),
    .out(_U1573_out)
);
assign _U1575_in = in1_hw_input_global_wrapper_stencil[3];
assign _U1575_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1575 (
    .in(_U1575_in),
    .clk(_U1575_clk),
    .out(_U1575_out)
);
assign _U1576_in = _U1575_out;
assign _U1576_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1576 (
    .in(_U1576_in),
    .clk(_U1576_clk),
    .out(_U1576_out)
);
assign _U1577_in = _U1576_out;
assign _U1577_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1577 (
    .in(_U1577_in),
    .clk(_U1577_clk),
    .out(_U1577_out)
);
assign _U1578_in = _U1583_out;
_U1578_pt__U1579 _U1578 (
    .in(_U1578_in),
    .out(_U1578_out)
);
assign _U1580_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U1580_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1580 (
    .in(_U1580_in),
    .clk(_U1580_clk),
    .out(_U1580_out)
);
assign _U1581_in = _U1580_out;
assign _U1581_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1581 (
    .in(_U1581_in),
    .clk(_U1581_clk),
    .out(_U1581_out)
);
assign _U1582_in = _U1581_out;
assign _U1582_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1582 (
    .in(_U1582_in),
    .clk(_U1582_clk),
    .out(_U1582_out)
);
assign _U1583_in = _U1582_out;
assign _U1583_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1583 (
    .in(_U1583_in),
    .clk(_U1583_clk),
    .out(_U1583_out)
);
assign _U1584_in = _U1589_out;
_U1584_pt__U1585 _U1584 (
    .in(_U1584_in),
    .out(_U1584_out)
);
assign _U1586_in = in1_hw_input_global_wrapper_stencil[4];
assign _U1586_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1586 (
    .in(_U1586_in),
    .clk(_U1586_clk),
    .out(_U1586_out)
);
assign _U1587_in = _U1586_out;
assign _U1587_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1587 (
    .in(_U1587_in),
    .clk(_U1587_clk),
    .out(_U1587_out)
);
assign _U1588_in = _U1587_out;
assign _U1588_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1588 (
    .in(_U1588_in),
    .clk(_U1588_clk),
    .out(_U1588_out)
);
assign _U1589_in = _U1588_out;
assign _U1589_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1589 (
    .in(_U1589_in),
    .clk(_U1589_clk),
    .out(_U1589_out)
);
assign _U1590_in = _U1596_out;
_U1590_pt__U1591 _U1590 (
    .in(_U1590_in),
    .out(_U1590_out)
);
assign _U1592_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U1592_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1592 (
    .in(_U1592_in),
    .clk(_U1592_clk),
    .out(_U1592_out)
);
assign _U1593_in = _U1592_out;
assign _U1593_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1593 (
    .in(_U1593_in),
    .clk(_U1593_clk),
    .out(_U1593_out)
);
assign _U1594_in = _U1593_out;
assign _U1594_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1594 (
    .in(_U1594_in),
    .clk(_U1594_clk),
    .out(_U1594_out)
);
assign _U1595_in = _U1594_out;
assign _U1595_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1595 (
    .in(_U1595_in),
    .clk(_U1595_clk),
    .out(_U1595_out)
);
assign _U1596_in = _U1595_out;
assign _U1596_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1596 (
    .in(_U1596_in),
    .clk(_U1596_clk),
    .out(_U1596_out)
);
assign _U1597_in = _U1604_out;
_U1597_pt__U1598 _U1597 (
    .in(_U1597_in),
    .out(_U1597_out)
);
assign _U1599_in = 16'(_U1578_out * _U1584_out);
assign _U1599_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1599 (
    .in(_U1599_in),
    .clk(_U1599_clk),
    .out(_U1599_out)
);
assign _U1600_in = _U1599_out;
assign _U1600_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1600 (
    .in(_U1600_in),
    .clk(_U1600_clk),
    .out(_U1600_out)
);
assign _U1601_in = _U1600_out;
assign _U1601_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1601 (
    .in(_U1601_in),
    .clk(_U1601_clk),
    .out(_U1601_out)
);
assign _U1602_in = _U1601_out;
assign _U1602_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1602 (
    .in(_U1602_in),
    .clk(_U1602_clk),
    .out(_U1602_out)
);
assign _U1603_in = _U1602_out;
assign _U1603_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1603 (
    .in(_U1603_in),
    .clk(_U1603_clk),
    .out(_U1603_out)
);
assign _U1604_in = _U1603_out;
assign _U1604_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1604 (
    .in(_U1604_in),
    .clk(_U1604_clk),
    .out(_U1604_out)
);
assign _U1605_in = _U1607_out;
_U1605_pt__U1606 _U1605 (
    .in(_U1605_in),
    .out(_U1605_out)
);
assign _U1607_in = 16'(_U1608_out + _U1614_out);
assign _U1607_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1607 (
    .in(_U1607_in),
    .clk(_U1607_clk),
    .out(_U1607_out)
);
assign _U1608_in = _U1613_out;
_U1608_pt__U1609 _U1608 (
    .in(_U1608_in),
    .out(_U1608_out)
);
assign _U1610_in = 16'(_U1590_out * _U1458_out);
assign _U1610_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1610 (
    .in(_U1610_in),
    .clk(_U1610_clk),
    .out(_U1610_out)
);
assign _U1611_in = _U1610_out;
assign _U1611_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1611 (
    .in(_U1611_in),
    .clk(_U1611_clk),
    .out(_U1611_out)
);
assign _U1612_in = _U1611_out;
assign _U1612_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1612 (
    .in(_U1612_in),
    .clk(_U1612_clk),
    .out(_U1612_out)
);
assign _U1613_in = _U1612_out;
assign _U1613_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1613 (
    .in(_U1613_in),
    .clk(_U1613_clk),
    .out(_U1613_out)
);
assign _U1614_in = _U1616_out;
_U1614_pt__U1615 _U1614 (
    .in(_U1614_in),
    .out(_U1614_out)
);
assign _U1616_in = 16'(_U1617_out + _U1621_out);
assign _U1616_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1616 (
    .in(_U1616_in),
    .clk(_U1616_clk),
    .out(_U1616_out)
);
assign _U1617_in = _U1620_out;
_U1617_pt__U1618 _U1617 (
    .in(_U1617_in),
    .out(_U1617_out)
);
assign _U1619_in = 16'(_U1465_out * _U1473_out);
assign _U1619_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1619 (
    .in(_U1619_in),
    .clk(_U1619_clk),
    .out(_U1619_out)
);
assign _U1620_in = _U1619_out;
assign _U1620_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1620 (
    .in(_U1620_in),
    .clk(_U1620_clk),
    .out(_U1620_out)
);
assign _U1621_in = _U1623_out;
_U1621_pt__U1622 _U1621 (
    .in(_U1621_in),
    .out(_U1621_out)
);
assign _U1623_in = 16'(_U1481_out * _U1490_out);
assign _U1623_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1623 (
    .in(_U1623_in),
    .clk(_U1623_clk),
    .out(_U1623_out)
);
assign _U1624_in = _U1639_out;
_U1624_pt__U1625 _U1624 (
    .in(_U1624_in),
    .out(_U1624_out)
);
assign _U1626_in = in0_conv_stencil[0];
assign _U1626_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1626 (
    .in(_U1626_in),
    .clk(_U1626_clk),
    .out(_U1626_out)
);
assign _U1627_in = _U1626_out;
assign _U1627_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1627 (
    .in(_U1627_in),
    .clk(_U1627_clk),
    .out(_U1627_out)
);
assign _U1628_in = _U1627_out;
assign _U1628_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1628 (
    .in(_U1628_in),
    .clk(_U1628_clk),
    .out(_U1628_out)
);
assign _U1629_in = _U1628_out;
assign _U1629_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1629 (
    .in(_U1629_in),
    .clk(_U1629_clk),
    .out(_U1629_out)
);
assign _U1630_in = _U1629_out;
assign _U1630_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1630 (
    .in(_U1630_in),
    .clk(_U1630_clk),
    .out(_U1630_out)
);
assign _U1631_in = _U1630_out;
assign _U1631_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1631 (
    .in(_U1631_in),
    .clk(_U1631_clk),
    .out(_U1631_out)
);
assign _U1632_in = _U1631_out;
assign _U1632_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1632 (
    .in(_U1632_in),
    .clk(_U1632_clk),
    .out(_U1632_out)
);
assign _U1633_in = _U1632_out;
assign _U1633_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1633 (
    .in(_U1633_in),
    .clk(_U1633_clk),
    .out(_U1633_out)
);
assign _U1634_in = _U1633_out;
assign _U1634_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1634 (
    .in(_U1634_in),
    .clk(_U1634_clk),
    .out(_U1634_out)
);
assign _U1635_in = _U1634_out;
assign _U1635_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1635 (
    .in(_U1635_in),
    .clk(_U1635_clk),
    .out(_U1635_out)
);
assign _U1636_in = _U1635_out;
assign _U1636_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1636 (
    .in(_U1636_in),
    .clk(_U1636_clk),
    .out(_U1636_out)
);
assign _U1637_in = _U1636_out;
assign _U1637_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1637 (
    .in(_U1637_in),
    .clk(_U1637_clk),
    .out(_U1637_out)
);
assign _U1638_in = _U1637_out;
assign _U1638_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1638 (
    .in(_U1638_in),
    .clk(_U1638_clk),
    .out(_U1638_out)
);
assign _U1639_in = _U1638_out;
assign _U1639_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1639 (
    .in(_U1639_in),
    .clk(_U1639_clk),
    .out(_U1639_out)
);
assign _U1640_in = in2_hw_kernel_global_wrapper_stencil[0];
_U1640_pt__U1641 _U1640 (
    .in(_U1640_in),
    .out(_U1640_out)
);
endmodule

module cu_op_hcompute_conv_stencil_15 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_15_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_15_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_15_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[0];
hcompute_conv_stencil_15_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_15_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U143_pt__U144 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1430_pt__U1431 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1427_pt__U1428 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U141_pt__U142 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1417_pt__U1418 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1414_pt__U1415 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1402_pt__U1403 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1399_pt__U1400 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U138_pt__U139 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1385_pt__U1386 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1382_pt__U1383 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1376_pt__U1377 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1370_pt__U1371 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1365_pt__U1366 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1360_pt__U1361 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1356_pt__U1357 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1352_pt__U1353 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1349_pt__U1350 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1346_pt__U1347 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1344_pt__U1345 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1335_pt__U1336 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1326_pt__U1327 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1318_pt__U1319 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1310_pt__U1311 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U12_pt__U13 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_6_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
wire [15:0] _U12_in;
assign _U12_in = in0_hw_input_stencil[0];
_U12_pt__U13 _U12 (
    .in(_U12_in),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil_6 (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read[0];
hcompute_hw_input_global_wrapper_stencil_6_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U1294_pt__U1295 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1289_pt__U1290 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1283_pt__U1284 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1280_pt__U1281 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1272_pt__U1273 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1270_pt__U1271 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1267_pt__U1268 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1260_pt__U1261 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1253_pt__U1254 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1250_pt__U1251 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1242_pt__U1243 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1240_pt__U1241 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_14_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U1240_in;
wire [15:0] _U1240_out;
wire [15:0] _U1242_in;
wire [15:0] _U1242_out;
wire [15:0] _U1244_in;
wire _U1244_clk;
wire [15:0] _U1244_out;
wire [15:0] _U1245_in;
wire _U1245_clk;
wire [15:0] _U1245_out;
wire [15:0] _U1246_in;
wire _U1246_clk;
wire [15:0] _U1246_out;
wire [15:0] _U1247_in;
wire _U1247_clk;
wire [15:0] _U1247_out;
wire [15:0] _U1248_in;
wire _U1248_clk;
wire [15:0] _U1248_out;
wire [15:0] _U1249_in;
wire _U1249_clk;
wire [15:0] _U1249_out;
wire [15:0] _U1250_in;
wire [15:0] _U1250_out;
wire [15:0] _U1252_in;
wire _U1252_clk;
wire [15:0] _U1252_out;
wire [15:0] _U1253_in;
wire [15:0] _U1253_out;
wire [15:0] _U1255_in;
wire _U1255_clk;
wire [15:0] _U1255_out;
wire [15:0] _U1256_in;
wire _U1256_clk;
wire [15:0] _U1256_out;
wire [15:0] _U1257_in;
wire _U1257_clk;
wire [15:0] _U1257_out;
wire [15:0] _U1258_in;
wire _U1258_clk;
wire [15:0] _U1258_out;
wire [15:0] _U1259_in;
wire _U1259_clk;
wire [15:0] _U1259_out;
wire [15:0] _U1260_in;
wire [15:0] _U1260_out;
wire [15:0] _U1262_in;
wire _U1262_clk;
wire [15:0] _U1262_out;
wire [15:0] _U1263_in;
wire _U1263_clk;
wire [15:0] _U1263_out;
wire [15:0] _U1264_in;
wire _U1264_clk;
wire [15:0] _U1264_out;
wire [15:0] _U1265_in;
wire _U1265_clk;
wire [15:0] _U1265_out;
wire [15:0] _U1266_in;
wire _U1266_clk;
wire [15:0] _U1266_out;
wire [15:0] _U1267_in;
wire [15:0] _U1267_out;
wire [15:0] _U1269_in;
wire _U1269_clk;
wire [15:0] _U1269_out;
wire [15:0] _U1270_in;
wire [15:0] _U1272_in;
wire [15:0] _U1272_out;
wire [15:0] _U1274_in;
wire _U1274_clk;
wire [15:0] _U1274_out;
wire [15:0] _U1275_in;
wire _U1275_clk;
wire [15:0] _U1275_out;
wire [15:0] _U1276_in;
wire _U1276_clk;
wire [15:0] _U1276_out;
wire [15:0] _U1277_in;
wire _U1277_clk;
wire [15:0] _U1277_out;
wire [15:0] _U1278_in;
wire _U1278_clk;
wire [15:0] _U1278_out;
wire [15:0] _U1279_in;
wire _U1279_clk;
wire [15:0] _U1279_out;
wire [15:0] _U1280_in;
wire [15:0] _U1280_out;
wire [15:0] _U1282_in;
wire _U1282_clk;
wire [15:0] _U1282_out;
wire [15:0] _U1283_in;
wire [15:0] _U1283_out;
wire [15:0] _U1285_in;
wire _U1285_clk;
wire [15:0] _U1285_out;
wire [15:0] _U1286_in;
wire _U1286_clk;
wire [15:0] _U1286_out;
wire [15:0] _U1287_in;
wire _U1287_clk;
wire [15:0] _U1287_out;
wire [15:0] _U1288_in;
wire _U1288_clk;
wire [15:0] _U1288_out;
wire [15:0] _U1289_in;
wire [15:0] _U1289_out;
wire [15:0] _U1291_in;
wire _U1291_clk;
wire [15:0] _U1291_out;
wire [15:0] _U1292_in;
wire _U1292_clk;
wire [15:0] _U1292_out;
wire [15:0] _U1293_in;
wire _U1293_clk;
wire [15:0] _U1293_out;
wire [15:0] _U1294_in;
wire [15:0] _U1294_out;
wire [15:0] _U1296_in;
wire _U1296_clk;
wire [15:0] _U1296_out;
wire [15:0] _U1297_in;
wire _U1297_clk;
wire [15:0] _U1297_out;
wire [15:0] _U1298_in;
wire _U1298_clk;
wire [15:0] _U1298_out;
wire [15:0] _U1299_in;
wire _U1299_clk;
wire [15:0] _U1299_out;
wire [15:0] _U1300_in;
wire _U1300_clk;
wire [15:0] _U1300_out;
wire [15:0] _U1301_in;
wire _U1301_clk;
wire [15:0] _U1301_out;
wire [15:0] _U1302_in;
wire _U1302_clk;
wire [15:0] _U1302_out;
wire [15:0] _U1303_in;
wire _U1303_clk;
wire [15:0] _U1303_out;
wire [15:0] _U1304_in;
wire _U1304_clk;
wire [15:0] _U1304_out;
wire [15:0] _U1305_in;
wire _U1305_clk;
wire [15:0] _U1305_out;
wire [15:0] _U1306_in;
wire _U1306_clk;
wire [15:0] _U1306_out;
wire [15:0] _U1307_in;
wire _U1307_clk;
wire [15:0] _U1307_out;
wire [15:0] _U1308_in;
wire _U1308_clk;
wire [15:0] _U1308_out;
wire [15:0] _U1309_in;
wire _U1309_clk;
wire [15:0] _U1309_out;
wire [15:0] _U1310_in;
wire [15:0] _U1310_out;
wire [15:0] _U1312_in;
wire _U1312_clk;
wire [15:0] _U1312_out;
wire [15:0] _U1313_in;
wire _U1313_clk;
wire [15:0] _U1313_out;
wire [15:0] _U1314_in;
wire _U1314_clk;
wire [15:0] _U1314_out;
wire [15:0] _U1315_in;
wire _U1315_clk;
wire [15:0] _U1315_out;
wire [15:0] _U1316_in;
wire _U1316_clk;
wire [15:0] _U1316_out;
wire [15:0] _U1317_in;
wire _U1317_clk;
wire [15:0] _U1317_out;
wire [15:0] _U1318_in;
wire [15:0] _U1318_out;
wire [15:0] _U1320_in;
wire _U1320_clk;
wire [15:0] _U1320_out;
wire [15:0] _U1321_in;
wire _U1321_clk;
wire [15:0] _U1321_out;
wire [15:0] _U1322_in;
wire _U1322_clk;
wire [15:0] _U1322_out;
wire [15:0] _U1323_in;
wire _U1323_clk;
wire [15:0] _U1323_out;
wire [15:0] _U1324_in;
wire _U1324_clk;
wire [15:0] _U1324_out;
wire [15:0] _U1325_in;
wire _U1325_clk;
wire [15:0] _U1325_out;
wire [15:0] _U1326_in;
wire [15:0] _U1326_out;
wire [15:0] _U1328_in;
wire _U1328_clk;
wire [15:0] _U1328_out;
wire [15:0] _U1329_in;
wire _U1329_clk;
wire [15:0] _U1329_out;
wire [15:0] _U1330_in;
wire _U1330_clk;
wire [15:0] _U1330_out;
wire [15:0] _U1331_in;
wire _U1331_clk;
wire [15:0] _U1331_out;
wire [15:0] _U1332_in;
wire _U1332_clk;
wire [15:0] _U1332_out;
wire [15:0] _U1333_in;
wire _U1333_clk;
wire [15:0] _U1333_out;
wire [15:0] _U1334_in;
wire _U1334_clk;
wire [15:0] _U1334_out;
wire [15:0] _U1335_in;
wire [15:0] _U1335_out;
wire [15:0] _U1337_in;
wire _U1337_clk;
wire [15:0] _U1337_out;
wire [15:0] _U1338_in;
wire _U1338_clk;
wire [15:0] _U1338_out;
wire [15:0] _U1339_in;
wire _U1339_clk;
wire [15:0] _U1339_out;
wire [15:0] _U1340_in;
wire _U1340_clk;
wire [15:0] _U1340_out;
wire [15:0] _U1341_in;
wire _U1341_clk;
wire [15:0] _U1341_out;
wire [15:0] _U1342_in;
wire _U1342_clk;
wire [15:0] _U1342_out;
wire [15:0] _U1343_in;
wire _U1343_clk;
wire [15:0] _U1343_out;
wire [15:0] _U1344_in;
wire [15:0] _U1344_out;
wire [15:0] _U1346_in;
wire [15:0] _U1346_out;
wire [15:0] _U1348_in;
wire _U1348_clk;
wire [15:0] _U1348_out;
wire [15:0] _U1349_in;
wire [15:0] _U1349_out;
wire [15:0] _U1351_in;
wire _U1351_clk;
wire [15:0] _U1351_out;
wire [15:0] _U1352_in;
wire [15:0] _U1352_out;
wire [15:0] _U1354_in;
wire _U1354_clk;
wire [15:0] _U1354_out;
wire [15:0] _U1355_in;
wire _U1355_clk;
wire [15:0] _U1355_out;
wire [15:0] _U1356_in;
wire [15:0] _U1356_out;
wire [15:0] _U1358_in;
wire _U1358_clk;
wire [15:0] _U1358_out;
wire [15:0] _U1359_in;
wire _U1359_clk;
wire [15:0] _U1359_out;
wire [15:0] _U1360_in;
wire [15:0] _U1360_out;
wire [15:0] _U1362_in;
wire _U1362_clk;
wire [15:0] _U1362_out;
wire [15:0] _U1363_in;
wire _U1363_clk;
wire [15:0] _U1363_out;
wire [15:0] _U1364_in;
wire _U1364_clk;
wire [15:0] _U1364_out;
wire [15:0] _U1365_in;
wire [15:0] _U1365_out;
wire [15:0] _U1367_in;
wire _U1367_clk;
wire [15:0] _U1367_out;
wire [15:0] _U1368_in;
wire _U1368_clk;
wire [15:0] _U1368_out;
wire [15:0] _U1369_in;
wire _U1369_clk;
wire [15:0] _U1369_out;
wire [15:0] _U1370_in;
wire [15:0] _U1370_out;
wire [15:0] _U1372_in;
wire _U1372_clk;
wire [15:0] _U1372_out;
wire [15:0] _U1373_in;
wire _U1373_clk;
wire [15:0] _U1373_out;
wire [15:0] _U1374_in;
wire _U1374_clk;
wire [15:0] _U1374_out;
wire [15:0] _U1375_in;
wire _U1375_clk;
wire [15:0] _U1375_out;
wire [15:0] _U1376_in;
wire [15:0] _U1376_out;
wire [15:0] _U1378_in;
wire _U1378_clk;
wire [15:0] _U1378_out;
wire [15:0] _U1379_in;
wire _U1379_clk;
wire [15:0] _U1379_out;
wire [15:0] _U1380_in;
wire _U1380_clk;
wire [15:0] _U1380_out;
wire [15:0] _U1381_in;
wire _U1381_clk;
wire [15:0] _U1381_out;
wire [15:0] _U1382_in;
wire [15:0] _U1382_out;
wire [15:0] _U1384_in;
wire _U1384_clk;
wire [15:0] _U1384_out;
wire [15:0] _U1385_in;
wire [15:0] _U1385_out;
wire [15:0] _U1387_in;
wire _U1387_clk;
wire [15:0] _U1387_out;
wire [15:0] _U1388_in;
wire _U1388_clk;
wire [15:0] _U1388_out;
wire [15:0] _U1389_in;
wire _U1389_clk;
wire [15:0] _U1389_out;
wire [15:0] _U1390_in;
wire _U1390_clk;
wire [15:0] _U1390_out;
wire [15:0] _U1391_in;
wire _U1391_clk;
wire [15:0] _U1391_out;
wire [15:0] _U1392_in;
wire _U1392_clk;
wire [15:0] _U1392_out;
wire [15:0] _U1393_in;
wire _U1393_clk;
wire [15:0] _U1393_out;
wire [15:0] _U1394_in;
wire _U1394_clk;
wire [15:0] _U1394_out;
wire [15:0] _U1395_in;
wire _U1395_clk;
wire [15:0] _U1395_out;
wire [15:0] _U1396_in;
wire _U1396_clk;
wire [15:0] _U1396_out;
wire [15:0] _U1397_in;
wire _U1397_clk;
wire [15:0] _U1397_out;
wire [15:0] _U1398_in;
wire _U1398_clk;
wire [15:0] _U1398_out;
wire [15:0] _U1399_in;
wire [15:0] _U1399_out;
wire [15:0] _U1401_in;
wire _U1401_clk;
wire [15:0] _U1401_out;
wire [15:0] _U1402_in;
wire [15:0] _U1402_out;
wire [15:0] _U1404_in;
wire _U1404_clk;
wire [15:0] _U1404_out;
wire [15:0] _U1405_in;
wire _U1405_clk;
wire [15:0] _U1405_out;
wire [15:0] _U1406_in;
wire _U1406_clk;
wire [15:0] _U1406_out;
wire [15:0] _U1407_in;
wire _U1407_clk;
wire [15:0] _U1407_out;
wire [15:0] _U1408_in;
wire _U1408_clk;
wire [15:0] _U1408_out;
wire [15:0] _U1409_in;
wire _U1409_clk;
wire [15:0] _U1409_out;
wire [15:0] _U1410_in;
wire _U1410_clk;
wire [15:0] _U1410_out;
wire [15:0] _U1411_in;
wire _U1411_clk;
wire [15:0] _U1411_out;
wire [15:0] _U1412_in;
wire _U1412_clk;
wire [15:0] _U1412_out;
wire [15:0] _U1413_in;
wire _U1413_clk;
wire [15:0] _U1413_out;
wire [15:0] _U1414_in;
wire [15:0] _U1414_out;
wire [15:0] _U1416_in;
wire _U1416_clk;
wire [15:0] _U1416_out;
wire [15:0] _U1417_in;
wire [15:0] _U1417_out;
wire [15:0] _U1419_in;
wire _U1419_clk;
wire [15:0] _U1419_out;
wire [15:0] _U1420_in;
wire _U1420_clk;
wire [15:0] _U1420_out;
wire [15:0] _U1421_in;
wire _U1421_clk;
wire [15:0] _U1421_out;
wire [15:0] _U1422_in;
wire _U1422_clk;
wire [15:0] _U1422_out;
wire [15:0] _U1423_in;
wire _U1423_clk;
wire [15:0] _U1423_out;
wire [15:0] _U1424_in;
wire _U1424_clk;
wire [15:0] _U1424_out;
wire [15:0] _U1425_in;
wire _U1425_clk;
wire [15:0] _U1425_out;
wire [15:0] _U1426_in;
wire _U1426_clk;
wire [15:0] _U1426_out;
wire [15:0] _U1427_in;
wire [15:0] _U1427_out;
wire [15:0] _U1429_in;
wire _U1429_clk;
wire [15:0] _U1429_out;
wire [15:0] _U1430_in;
wire [15:0] _U1430_out;
wire [15:0] _U1432_in;
wire _U1432_clk;
wire [15:0] _U1432_out;
wire [15:0] _U1433_in;
wire _U1433_clk;
wire [15:0] _U1433_out;
wire [15:0] _U1434_in;
wire _U1434_clk;
wire [15:0] _U1434_out;
wire [15:0] _U1435_in;
wire _U1435_clk;
wire [15:0] _U1435_out;
wire [15:0] _U1436_in;
wire _U1436_clk;
wire [15:0] _U1436_out;
wire [15:0] _U1437_in;
wire _U1437_clk;
wire [15:0] _U1437_out;
wire [15:0] _U1438_in;
wire _U1438_clk;
wire [15:0] _U1438_out;
wire [15:0] _U1439_in;
wire _U1439_clk;
wire [15:0] _U1439_out;
wire [15:0] _U1440_in;
wire _U1440_clk;
wire [15:0] _U1440_out;
assign _U1240_in = in2_hw_kernel_global_wrapper_stencil[2];
_U1240_pt__U1241 _U1240 (
    .in(_U1240_in),
    .out(_U1240_out)
);
assign _U1242_in = _U1249_out;
_U1242_pt__U1243 _U1242 (
    .in(_U1242_in),
    .out(_U1242_out)
);
assign _U1244_in = 16'(_U1360_out * _U1365_out);
assign _U1244_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1244 (
    .in(_U1244_in),
    .clk(_U1244_clk),
    .out(_U1244_out)
);
assign _U1245_in = _U1244_out;
assign _U1245_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1245 (
    .in(_U1245_in),
    .clk(_U1245_clk),
    .out(_U1245_out)
);
assign _U1246_in = _U1245_out;
assign _U1246_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1246 (
    .in(_U1246_in),
    .clk(_U1246_clk),
    .out(_U1246_out)
);
assign _U1247_in = _U1246_out;
assign _U1247_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1247 (
    .in(_U1247_in),
    .clk(_U1247_clk),
    .out(_U1247_out)
);
assign _U1248_in = _U1247_out;
assign _U1248_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1248 (
    .in(_U1248_in),
    .clk(_U1248_clk),
    .out(_U1248_out)
);
assign _U1249_in = _U1248_out;
assign _U1249_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1249 (
    .in(_U1249_in),
    .clk(_U1249_clk),
    .out(_U1249_out)
);
assign _U1250_in = _U1252_out;
_U1250_pt__U1251 _U1250 (
    .in(_U1250_in),
    .out(_U1250_out)
);
assign _U1252_in = 16'(_U1385_out + _U1399_out);
assign _U1252_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1252 (
    .in(_U1252_in),
    .clk(_U1252_clk),
    .out(_U1252_out)
);
assign _U1253_in = _U1259_out;
_U1253_pt__U1254 _U1253 (
    .in(_U1253_in),
    .out(_U1253_out)
);
assign _U1255_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U1255_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1255 (
    .in(_U1255_in),
    .clk(_U1255_clk),
    .out(_U1255_out)
);
assign _U1256_in = _U1255_out;
assign _U1256_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1256 (
    .in(_U1256_in),
    .clk(_U1256_clk),
    .out(_U1256_out)
);
assign _U1257_in = _U1256_out;
assign _U1257_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1257 (
    .in(_U1257_in),
    .clk(_U1257_clk),
    .out(_U1257_out)
);
assign _U1258_in = _U1257_out;
assign _U1258_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1258 (
    .in(_U1258_in),
    .clk(_U1258_clk),
    .out(_U1258_out)
);
assign _U1259_in = _U1258_out;
assign _U1259_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1259 (
    .in(_U1259_in),
    .clk(_U1259_clk),
    .out(_U1259_out)
);
assign _U1260_in = _U1266_out;
_U1260_pt__U1261 _U1260 (
    .in(_U1260_in),
    .out(_U1260_out)
);
assign _U1262_in = in1_hw_input_global_wrapper_stencil[7];
assign _U1262_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1262 (
    .in(_U1262_in),
    .clk(_U1262_clk),
    .out(_U1262_out)
);
assign _U1263_in = _U1262_out;
assign _U1263_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1263 (
    .in(_U1263_in),
    .clk(_U1263_clk),
    .out(_U1263_out)
);
assign _U1264_in = _U1263_out;
assign _U1264_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1264 (
    .in(_U1264_in),
    .clk(_U1264_clk),
    .out(_U1264_out)
);
assign _U1265_in = _U1264_out;
assign _U1265_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1265 (
    .in(_U1265_in),
    .clk(_U1265_clk),
    .out(_U1265_out)
);
assign _U1266_in = _U1265_out;
assign _U1266_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1266 (
    .in(_U1266_in),
    .clk(_U1266_clk),
    .out(_U1266_out)
);
assign _U1267_in = _U1269_out;
_U1267_pt__U1268 _U1267 (
    .in(_U1267_in),
    .out(_U1267_out)
);
assign _U1269_in = 16'(_U1294_out + _U1382_out);
assign _U1269_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1269 (
    .in(_U1269_in),
    .clk(_U1269_clk),
    .out(_U1269_out)
);
assign _U1270_in = 16'(_U1430_out + _U1267_out);
_U1270_pt__U1271 _U1270 (
    .in(_U1270_in),
    .out(out_conv_stencil)
);
assign _U1272_in = _U1279_out;
_U1272_pt__U1273 _U1272 (
    .in(_U1272_in),
    .out(_U1272_out)
);
assign _U1274_in = 16'(_U1326_out * _U1335_out);
assign _U1274_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1274 (
    .in(_U1274_in),
    .clk(_U1274_clk),
    .out(_U1274_out)
);
assign _U1275_in = _U1274_out;
assign _U1275_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1275 (
    .in(_U1275_in),
    .clk(_U1275_clk),
    .out(_U1275_out)
);
assign _U1276_in = _U1275_out;
assign _U1276_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1276 (
    .in(_U1276_in),
    .clk(_U1276_clk),
    .out(_U1276_out)
);
assign _U1277_in = _U1276_out;
assign _U1277_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1277 (
    .in(_U1277_in),
    .clk(_U1277_clk),
    .out(_U1277_out)
);
assign _U1278_in = _U1277_out;
assign _U1278_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1278 (
    .in(_U1278_in),
    .clk(_U1278_clk),
    .out(_U1278_out)
);
assign _U1279_in = _U1278_out;
assign _U1279_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1279 (
    .in(_U1279_in),
    .clk(_U1279_clk),
    .out(_U1279_out)
);
assign _U1280_in = _U1282_out;
_U1280_pt__U1281 _U1280 (
    .in(_U1280_in),
    .out(_U1280_out)
);
assign _U1282_in = 16'(_U1283_out + _U1289_out);
assign _U1282_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1282 (
    .in(_U1282_in),
    .clk(_U1282_clk),
    .out(_U1282_out)
);
assign _U1283_in = _U1288_out;
_U1283_pt__U1284 _U1283 (
    .in(_U1283_in),
    .out(_U1283_out)
);
assign _U1285_in = 16'(_U1370_out * _U1376_out);
assign _U1285_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1285 (
    .in(_U1285_in),
    .clk(_U1285_clk),
    .out(_U1285_out)
);
assign _U1286_in = _U1285_out;
assign _U1286_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1286 (
    .in(_U1286_in),
    .clk(_U1286_clk),
    .out(_U1286_out)
);
assign _U1287_in = _U1286_out;
assign _U1287_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1287 (
    .in(_U1287_in),
    .clk(_U1287_clk),
    .out(_U1287_out)
);
assign _U1288_in = _U1287_out;
assign _U1288_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1288 (
    .in(_U1288_in),
    .clk(_U1288_clk),
    .out(_U1288_out)
);
assign _U1289_in = _U1293_out;
_U1289_pt__U1290 _U1289 (
    .in(_U1289_in),
    .out(_U1289_out)
);
assign _U1291_in = 16'(_U1253_out * _U1260_out);
assign _U1291_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1291 (
    .in(_U1291_in),
    .clk(_U1291_clk),
    .out(_U1291_out)
);
assign _U1292_in = _U1291_out;
assign _U1292_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1292 (
    .in(_U1292_in),
    .clk(_U1292_clk),
    .out(_U1292_out)
);
assign _U1293_in = _U1292_out;
assign _U1293_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1293 (
    .in(_U1293_in),
    .clk(_U1293_clk),
    .out(_U1293_out)
);
assign _U1294_in = _U1309_out;
_U1294_pt__U1295 _U1294 (
    .in(_U1294_in),
    .out(_U1294_out)
);
assign _U1296_in = in0_conv_stencil[0];
assign _U1296_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1296 (
    .in(_U1296_in),
    .clk(_U1296_clk),
    .out(_U1296_out)
);
assign _U1297_in = _U1296_out;
assign _U1297_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1297 (
    .in(_U1297_in),
    .clk(_U1297_clk),
    .out(_U1297_out)
);
assign _U1298_in = _U1297_out;
assign _U1298_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1298 (
    .in(_U1298_in),
    .clk(_U1298_clk),
    .out(_U1298_out)
);
assign _U1299_in = _U1298_out;
assign _U1299_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1299 (
    .in(_U1299_in),
    .clk(_U1299_clk),
    .out(_U1299_out)
);
assign _U1300_in = _U1299_out;
assign _U1300_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1300 (
    .in(_U1300_in),
    .clk(_U1300_clk),
    .out(_U1300_out)
);
assign _U1301_in = _U1300_out;
assign _U1301_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1301 (
    .in(_U1301_in),
    .clk(_U1301_clk),
    .out(_U1301_out)
);
assign _U1302_in = _U1301_out;
assign _U1302_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1302 (
    .in(_U1302_in),
    .clk(_U1302_clk),
    .out(_U1302_out)
);
assign _U1303_in = _U1302_out;
assign _U1303_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1303 (
    .in(_U1303_in),
    .clk(_U1303_clk),
    .out(_U1303_out)
);
assign _U1304_in = _U1303_out;
assign _U1304_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1304 (
    .in(_U1304_in),
    .clk(_U1304_clk),
    .out(_U1304_out)
);
assign _U1305_in = _U1304_out;
assign _U1305_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1305 (
    .in(_U1305_in),
    .clk(_U1305_clk),
    .out(_U1305_out)
);
assign _U1306_in = _U1305_out;
assign _U1306_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1306 (
    .in(_U1306_in),
    .clk(_U1306_clk),
    .out(_U1306_out)
);
assign _U1307_in = _U1306_out;
assign _U1307_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1307 (
    .in(_U1307_in),
    .clk(_U1307_clk),
    .out(_U1307_out)
);
assign _U1308_in = _U1307_out;
assign _U1308_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1308 (
    .in(_U1308_in),
    .clk(_U1308_clk),
    .out(_U1308_out)
);
assign _U1309_in = _U1308_out;
assign _U1309_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1309 (
    .in(_U1309_in),
    .clk(_U1309_clk),
    .out(_U1309_out)
);
assign _U1310_in = _U1317_out;
_U1310_pt__U1311 _U1310 (
    .in(_U1310_in),
    .out(_U1310_out)
);
assign _U1312_in = in2_hw_kernel_global_wrapper_stencil[0];
assign _U1312_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1312 (
    .in(_U1312_in),
    .clk(_U1312_clk),
    .out(_U1312_out)
);
assign _U1313_in = _U1312_out;
assign _U1313_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1313 (
    .in(_U1313_in),
    .clk(_U1313_clk),
    .out(_U1313_out)
);
assign _U1314_in = _U1313_out;
assign _U1314_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1314 (
    .in(_U1314_in),
    .clk(_U1314_clk),
    .out(_U1314_out)
);
assign _U1315_in = _U1314_out;
assign _U1315_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1315 (
    .in(_U1315_in),
    .clk(_U1315_clk),
    .out(_U1315_out)
);
assign _U1316_in = _U1315_out;
assign _U1316_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1316 (
    .in(_U1316_in),
    .clk(_U1316_clk),
    .out(_U1316_out)
);
assign _U1317_in = _U1316_out;
assign _U1317_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1317 (
    .in(_U1317_in),
    .clk(_U1317_clk),
    .out(_U1317_out)
);
assign _U1318_in = _U1325_out;
_U1318_pt__U1319 _U1318 (
    .in(_U1318_in),
    .out(_U1318_out)
);
assign _U1320_in = in1_hw_input_global_wrapper_stencil[0];
assign _U1320_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1320 (
    .in(_U1320_in),
    .clk(_U1320_clk),
    .out(_U1320_out)
);
assign _U1321_in = _U1320_out;
assign _U1321_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1321 (
    .in(_U1321_in),
    .clk(_U1321_clk),
    .out(_U1321_out)
);
assign _U1322_in = _U1321_out;
assign _U1322_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1322 (
    .in(_U1322_in),
    .clk(_U1322_clk),
    .out(_U1322_out)
);
assign _U1323_in = _U1322_out;
assign _U1323_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1323 (
    .in(_U1323_in),
    .clk(_U1323_clk),
    .out(_U1323_out)
);
assign _U1324_in = _U1323_out;
assign _U1324_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1324 (
    .in(_U1324_in),
    .clk(_U1324_clk),
    .out(_U1324_out)
);
assign _U1325_in = _U1324_out;
assign _U1325_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1325 (
    .in(_U1325_in),
    .clk(_U1325_clk),
    .out(_U1325_out)
);
assign _U1326_in = _U1334_out;
_U1326_pt__U1327 _U1326 (
    .in(_U1326_in),
    .out(_U1326_out)
);
assign _U1328_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U1328_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1328 (
    .in(_U1328_in),
    .clk(_U1328_clk),
    .out(_U1328_out)
);
assign _U1329_in = _U1328_out;
assign _U1329_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1329 (
    .in(_U1329_in),
    .clk(_U1329_clk),
    .out(_U1329_out)
);
assign _U1330_in = _U1329_out;
assign _U1330_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1330 (
    .in(_U1330_in),
    .clk(_U1330_clk),
    .out(_U1330_out)
);
assign _U1331_in = _U1330_out;
assign _U1331_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1331 (
    .in(_U1331_in),
    .clk(_U1331_clk),
    .out(_U1331_out)
);
assign _U1332_in = _U1331_out;
assign _U1332_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1332 (
    .in(_U1332_in),
    .clk(_U1332_clk),
    .out(_U1332_out)
);
assign _U1333_in = _U1332_out;
assign _U1333_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1333 (
    .in(_U1333_in),
    .clk(_U1333_clk),
    .out(_U1333_out)
);
assign _U1334_in = _U1333_out;
assign _U1334_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1334 (
    .in(_U1334_in),
    .clk(_U1334_clk),
    .out(_U1334_out)
);
assign _U1335_in = _U1343_out;
_U1335_pt__U1336 _U1335 (
    .in(_U1335_in),
    .out(_U1335_out)
);
assign _U1337_in = in1_hw_input_global_wrapper_stencil[1];
assign _U1337_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1337 (
    .in(_U1337_in),
    .clk(_U1337_clk),
    .out(_U1337_out)
);
assign _U1338_in = _U1337_out;
assign _U1338_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1338 (
    .in(_U1338_in),
    .clk(_U1338_clk),
    .out(_U1338_out)
);
assign _U1339_in = _U1338_out;
assign _U1339_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1339 (
    .in(_U1339_in),
    .clk(_U1339_clk),
    .out(_U1339_out)
);
assign _U1340_in = _U1339_out;
assign _U1340_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1340 (
    .in(_U1340_in),
    .clk(_U1340_clk),
    .out(_U1340_out)
);
assign _U1341_in = _U1340_out;
assign _U1341_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1341 (
    .in(_U1341_in),
    .clk(_U1341_clk),
    .out(_U1341_out)
);
assign _U1342_in = _U1341_out;
assign _U1342_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1342 (
    .in(_U1342_in),
    .clk(_U1342_clk),
    .out(_U1342_out)
);
assign _U1343_in = _U1342_out;
assign _U1343_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1343 (
    .in(_U1343_in),
    .clk(_U1343_clk),
    .out(_U1343_out)
);
assign _U1344_in = in1_hw_input_global_wrapper_stencil[2];
_U1344_pt__U1345 _U1344 (
    .in(_U1344_in),
    .out(_U1344_out)
);
assign _U1346_in = _U1348_out;
_U1346_pt__U1347 _U1346 (
    .in(_U1346_in),
    .out(_U1346_out)
);
assign _U1348_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U1348_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1348 (
    .in(_U1348_in),
    .clk(_U1348_clk),
    .out(_U1348_out)
);
assign _U1349_in = _U1351_out;
_U1349_pt__U1350 _U1349 (
    .in(_U1349_in),
    .out(_U1349_out)
);
assign _U1351_in = in1_hw_input_global_wrapper_stencil[3];
assign _U1351_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1351 (
    .in(_U1351_in),
    .clk(_U1351_clk),
    .out(_U1351_out)
);
assign _U1352_in = _U1355_out;
_U1352_pt__U1353 _U1352 (
    .in(_U1352_in),
    .out(_U1352_out)
);
assign _U1354_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U1354_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1354 (
    .in(_U1354_in),
    .clk(_U1354_clk),
    .out(_U1354_out)
);
assign _U1355_in = _U1354_out;
assign _U1355_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1355 (
    .in(_U1355_in),
    .clk(_U1355_clk),
    .out(_U1355_out)
);
assign _U1356_in = _U1359_out;
_U1356_pt__U1357 _U1356 (
    .in(_U1356_in),
    .out(_U1356_out)
);
assign _U1358_in = in1_hw_input_global_wrapper_stencil[4];
assign _U1358_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1358 (
    .in(_U1358_in),
    .clk(_U1358_clk),
    .out(_U1358_out)
);
assign _U1359_in = _U1358_out;
assign _U1359_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1359 (
    .in(_U1359_in),
    .clk(_U1359_clk),
    .out(_U1359_out)
);
assign _U1360_in = _U1364_out;
_U1360_pt__U1361 _U1360 (
    .in(_U1360_in),
    .out(_U1360_out)
);
assign _U1362_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U1362_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1362 (
    .in(_U1362_in),
    .clk(_U1362_clk),
    .out(_U1362_out)
);
assign _U1363_in = _U1362_out;
assign _U1363_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1363 (
    .in(_U1363_in),
    .clk(_U1363_clk),
    .out(_U1363_out)
);
assign _U1364_in = _U1363_out;
assign _U1364_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1364 (
    .in(_U1364_in),
    .clk(_U1364_clk),
    .out(_U1364_out)
);
assign _U1365_in = _U1369_out;
_U1365_pt__U1366 _U1365 (
    .in(_U1365_in),
    .out(_U1365_out)
);
assign _U1367_in = in1_hw_input_global_wrapper_stencil[5];
assign _U1367_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1367 (
    .in(_U1367_in),
    .clk(_U1367_clk),
    .out(_U1367_out)
);
assign _U1368_in = _U1367_out;
assign _U1368_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1368 (
    .in(_U1368_in),
    .clk(_U1368_clk),
    .out(_U1368_out)
);
assign _U1369_in = _U1368_out;
assign _U1369_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1369 (
    .in(_U1369_in),
    .clk(_U1369_clk),
    .out(_U1369_out)
);
assign _U1370_in = _U1375_out;
_U1370_pt__U1371 _U1370 (
    .in(_U1370_in),
    .out(_U1370_out)
);
assign _U1372_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U1372_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1372 (
    .in(_U1372_in),
    .clk(_U1372_clk),
    .out(_U1372_out)
);
assign _U1373_in = _U1372_out;
assign _U1373_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1373 (
    .in(_U1373_in),
    .clk(_U1373_clk),
    .out(_U1373_out)
);
assign _U1374_in = _U1373_out;
assign _U1374_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1374 (
    .in(_U1374_in),
    .clk(_U1374_clk),
    .out(_U1374_out)
);
assign _U1375_in = _U1374_out;
assign _U1375_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1375 (
    .in(_U1375_in),
    .clk(_U1375_clk),
    .out(_U1375_out)
);
assign _U1376_in = _U1381_out;
_U1376_pt__U1377 _U1376 (
    .in(_U1376_in),
    .out(_U1376_out)
);
assign _U1378_in = in1_hw_input_global_wrapper_stencil[6];
assign _U1378_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1378 (
    .in(_U1378_in),
    .clk(_U1378_clk),
    .out(_U1378_out)
);
assign _U1379_in = _U1378_out;
assign _U1379_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1379 (
    .in(_U1379_in),
    .clk(_U1379_clk),
    .out(_U1379_out)
);
assign _U1380_in = _U1379_out;
assign _U1380_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1380 (
    .in(_U1380_in),
    .clk(_U1380_clk),
    .out(_U1380_out)
);
assign _U1381_in = _U1380_out;
assign _U1381_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1381 (
    .in(_U1381_in),
    .clk(_U1381_clk),
    .out(_U1381_out)
);
assign _U1382_in = _U1384_out;
_U1382_pt__U1383 _U1382 (
    .in(_U1382_in),
    .out(_U1382_out)
);
assign _U1384_in = 16'(_U1272_out + _U1250_out);
assign _U1384_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1384 (
    .in(_U1384_in),
    .clk(_U1384_clk),
    .out(_U1384_out)
);
assign _U1385_in = _U1398_out;
_U1385_pt__U1386 _U1385 (
    .in(_U1385_in),
    .out(_U1385_out)
);
assign _U1387_in = 16'(_U1240_out * _U1344_out);
assign _U1387_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1387 (
    .in(_U1387_in),
    .clk(_U1387_clk),
    .out(_U1387_out)
);
assign _U1388_in = _U1387_out;
assign _U1388_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1388 (
    .in(_U1388_in),
    .clk(_U1388_clk),
    .out(_U1388_out)
);
assign _U1389_in = _U1388_out;
assign _U1389_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1389 (
    .in(_U1389_in),
    .clk(_U1389_clk),
    .out(_U1389_out)
);
assign _U1390_in = _U1389_out;
assign _U1390_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1390 (
    .in(_U1390_in),
    .clk(_U1390_clk),
    .out(_U1390_out)
);
assign _U1391_in = _U1390_out;
assign _U1391_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1391 (
    .in(_U1391_in),
    .clk(_U1391_clk),
    .out(_U1391_out)
);
assign _U1392_in = _U1391_out;
assign _U1392_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1392 (
    .in(_U1392_in),
    .clk(_U1392_clk),
    .out(_U1392_out)
);
assign _U1393_in = _U1392_out;
assign _U1393_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1393 (
    .in(_U1393_in),
    .clk(_U1393_clk),
    .out(_U1393_out)
);
assign _U1394_in = _U1393_out;
assign _U1394_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1394 (
    .in(_U1394_in),
    .clk(_U1394_clk),
    .out(_U1394_out)
);
assign _U1395_in = _U1394_out;
assign _U1395_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1395 (
    .in(_U1395_in),
    .clk(_U1395_clk),
    .out(_U1395_out)
);
assign _U1396_in = _U1395_out;
assign _U1396_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1396 (
    .in(_U1396_in),
    .clk(_U1396_clk),
    .out(_U1396_out)
);
assign _U1397_in = _U1396_out;
assign _U1397_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1397 (
    .in(_U1397_in),
    .clk(_U1397_clk),
    .out(_U1397_out)
);
assign _U1398_in = _U1397_out;
assign _U1398_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1398 (
    .in(_U1398_in),
    .clk(_U1398_clk),
    .out(_U1398_out)
);
assign _U1399_in = _U1401_out;
_U1399_pt__U1400 _U1399 (
    .in(_U1399_in),
    .out(_U1399_out)
);
assign _U1401_in = 16'(_U1402_out + _U1414_out);
assign _U1401_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1401 (
    .in(_U1401_in),
    .clk(_U1401_clk),
    .out(_U1401_out)
);
assign _U1402_in = _U1413_out;
_U1402_pt__U1403 _U1402 (
    .in(_U1402_in),
    .out(_U1402_out)
);
assign _U1404_in = 16'(_U1346_out * _U1349_out);
assign _U1404_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1404 (
    .in(_U1404_in),
    .clk(_U1404_clk),
    .out(_U1404_out)
);
assign _U1405_in = _U1404_out;
assign _U1405_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1405 (
    .in(_U1405_in),
    .clk(_U1405_clk),
    .out(_U1405_out)
);
assign _U1406_in = _U1405_out;
assign _U1406_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1406 (
    .in(_U1406_in),
    .clk(_U1406_clk),
    .out(_U1406_out)
);
assign _U1407_in = _U1406_out;
assign _U1407_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1407 (
    .in(_U1407_in),
    .clk(_U1407_clk),
    .out(_U1407_out)
);
assign _U1408_in = _U1407_out;
assign _U1408_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1408 (
    .in(_U1408_in),
    .clk(_U1408_clk),
    .out(_U1408_out)
);
assign _U1409_in = _U1408_out;
assign _U1409_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1409 (
    .in(_U1409_in),
    .clk(_U1409_clk),
    .out(_U1409_out)
);
assign _U1410_in = _U1409_out;
assign _U1410_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1410 (
    .in(_U1410_in),
    .clk(_U1410_clk),
    .out(_U1410_out)
);
assign _U1411_in = _U1410_out;
assign _U1411_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1411 (
    .in(_U1411_in),
    .clk(_U1411_clk),
    .out(_U1411_out)
);
assign _U1412_in = _U1411_out;
assign _U1412_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1412 (
    .in(_U1412_in),
    .clk(_U1412_clk),
    .out(_U1412_out)
);
assign _U1413_in = _U1412_out;
assign _U1413_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1413 (
    .in(_U1413_in),
    .clk(_U1413_clk),
    .out(_U1413_out)
);
assign _U1414_in = _U1416_out;
_U1414_pt__U1415 _U1414 (
    .in(_U1414_in),
    .out(_U1414_out)
);
assign _U1416_in = 16'(_U1417_out + _U1427_out);
assign _U1416_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1416 (
    .in(_U1416_in),
    .clk(_U1416_clk),
    .out(_U1416_out)
);
assign _U1417_in = _U1426_out;
_U1417_pt__U1418 _U1417 (
    .in(_U1417_in),
    .out(_U1417_out)
);
assign _U1419_in = 16'(_U1352_out * _U1356_out);
assign _U1419_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1419 (
    .in(_U1419_in),
    .clk(_U1419_clk),
    .out(_U1419_out)
);
assign _U1420_in = _U1419_out;
assign _U1420_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1420 (
    .in(_U1420_in),
    .clk(_U1420_clk),
    .out(_U1420_out)
);
assign _U1421_in = _U1420_out;
assign _U1421_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1421 (
    .in(_U1421_in),
    .clk(_U1421_clk),
    .out(_U1421_out)
);
assign _U1422_in = _U1421_out;
assign _U1422_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1422 (
    .in(_U1422_in),
    .clk(_U1422_clk),
    .out(_U1422_out)
);
assign _U1423_in = _U1422_out;
assign _U1423_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1423 (
    .in(_U1423_in),
    .clk(_U1423_clk),
    .out(_U1423_out)
);
assign _U1424_in = _U1423_out;
assign _U1424_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1424 (
    .in(_U1424_in),
    .clk(_U1424_clk),
    .out(_U1424_out)
);
assign _U1425_in = _U1424_out;
assign _U1425_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1425 (
    .in(_U1425_in),
    .clk(_U1425_clk),
    .out(_U1425_out)
);
assign _U1426_in = _U1425_out;
assign _U1426_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1426 (
    .in(_U1426_in),
    .clk(_U1426_clk),
    .out(_U1426_out)
);
assign _U1427_in = _U1429_out;
_U1427_pt__U1428 _U1427 (
    .in(_U1427_in),
    .out(_U1427_out)
);
assign _U1429_in = 16'(_U1242_out + _U1280_out);
assign _U1429_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1429 (
    .in(_U1429_in),
    .clk(_U1429_clk),
    .out(_U1429_out)
);
assign _U1430_in = _U1440_out;
_U1430_pt__U1431 _U1430 (
    .in(_U1430_in),
    .out(_U1430_out)
);
assign _U1432_in = 16'(_U1310_out * _U1318_out);
assign _U1432_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1432 (
    .in(_U1432_in),
    .clk(_U1432_clk),
    .out(_U1432_out)
);
assign _U1433_in = _U1432_out;
assign _U1433_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1433 (
    .in(_U1433_in),
    .clk(_U1433_clk),
    .out(_U1433_out)
);
assign _U1434_in = _U1433_out;
assign _U1434_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1434 (
    .in(_U1434_in),
    .clk(_U1434_clk),
    .out(_U1434_out)
);
assign _U1435_in = _U1434_out;
assign _U1435_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1435 (
    .in(_U1435_in),
    .clk(_U1435_clk),
    .out(_U1435_out)
);
assign _U1436_in = _U1435_out;
assign _U1436_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1436 (
    .in(_U1436_in),
    .clk(_U1436_clk),
    .out(_U1436_out)
);
assign _U1437_in = _U1436_out;
assign _U1437_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1437 (
    .in(_U1437_in),
    .clk(_U1437_clk),
    .out(_U1437_out)
);
assign _U1438_in = _U1437_out;
assign _U1438_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1438 (
    .in(_U1438_in),
    .clk(_U1438_clk),
    .out(_U1438_out)
);
assign _U1439_in = _U1438_out;
assign _U1439_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1439 (
    .in(_U1439_in),
    .clk(_U1439_clk),
    .out(_U1439_out)
);
assign _U1440_in = _U1439_out;
assign _U1440_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1440 (
    .in(_U1440_in),
    .clk(_U1440_clk),
    .out(_U1440_out)
);
endmodule

module cu_op_hcompute_conv_stencil_14 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_14_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_14_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_14_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[0];
hcompute_conv_stencil_14_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_14_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U1232_pt__U1233 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1229_pt__U1230 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U121_pt__U122 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1219_pt__U1220 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1216_pt__U1217 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1204_pt__U1205 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1199_pt__U1200 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1195_pt__U1196 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1191_pt__U1192 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1188_pt__U1189 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1185_pt__U1186 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1183_pt__U1184 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1181_pt__U1182 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1172_pt__U1173 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1163_pt__U1164 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1155_pt__U1156 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1147_pt__U1148 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1140_pt__U1141 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1138_pt__U1139 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1135_pt__U1136 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1132_pt__U1133 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U112_pt__U113 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1126_pt__U1127 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1123_pt__U1124 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1115_pt__U1116 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1112_pt__U1113 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1109_pt__U1110 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1102_pt__U1103 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U10_pt__U11 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_5_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
wire [15:0] _U10_in;
assign _U10_in = in0_hw_input_stencil[0];
_U10_pt__U11 _U10 (
    .in(_U10_in),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil_5 (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read[0];
hcompute_hw_input_global_wrapper_stencil_5_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U1096_pt__U1097 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1090_pt__U1091 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1074_pt__U1075 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1067_pt__U1068 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1054_pt__U1055 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1049_pt__U1050 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U103_pt__U104 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_8_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U100_in;
wire _U100_clk;
wire [15:0] _U100_out;
wire [15:0] _U101_in;
wire _U101_clk;
wire [15:0] _U101_out;
wire [15:0] _U102_in;
wire _U102_clk;
wire [15:0] _U102_out;
wire [15:0] _U103_in;
wire [15:0] _U103_out;
wire [15:0] _U105_in;
wire _U105_clk;
wire [15:0] _U105_out;
wire [15:0] _U106_in;
wire _U106_clk;
wire [15:0] _U106_out;
wire [15:0] _U107_in;
wire _U107_clk;
wire [15:0] _U107_out;
wire [15:0] _U108_in;
wire _U108_clk;
wire [15:0] _U108_out;
wire [15:0] _U109_in;
wire _U109_clk;
wire [15:0] _U109_out;
wire [15:0] _U110_in;
wire _U110_clk;
wire [15:0] _U110_out;
wire [15:0] _U111_in;
wire _U111_clk;
wire [15:0] _U111_out;
wire [15:0] _U112_in;
wire [15:0] _U112_out;
wire [15:0] _U114_in;
wire _U114_clk;
wire [15:0] _U114_out;
wire [15:0] _U115_in;
wire _U115_clk;
wire [15:0] _U115_out;
wire [15:0] _U116_in;
wire _U116_clk;
wire [15:0] _U116_out;
wire [15:0] _U117_in;
wire _U117_clk;
wire [15:0] _U117_out;
wire [15:0] _U118_in;
wire _U118_clk;
wire [15:0] _U118_out;
wire [15:0] _U119_in;
wire _U119_clk;
wire [15:0] _U119_out;
wire [15:0] _U120_in;
wire _U120_clk;
wire [15:0] _U120_out;
wire [15:0] _U121_in;
wire [15:0] _U121_out;
wire [15:0] _U123_in;
wire _U123_clk;
wire [15:0] _U123_out;
wire [15:0] _U124_in;
wire _U124_clk;
wire [15:0] _U124_out;
wire [15:0] _U125_in;
wire _U125_clk;
wire [15:0] _U125_out;
wire [15:0] _U126_in;
wire _U126_clk;
wire [15:0] _U126_out;
wire [15:0] _U127_in;
wire _U127_clk;
wire [15:0] _U127_out;
wire [15:0] _U128_in;
wire _U128_clk;
wire [15:0] _U128_out;
wire [15:0] _U129_in;
wire _U129_clk;
wire [15:0] _U129_out;
wire [15:0] _U130_in;
wire _U130_clk;
wire [15:0] _U130_out;
wire [15:0] _U131_in;
wire _U131_clk;
wire [15:0] _U131_out;
wire [15:0] _U132_in;
wire _U132_clk;
wire [15:0] _U132_out;
wire [15:0] _U133_in;
wire _U133_clk;
wire [15:0] _U133_out;
wire [15:0] _U134_in;
wire _U134_clk;
wire [15:0] _U134_out;
wire [15:0] _U135_in;
wire _U135_clk;
wire [15:0] _U135_out;
wire [15:0] _U136_in;
wire _U136_clk;
wire [15:0] _U136_out;
wire [15:0] _U137_in;
wire _U137_clk;
wire [15:0] _U137_out;
wire [15:0] _U138_in;
wire [15:0] _U138_out;
wire [15:0] _U140_in;
wire _U140_clk;
wire [15:0] _U140_out;
wire [15:0] _U141_in;
wire [15:0] _U143_in;
wire [15:0] _U143_out;
wire [15:0] _U145_in;
wire _U145_clk;
wire [15:0] _U145_out;
wire [15:0] _U146_in;
wire _U146_clk;
wire [15:0] _U146_out;
wire [15:0] _U147_in;
wire _U147_clk;
wire [15:0] _U147_out;
wire [15:0] _U148_in;
wire _U148_clk;
wire [15:0] _U148_out;
wire [15:0] _U149_in;
wire _U149_clk;
wire [15:0] _U149_out;
wire [15:0] _U150_in;
wire _U150_clk;
wire [15:0] _U150_out;
wire [15:0] _U151_in;
wire _U151_clk;
wire [15:0] _U151_out;
wire [15:0] _U152_in;
wire _U152_clk;
wire [15:0] _U152_out;
wire [15:0] _U153_in;
wire _U153_clk;
wire [15:0] _U153_out;
wire [15:0] _U154_in;
wire _U154_clk;
wire [15:0] _U154_out;
wire [15:0] _U155_in;
wire _U155_clk;
wire [15:0] _U155_out;
wire [15:0] _U156_in;
wire _U156_clk;
wire [15:0] _U156_out;
wire [15:0] _U157_in;
wire [15:0] _U157_out;
wire [15:0] _U159_in;
wire _U159_clk;
wire [15:0] _U159_out;
wire [15:0] _U160_in;
wire [15:0] _U160_out;
wire [15:0] _U162_in;
wire _U162_clk;
wire [15:0] _U162_out;
wire [15:0] _U163_in;
wire _U163_clk;
wire [15:0] _U163_out;
wire [15:0] _U164_in;
wire _U164_clk;
wire [15:0] _U164_out;
wire [15:0] _U165_in;
wire _U165_clk;
wire [15:0] _U165_out;
wire [15:0] _U166_in;
wire _U166_clk;
wire [15:0] _U166_out;
wire [15:0] _U167_in;
wire _U167_clk;
wire [15:0] _U167_out;
wire [15:0] _U168_in;
wire _U168_clk;
wire [15:0] _U168_out;
wire [15:0] _U169_in;
wire _U169_clk;
wire [15:0] _U169_out;
wire [15:0] _U170_in;
wire _U170_clk;
wire [15:0] _U170_out;
wire [15:0] _U171_in;
wire _U171_clk;
wire [15:0] _U171_out;
wire [15:0] _U172_in;
wire [15:0] _U172_out;
wire [15:0] _U174_in;
wire _U174_clk;
wire [15:0] _U174_out;
wire [15:0] _U175_in;
wire [15:0] _U175_out;
wire [15:0] _U177_in;
wire _U177_clk;
wire [15:0] _U177_out;
wire [15:0] _U178_in;
wire _U178_clk;
wire [15:0] _U178_out;
wire [15:0] _U179_in;
wire _U179_clk;
wire [15:0] _U179_out;
wire [15:0] _U180_in;
wire _U180_clk;
wire [15:0] _U180_out;
wire [15:0] _U181_in;
wire _U181_clk;
wire [15:0] _U181_out;
wire [15:0] _U182_in;
wire _U182_clk;
wire [15:0] _U182_out;
wire [15:0] _U183_in;
wire _U183_clk;
wire [15:0] _U183_out;
wire [15:0] _U184_in;
wire _U184_clk;
wire [15:0] _U184_out;
wire [15:0] _U185_in;
wire [15:0] _U185_out;
wire [15:0] _U187_in;
wire _U187_clk;
wire [15:0] _U187_out;
wire [15:0] _U188_in;
wire [15:0] _U188_out;
wire [15:0] _U190_in;
wire _U190_clk;
wire [15:0] _U190_out;
wire [15:0] _U191_in;
wire _U191_clk;
wire [15:0] _U191_out;
wire [15:0] _U192_in;
wire _U192_clk;
wire [15:0] _U192_out;
wire [15:0] _U193_in;
wire _U193_clk;
wire [15:0] _U193_out;
wire [15:0] _U194_in;
wire _U194_clk;
wire [15:0] _U194_out;
wire [15:0] _U195_in;
wire _U195_clk;
wire [15:0] _U195_out;
wire [15:0] _U196_in;
wire [15:0] _U196_out;
wire [15:0] _U198_in;
wire _U198_clk;
wire [15:0] _U198_out;
wire [15:0] _U199_in;
wire [15:0] _U199_out;
wire [15:0] _U201_in;
wire _U201_clk;
wire [15:0] _U201_out;
wire [15:0] _U202_in;
wire _U202_clk;
wire [15:0] _U202_out;
wire [15:0] _U203_in;
wire _U203_clk;
wire [15:0] _U203_out;
wire [15:0] _U204_in;
wire _U204_clk;
wire [15:0] _U204_out;
wire [15:0] _U205_in;
wire [15:0] _U205_out;
wire [15:0] _U207_in;
wire _U207_clk;
wire [15:0] _U207_out;
wire [15:0] _U208_in;
wire [15:0] _U208_out;
wire [15:0] _U210_in;
wire _U210_clk;
wire [15:0] _U210_out;
wire [15:0] _U211_in;
wire _U211_clk;
wire [15:0] _U211_out;
wire [15:0] _U212_in;
wire [15:0] _U212_out;
wire [15:0] _U214_in;
wire _U214_clk;
wire [15:0] _U214_out;
wire [15:0] _U215_in;
wire [15:0] _U215_out;
wire [15:0] _U217_in;
wire _U217_clk;
wire [15:0] _U217_out;
wire [15:0] _U218_in;
wire _U218_clk;
wire [15:0] _U218_out;
wire [15:0] _U219_in;
wire _U219_clk;
wire [15:0] _U219_out;
wire [15:0] _U220_in;
wire _U220_clk;
wire [15:0] _U220_out;
wire [15:0] _U221_in;
wire _U221_clk;
wire [15:0] _U221_out;
wire [15:0] _U222_in;
wire _U222_clk;
wire [15:0] _U222_out;
wire [15:0] _U223_in;
wire _U223_clk;
wire [15:0] _U223_out;
wire [15:0] _U224_in;
wire _U224_clk;
wire [15:0] _U224_out;
wire [15:0] _U225_in;
wire _U225_clk;
wire [15:0] _U225_out;
wire [15:0] _U226_in;
wire _U226_clk;
wire [15:0] _U226_out;
wire [15:0] _U227_in;
wire _U227_clk;
wire [15:0] _U227_out;
wire [15:0] _U228_in;
wire _U228_clk;
wire [15:0] _U228_out;
wire [15:0] _U229_in;
wire _U229_clk;
wire [15:0] _U229_out;
wire [15:0] _U230_in;
wire _U230_clk;
wire [15:0] _U230_out;
wire [15:0] _U231_in;
wire [15:0] _U231_out;
wire [15:0] _U233_in;
wire [15:0] _U233_out;
wire [15:0] _U34_in;
wire [15:0] _U34_out;
wire [15:0] _U36_in;
wire _U36_clk;
wire [15:0] _U36_out;
wire [15:0] _U37_in;
wire [15:0] _U37_out;
wire [15:0] _U39_in;
wire _U39_clk;
wire [15:0] _U39_out;
wire [15:0] _U40_in;
wire [15:0] _U40_out;
wire [15:0] _U42_in;
wire _U42_clk;
wire [15:0] _U42_out;
wire [15:0] _U43_in;
wire [15:0] _U43_out;
wire [15:0] _U45_in;
wire _U45_clk;
wire [15:0] _U45_out;
wire [15:0] _U46_in;
wire _U46_clk;
wire [15:0] _U46_out;
wire [15:0] _U47_in;
wire [15:0] _U47_out;
wire [15:0] _U49_in;
wire _U49_clk;
wire [15:0] _U49_out;
wire [15:0] _U50_in;
wire _U50_clk;
wire [15:0] _U50_out;
wire [15:0] _U51_in;
wire [15:0] _U51_out;
wire [15:0] _U53_in;
wire _U53_clk;
wire [15:0] _U53_out;
wire [15:0] _U54_in;
wire _U54_clk;
wire [15:0] _U54_out;
wire [15:0] _U55_in;
wire _U55_clk;
wire [15:0] _U55_out;
wire [15:0] _U56_in;
wire [15:0] _U56_out;
wire [15:0] _U58_in;
wire _U58_clk;
wire [15:0] _U58_out;
wire [15:0] _U59_in;
wire _U59_clk;
wire [15:0] _U59_out;
wire [15:0] _U60_in;
wire _U60_clk;
wire [15:0] _U60_out;
wire [15:0] _U61_in;
wire [15:0] _U61_out;
wire [15:0] _U63_in;
wire _U63_clk;
wire [15:0] _U63_out;
wire [15:0] _U64_in;
wire _U64_clk;
wire [15:0] _U64_out;
wire [15:0] _U65_in;
wire _U65_clk;
wire [15:0] _U65_out;
wire [15:0] _U66_in;
wire _U66_clk;
wire [15:0] _U66_out;
wire [15:0] _U67_in;
wire [15:0] _U67_out;
wire [15:0] _U69_in;
wire _U69_clk;
wire [15:0] _U69_out;
wire [15:0] _U70_in;
wire _U70_clk;
wire [15:0] _U70_out;
wire [15:0] _U71_in;
wire _U71_clk;
wire [15:0] _U71_out;
wire [15:0] _U72_in;
wire _U72_clk;
wire [15:0] _U72_out;
wire [15:0] _U73_in;
wire [15:0] _U73_out;
wire [15:0] _U75_in;
wire _U75_clk;
wire [15:0] _U75_out;
wire [15:0] _U76_in;
wire _U76_clk;
wire [15:0] _U76_out;
wire [15:0] _U77_in;
wire _U77_clk;
wire [15:0] _U77_out;
wire [15:0] _U78_in;
wire _U78_clk;
wire [15:0] _U78_out;
wire [15:0] _U79_in;
wire _U79_clk;
wire [15:0] _U79_out;
wire [15:0] _U80_in;
wire [15:0] _U80_out;
wire [15:0] _U82_in;
wire _U82_clk;
wire [15:0] _U82_out;
wire [15:0] _U83_in;
wire _U83_clk;
wire [15:0] _U83_out;
wire [15:0] _U84_in;
wire _U84_clk;
wire [15:0] _U84_out;
wire [15:0] _U85_in;
wire _U85_clk;
wire [15:0] _U85_out;
wire [15:0] _U86_in;
wire _U86_clk;
wire [15:0] _U86_out;
wire [15:0] _U87_in;
wire [15:0] _U87_out;
wire [15:0] _U89_in;
wire _U89_clk;
wire [15:0] _U89_out;
wire [15:0] _U90_in;
wire _U90_clk;
wire [15:0] _U90_out;
wire [15:0] _U91_in;
wire _U91_clk;
wire [15:0] _U91_out;
wire [15:0] _U92_in;
wire _U92_clk;
wire [15:0] _U92_out;
wire [15:0] _U93_in;
wire _U93_clk;
wire [15:0] _U93_out;
wire [15:0] _U94_in;
wire _U94_clk;
wire [15:0] _U94_out;
wire [15:0] _U95_in;
wire [15:0] _U95_out;
wire [15:0] _U97_in;
wire _U97_clk;
wire [15:0] _U97_out;
wire [15:0] _U98_in;
wire _U98_clk;
wire [15:0] _U98_out;
wire [15:0] _U99_in;
wire _U99_clk;
wire [15:0] _U99_out;
assign _U100_in = _U99_out;
assign _U100_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U100 (
    .in(_U100_in),
    .clk(_U100_clk),
    .out(_U100_out)
);
assign _U101_in = _U100_out;
assign _U101_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U101 (
    .in(_U101_in),
    .clk(_U101_clk),
    .out(_U101_out)
);
assign _U102_in = _U101_out;
assign _U102_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U102 (
    .in(_U102_in),
    .clk(_U102_clk),
    .out(_U102_out)
);
assign _U103_in = _U111_out;
_U103_pt__U104 _U103 (
    .in(_U103_in),
    .out(_U103_out)
);
assign _U105_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U105_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U105 (
    .in(_U105_in),
    .clk(_U105_clk),
    .out(_U105_out)
);
assign _U106_in = _U105_out;
assign _U106_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U106 (
    .in(_U106_in),
    .clk(_U106_clk),
    .out(_U106_out)
);
assign _U107_in = _U106_out;
assign _U107_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U107 (
    .in(_U107_in),
    .clk(_U107_clk),
    .out(_U107_out)
);
assign _U108_in = _U107_out;
assign _U108_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U108 (
    .in(_U108_in),
    .clk(_U108_clk),
    .out(_U108_out)
);
assign _U109_in = _U108_out;
assign _U109_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U109 (
    .in(_U109_in),
    .clk(_U109_clk),
    .out(_U109_out)
);
assign _U110_in = _U109_out;
assign _U110_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U110 (
    .in(_U110_in),
    .clk(_U110_clk),
    .out(_U110_out)
);
assign _U111_in = _U110_out;
assign _U111_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U111 (
    .in(_U111_in),
    .clk(_U111_clk),
    .out(_U111_out)
);
assign _U112_in = _U120_out;
_U112_pt__U113 _U112 (
    .in(_U112_in),
    .out(_U112_out)
);
assign _U114_in = in1_hw_input_global_wrapper_stencil[7];
assign _U114_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U114 (
    .in(_U114_in),
    .clk(_U114_clk),
    .out(_U114_out)
);
assign _U115_in = _U114_out;
assign _U115_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U115 (
    .in(_U115_in),
    .clk(_U115_clk),
    .out(_U115_out)
);
assign _U116_in = _U115_out;
assign _U116_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U116 (
    .in(_U116_in),
    .clk(_U116_clk),
    .out(_U116_out)
);
assign _U117_in = _U116_out;
assign _U117_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U117 (
    .in(_U117_in),
    .clk(_U117_clk),
    .out(_U117_out)
);
assign _U118_in = _U117_out;
assign _U118_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U118 (
    .in(_U118_in),
    .clk(_U118_clk),
    .out(_U118_out)
);
assign _U119_in = _U118_out;
assign _U119_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U119 (
    .in(_U119_in),
    .clk(_U119_clk),
    .out(_U119_out)
);
assign _U120_in = _U119_out;
assign _U120_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U120 (
    .in(_U120_in),
    .clk(_U120_clk),
    .out(_U120_out)
);
assign _U121_in = _U137_out;
_U121_pt__U122 _U121 (
    .in(_U121_in),
    .out(_U121_out)
);
assign _U123_in = 16'(_U231_out * _U233_out);
assign _U123_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U123 (
    .in(_U123_in),
    .clk(_U123_clk),
    .out(_U123_out)
);
assign _U124_in = _U123_out;
assign _U124_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U124 (
    .in(_U124_in),
    .clk(_U124_clk),
    .out(_U124_out)
);
assign _U125_in = _U124_out;
assign _U125_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U125 (
    .in(_U125_in),
    .clk(_U125_clk),
    .out(_U125_out)
);
assign _U126_in = _U125_out;
assign _U126_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U126 (
    .in(_U126_in),
    .clk(_U126_clk),
    .out(_U126_out)
);
assign _U127_in = _U126_out;
assign _U127_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U127 (
    .in(_U127_in),
    .clk(_U127_clk),
    .out(_U127_out)
);
assign _U128_in = _U127_out;
assign _U128_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U128 (
    .in(_U128_in),
    .clk(_U128_clk),
    .out(_U128_out)
);
assign _U129_in = _U128_out;
assign _U129_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U129 (
    .in(_U129_in),
    .clk(_U129_clk),
    .out(_U129_out)
);
assign _U130_in = _U129_out;
assign _U130_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U130 (
    .in(_U130_in),
    .clk(_U130_clk),
    .out(_U130_out)
);
assign _U131_in = _U130_out;
assign _U131_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U131 (
    .in(_U131_in),
    .clk(_U131_clk),
    .out(_U131_out)
);
assign _U132_in = _U131_out;
assign _U132_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U132 (
    .in(_U132_in),
    .clk(_U132_clk),
    .out(_U132_out)
);
assign _U133_in = _U132_out;
assign _U133_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U133 (
    .in(_U133_in),
    .clk(_U133_clk),
    .out(_U133_out)
);
assign _U134_in = _U133_out;
assign _U134_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U134 (
    .in(_U134_in),
    .clk(_U134_clk),
    .out(_U134_out)
);
assign _U135_in = _U134_out;
assign _U135_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U135 (
    .in(_U135_in),
    .clk(_U135_clk),
    .out(_U135_out)
);
assign _U136_in = _U135_out;
assign _U136_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U136 (
    .in(_U136_in),
    .clk(_U136_clk),
    .out(_U136_out)
);
assign _U137_in = _U136_out;
assign _U137_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U137 (
    .in(_U137_in),
    .clk(_U137_clk),
    .out(_U137_out)
);
assign _U138_in = _U140_out;
_U138_pt__U139 _U138 (
    .in(_U138_in),
    .out(_U138_out)
);
assign _U140_in = 16'(_U215_out + _U34_out);
assign _U140_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U140 (
    .in(_U140_in),
    .clk(_U140_clk),
    .out(_U140_out)
);
assign _U141_in = 16'(_U121_out + _U138_out);
_U141_pt__U142 _U141 (
    .in(_U141_in),
    .out(out_conv_stencil)
);
assign _U143_in = _U156_out;
_U143_pt__U144 _U143 (
    .in(_U143_in),
    .out(_U143_out)
);
assign _U145_in = 16'(_U37_out * _U40_out);
assign _U145_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U145 (
    .in(_U145_in),
    .clk(_U145_clk),
    .out(_U145_out)
);
assign _U146_in = _U145_out;
assign _U146_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U146 (
    .in(_U146_in),
    .clk(_U146_clk),
    .out(_U146_out)
);
assign _U147_in = _U146_out;
assign _U147_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U147 (
    .in(_U147_in),
    .clk(_U147_clk),
    .out(_U147_out)
);
assign _U148_in = _U147_out;
assign _U148_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U148 (
    .in(_U148_in),
    .clk(_U148_clk),
    .out(_U148_out)
);
assign _U149_in = _U148_out;
assign _U149_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U149 (
    .in(_U149_in),
    .clk(_U149_clk),
    .out(_U149_out)
);
assign _U150_in = _U149_out;
assign _U150_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U150 (
    .in(_U150_in),
    .clk(_U150_clk),
    .out(_U150_out)
);
assign _U151_in = _U150_out;
assign _U151_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U151 (
    .in(_U151_in),
    .clk(_U151_clk),
    .out(_U151_out)
);
assign _U152_in = _U151_out;
assign _U152_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U152 (
    .in(_U152_in),
    .clk(_U152_clk),
    .out(_U152_out)
);
assign _U153_in = _U152_out;
assign _U153_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U153 (
    .in(_U153_in),
    .clk(_U153_clk),
    .out(_U153_out)
);
assign _U154_in = _U153_out;
assign _U154_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U154 (
    .in(_U154_in),
    .clk(_U154_clk),
    .out(_U154_out)
);
assign _U155_in = _U154_out;
assign _U155_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U155 (
    .in(_U155_in),
    .clk(_U155_clk),
    .out(_U155_out)
);
assign _U156_in = _U155_out;
assign _U156_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U156 (
    .in(_U156_in),
    .clk(_U156_clk),
    .out(_U156_out)
);
assign _U157_in = _U159_out;
_U157_pt__U158 _U157 (
    .in(_U157_in),
    .out(_U157_out)
);
assign _U159_in = 16'(_U160_out + _U172_out);
assign _U159_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U159 (
    .in(_U159_in),
    .clk(_U159_clk),
    .out(_U159_out)
);
assign _U160_in = _U171_out;
_U160_pt__U161 _U160 (
    .in(_U160_in),
    .out(_U160_out)
);
assign _U162_in = 16'(_U43_out * _U47_out);
assign _U162_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U162 (
    .in(_U162_in),
    .clk(_U162_clk),
    .out(_U162_out)
);
assign _U163_in = _U162_out;
assign _U163_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U163 (
    .in(_U163_in),
    .clk(_U163_clk),
    .out(_U163_out)
);
assign _U164_in = _U163_out;
assign _U164_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U164 (
    .in(_U164_in),
    .clk(_U164_clk),
    .out(_U164_out)
);
assign _U165_in = _U164_out;
assign _U165_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U165 (
    .in(_U165_in),
    .clk(_U165_clk),
    .out(_U165_out)
);
assign _U166_in = _U165_out;
assign _U166_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U166 (
    .in(_U166_in),
    .clk(_U166_clk),
    .out(_U166_out)
);
assign _U167_in = _U166_out;
assign _U167_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U167 (
    .in(_U167_in),
    .clk(_U167_clk),
    .out(_U167_out)
);
assign _U168_in = _U167_out;
assign _U168_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U168 (
    .in(_U168_in),
    .clk(_U168_clk),
    .out(_U168_out)
);
assign _U169_in = _U168_out;
assign _U169_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U169 (
    .in(_U169_in),
    .clk(_U169_clk),
    .out(_U169_out)
);
assign _U170_in = _U169_out;
assign _U170_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U170 (
    .in(_U170_in),
    .clk(_U170_clk),
    .out(_U170_out)
);
assign _U171_in = _U170_out;
assign _U171_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U171 (
    .in(_U171_in),
    .clk(_U171_clk),
    .out(_U171_out)
);
assign _U172_in = _U174_out;
_U172_pt__U173 _U172 (
    .in(_U172_in),
    .out(_U172_out)
);
assign _U174_in = 16'(_U175_out + _U185_out);
assign _U174_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U174 (
    .in(_U174_in),
    .clk(_U174_clk),
    .out(_U174_out)
);
assign _U175_in = _U184_out;
_U175_pt__U176 _U175 (
    .in(_U175_in),
    .out(_U175_out)
);
assign _U177_in = 16'(_U51_out * _U56_out);
assign _U177_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U177 (
    .in(_U177_in),
    .clk(_U177_clk),
    .out(_U177_out)
);
assign _U178_in = _U177_out;
assign _U178_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U178 (
    .in(_U178_in),
    .clk(_U178_clk),
    .out(_U178_out)
);
assign _U179_in = _U178_out;
assign _U179_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U179 (
    .in(_U179_in),
    .clk(_U179_clk),
    .out(_U179_out)
);
assign _U180_in = _U179_out;
assign _U180_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U180 (
    .in(_U180_in),
    .clk(_U180_clk),
    .out(_U180_out)
);
assign _U181_in = _U180_out;
assign _U181_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U181 (
    .in(_U181_in),
    .clk(_U181_clk),
    .out(_U181_out)
);
assign _U182_in = _U181_out;
assign _U182_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U182 (
    .in(_U182_in),
    .clk(_U182_clk),
    .out(_U182_out)
);
assign _U183_in = _U182_out;
assign _U183_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U183 (
    .in(_U183_in),
    .clk(_U183_clk),
    .out(_U183_out)
);
assign _U184_in = _U183_out;
assign _U184_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U184 (
    .in(_U184_in),
    .clk(_U184_clk),
    .out(_U184_out)
);
assign _U185_in = _U187_out;
_U185_pt__U186 _U185 (
    .in(_U185_in),
    .out(_U185_out)
);
assign _U187_in = 16'(_U188_out + _U196_out);
assign _U187_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U187 (
    .in(_U187_in),
    .clk(_U187_clk),
    .out(_U187_out)
);
assign _U188_in = _U195_out;
_U188_pt__U189 _U188 (
    .in(_U188_in),
    .out(_U188_out)
);
assign _U190_in = 16'(_U61_out * _U67_out);
assign _U190_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U190 (
    .in(_U190_in),
    .clk(_U190_clk),
    .out(_U190_out)
);
assign _U191_in = _U190_out;
assign _U191_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U191 (
    .in(_U191_in),
    .clk(_U191_clk),
    .out(_U191_out)
);
assign _U192_in = _U191_out;
assign _U192_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U192 (
    .in(_U192_in),
    .clk(_U192_clk),
    .out(_U192_out)
);
assign _U193_in = _U192_out;
assign _U193_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U193 (
    .in(_U193_in),
    .clk(_U193_clk),
    .out(_U193_out)
);
assign _U194_in = _U193_out;
assign _U194_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U194 (
    .in(_U194_in),
    .clk(_U194_clk),
    .out(_U194_out)
);
assign _U195_in = _U194_out;
assign _U195_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U195 (
    .in(_U195_in),
    .clk(_U195_clk),
    .out(_U195_out)
);
assign _U196_in = _U198_out;
_U196_pt__U197 _U196 (
    .in(_U196_in),
    .out(_U196_out)
);
assign _U198_in = 16'(_U199_out + _U205_out);
assign _U198_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U198 (
    .in(_U198_in),
    .clk(_U198_clk),
    .out(_U198_out)
);
assign _U199_in = _U204_out;
_U199_pt__U200 _U199 (
    .in(_U199_in),
    .out(_U199_out)
);
assign _U201_in = 16'(_U73_out * _U80_out);
assign _U201_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U201 (
    .in(_U201_in),
    .clk(_U201_clk),
    .out(_U201_out)
);
assign _U202_in = _U201_out;
assign _U202_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U202 (
    .in(_U202_in),
    .clk(_U202_clk),
    .out(_U202_out)
);
assign _U203_in = _U202_out;
assign _U203_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U203 (
    .in(_U203_in),
    .clk(_U203_clk),
    .out(_U203_out)
);
assign _U204_in = _U203_out;
assign _U204_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U204 (
    .in(_U204_in),
    .clk(_U204_clk),
    .out(_U204_out)
);
assign _U205_in = _U207_out;
_U205_pt__U206 _U205 (
    .in(_U205_in),
    .out(_U205_out)
);
assign _U207_in = 16'(_U208_out + _U212_out);
assign _U207_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U207 (
    .in(_U207_in),
    .clk(_U207_clk),
    .out(_U207_out)
);
assign _U208_in = _U211_out;
_U208_pt__U209 _U208 (
    .in(_U208_in),
    .out(_U208_out)
);
assign _U210_in = 16'(_U87_out * _U95_out);
assign _U210_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U210 (
    .in(_U210_in),
    .clk(_U210_clk),
    .out(_U210_out)
);
assign _U211_in = _U210_out;
assign _U211_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U211 (
    .in(_U211_in),
    .clk(_U211_clk),
    .out(_U211_out)
);
assign _U212_in = _U214_out;
_U212_pt__U213 _U212 (
    .in(_U212_in),
    .out(_U212_out)
);
assign _U214_in = 16'(_U103_out * _U112_out);
assign _U214_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U214 (
    .in(_U214_in),
    .clk(_U214_clk),
    .out(_U214_out)
);
assign _U215_in = _U230_out;
_U215_pt__U216 _U215 (
    .in(_U215_in),
    .out(_U215_out)
);
assign _U217_in = in0_conv_stencil[0];
assign _U217_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U217 (
    .in(_U217_in),
    .clk(_U217_clk),
    .out(_U217_out)
);
assign _U218_in = _U217_out;
assign _U218_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U218 (
    .in(_U218_in),
    .clk(_U218_clk),
    .out(_U218_out)
);
assign _U219_in = _U218_out;
assign _U219_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U219 (
    .in(_U219_in),
    .clk(_U219_clk),
    .out(_U219_out)
);
assign _U220_in = _U219_out;
assign _U220_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U220 (
    .in(_U220_in),
    .clk(_U220_clk),
    .out(_U220_out)
);
assign _U221_in = _U220_out;
assign _U221_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U221 (
    .in(_U221_in),
    .clk(_U221_clk),
    .out(_U221_out)
);
assign _U222_in = _U221_out;
assign _U222_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U222 (
    .in(_U222_in),
    .clk(_U222_clk),
    .out(_U222_out)
);
assign _U223_in = _U222_out;
assign _U223_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U223 (
    .in(_U223_in),
    .clk(_U223_clk),
    .out(_U223_out)
);
assign _U224_in = _U223_out;
assign _U224_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U224 (
    .in(_U224_in),
    .clk(_U224_clk),
    .out(_U224_out)
);
assign _U225_in = _U224_out;
assign _U225_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U225 (
    .in(_U225_in),
    .clk(_U225_clk),
    .out(_U225_out)
);
assign _U226_in = _U225_out;
assign _U226_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U226 (
    .in(_U226_in),
    .clk(_U226_clk),
    .out(_U226_out)
);
assign _U227_in = _U226_out;
assign _U227_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U227 (
    .in(_U227_in),
    .clk(_U227_clk),
    .out(_U227_out)
);
assign _U228_in = _U227_out;
assign _U228_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U228 (
    .in(_U228_in),
    .clk(_U228_clk),
    .out(_U228_out)
);
assign _U229_in = _U228_out;
assign _U229_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U229 (
    .in(_U229_in),
    .clk(_U229_clk),
    .out(_U229_out)
);
assign _U230_in = _U229_out;
assign _U230_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U230 (
    .in(_U230_in),
    .clk(_U230_clk),
    .out(_U230_out)
);
assign _U231_in = in2_hw_kernel_global_wrapper_stencil[0];
_U231_pt__U232 _U231 (
    .in(_U231_in),
    .out(_U231_out)
);
assign _U233_in = in1_hw_input_global_wrapper_stencil[0];
_U233_pt__U234 _U233 (
    .in(_U233_in),
    .out(_U233_out)
);
assign _U34_in = _U36_out;
_U34_pt__U35 _U34 (
    .in(_U34_in),
    .out(_U34_out)
);
assign _U36_in = 16'(_U143_out + _U157_out);
assign _U36_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U36 (
    .in(_U36_in),
    .clk(_U36_clk),
    .out(_U36_out)
);
assign _U37_in = _U39_out;
_U37_pt__U38 _U37 (
    .in(_U37_in),
    .out(_U37_out)
);
assign _U39_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U39_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U39 (
    .in(_U39_in),
    .clk(_U39_clk),
    .out(_U39_out)
);
assign _U40_in = _U42_out;
_U40_pt__U41 _U40 (
    .in(_U40_in),
    .out(_U40_out)
);
assign _U42_in = in1_hw_input_global_wrapper_stencil[1];
assign _U42_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U42 (
    .in(_U42_in),
    .clk(_U42_clk),
    .out(_U42_out)
);
assign _U43_in = _U46_out;
_U43_pt__U44 _U43 (
    .in(_U43_in),
    .out(_U43_out)
);
assign _U45_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U45_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U45 (
    .in(_U45_in),
    .clk(_U45_clk),
    .out(_U45_out)
);
assign _U46_in = _U45_out;
assign _U46_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U46 (
    .in(_U46_in),
    .clk(_U46_clk),
    .out(_U46_out)
);
assign _U47_in = _U50_out;
_U47_pt__U48 _U47 (
    .in(_U47_in),
    .out(_U47_out)
);
assign _U49_in = in1_hw_input_global_wrapper_stencil[2];
assign _U49_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U49 (
    .in(_U49_in),
    .clk(_U49_clk),
    .out(_U49_out)
);
assign _U50_in = _U49_out;
assign _U50_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U50 (
    .in(_U50_in),
    .clk(_U50_clk),
    .out(_U50_out)
);
assign _U51_in = _U55_out;
_U51_pt__U52 _U51 (
    .in(_U51_in),
    .out(_U51_out)
);
assign _U53_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U53_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U53 (
    .in(_U53_in),
    .clk(_U53_clk),
    .out(_U53_out)
);
assign _U54_in = _U53_out;
assign _U54_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U54 (
    .in(_U54_in),
    .clk(_U54_clk),
    .out(_U54_out)
);
assign _U55_in = _U54_out;
assign _U55_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U55 (
    .in(_U55_in),
    .clk(_U55_clk),
    .out(_U55_out)
);
assign _U56_in = _U60_out;
_U56_pt__U57 _U56 (
    .in(_U56_in),
    .out(_U56_out)
);
assign _U58_in = in1_hw_input_global_wrapper_stencil[3];
assign _U58_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U58 (
    .in(_U58_in),
    .clk(_U58_clk),
    .out(_U58_out)
);
assign _U59_in = _U58_out;
assign _U59_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U59 (
    .in(_U59_in),
    .clk(_U59_clk),
    .out(_U59_out)
);
assign _U60_in = _U59_out;
assign _U60_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U60 (
    .in(_U60_in),
    .clk(_U60_clk),
    .out(_U60_out)
);
assign _U61_in = _U66_out;
_U61_pt__U62 _U61 (
    .in(_U61_in),
    .out(_U61_out)
);
assign _U63_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U63_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U63 (
    .in(_U63_in),
    .clk(_U63_clk),
    .out(_U63_out)
);
assign _U64_in = _U63_out;
assign _U64_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U64 (
    .in(_U64_in),
    .clk(_U64_clk),
    .out(_U64_out)
);
assign _U65_in = _U64_out;
assign _U65_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U65 (
    .in(_U65_in),
    .clk(_U65_clk),
    .out(_U65_out)
);
assign _U66_in = _U65_out;
assign _U66_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U66 (
    .in(_U66_in),
    .clk(_U66_clk),
    .out(_U66_out)
);
assign _U67_in = _U72_out;
_U67_pt__U68 _U67 (
    .in(_U67_in),
    .out(_U67_out)
);
assign _U69_in = in1_hw_input_global_wrapper_stencil[4];
assign _U69_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U69 (
    .in(_U69_in),
    .clk(_U69_clk),
    .out(_U69_out)
);
assign _U70_in = _U69_out;
assign _U70_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U70 (
    .in(_U70_in),
    .clk(_U70_clk),
    .out(_U70_out)
);
assign _U71_in = _U70_out;
assign _U71_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U71 (
    .in(_U71_in),
    .clk(_U71_clk),
    .out(_U71_out)
);
assign _U72_in = _U71_out;
assign _U72_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U72 (
    .in(_U72_in),
    .clk(_U72_clk),
    .out(_U72_out)
);
assign _U73_in = _U79_out;
_U73_pt__U74 _U73 (
    .in(_U73_in),
    .out(_U73_out)
);
assign _U75_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U75_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U75 (
    .in(_U75_in),
    .clk(_U75_clk),
    .out(_U75_out)
);
assign _U76_in = _U75_out;
assign _U76_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U76 (
    .in(_U76_in),
    .clk(_U76_clk),
    .out(_U76_out)
);
assign _U77_in = _U76_out;
assign _U77_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U77 (
    .in(_U77_in),
    .clk(_U77_clk),
    .out(_U77_out)
);
assign _U78_in = _U77_out;
assign _U78_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U78 (
    .in(_U78_in),
    .clk(_U78_clk),
    .out(_U78_out)
);
assign _U79_in = _U78_out;
assign _U79_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U79 (
    .in(_U79_in),
    .clk(_U79_clk),
    .out(_U79_out)
);
assign _U80_in = _U86_out;
_U80_pt__U81 _U80 (
    .in(_U80_in),
    .out(_U80_out)
);
assign _U82_in = in1_hw_input_global_wrapper_stencil[5];
assign _U82_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U82 (
    .in(_U82_in),
    .clk(_U82_clk),
    .out(_U82_out)
);
assign _U83_in = _U82_out;
assign _U83_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U83 (
    .in(_U83_in),
    .clk(_U83_clk),
    .out(_U83_out)
);
assign _U84_in = _U83_out;
assign _U84_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U84 (
    .in(_U84_in),
    .clk(_U84_clk),
    .out(_U84_out)
);
assign _U85_in = _U84_out;
assign _U85_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U85 (
    .in(_U85_in),
    .clk(_U85_clk),
    .out(_U85_out)
);
assign _U86_in = _U85_out;
assign _U86_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U86 (
    .in(_U86_in),
    .clk(_U86_clk),
    .out(_U86_out)
);
assign _U87_in = _U94_out;
_U87_pt__U88 _U87 (
    .in(_U87_in),
    .out(_U87_out)
);
assign _U89_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U89_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U89 (
    .in(_U89_in),
    .clk(_U89_clk),
    .out(_U89_out)
);
assign _U90_in = _U89_out;
assign _U90_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U90 (
    .in(_U90_in),
    .clk(_U90_clk),
    .out(_U90_out)
);
assign _U91_in = _U90_out;
assign _U91_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U91 (
    .in(_U91_in),
    .clk(_U91_clk),
    .out(_U91_out)
);
assign _U92_in = _U91_out;
assign _U92_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U92 (
    .in(_U92_in),
    .clk(_U92_clk),
    .out(_U92_out)
);
assign _U93_in = _U92_out;
assign _U93_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U93 (
    .in(_U93_in),
    .clk(_U93_clk),
    .out(_U93_out)
);
assign _U94_in = _U93_out;
assign _U94_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U94 (
    .in(_U94_in),
    .clk(_U94_clk),
    .out(_U94_out)
);
assign _U95_in = _U102_out;
_U95_pt__U96 _U95 (
    .in(_U95_in),
    .out(_U95_out)
);
assign _U97_in = in1_hw_input_global_wrapper_stencil[6];
assign _U97_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U97 (
    .in(_U97_in),
    .clk(_U97_clk),
    .out(_U97_out)
);
assign _U98_in = _U97_out;
assign _U98_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U98 (
    .in(_U98_in),
    .clk(_U98_clk),
    .out(_U98_out)
);
assign _U99_in = _U98_out;
assign _U99_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U99 (
    .in(_U99_in),
    .clk(_U99_clk),
    .out(_U99_out)
);
endmodule

module cu_op_hcompute_conv_stencil_8 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_8_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_8_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_8_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[0];
hcompute_conv_stencil_8_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_8_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U1039_pt__U1040 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_13_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U1039_in;
wire [15:0] _U1039_out;
wire [15:0] _U1041_in;
wire _U1041_clk;
wire [15:0] _U1041_out;
wire [15:0] _U1042_in;
wire _U1042_clk;
wire [15:0] _U1042_out;
wire [15:0] _U1043_in;
wire _U1043_clk;
wire [15:0] _U1043_out;
wire [15:0] _U1044_in;
wire _U1044_clk;
wire [15:0] _U1044_out;
wire [15:0] _U1045_in;
wire _U1045_clk;
wire [15:0] _U1045_out;
wire [15:0] _U1046_in;
wire _U1046_clk;
wire [15:0] _U1046_out;
wire [15:0] _U1047_in;
wire _U1047_clk;
wire [15:0] _U1047_out;
wire [15:0] _U1048_in;
wire _U1048_clk;
wire [15:0] _U1048_out;
wire [15:0] _U1049_in;
wire [15:0] _U1049_out;
wire [15:0] _U1051_in;
wire _U1051_clk;
wire [15:0] _U1051_out;
wire [15:0] _U1052_in;
wire _U1052_clk;
wire [15:0] _U1052_out;
wire [15:0] _U1053_in;
wire _U1053_clk;
wire [15:0] _U1053_out;
wire [15:0] _U1054_in;
wire [15:0] _U1054_out;
wire [15:0] _U1056_in;
wire _U1056_clk;
wire [15:0] _U1056_out;
wire [15:0] _U1057_in;
wire _U1057_clk;
wire [15:0] _U1057_out;
wire [15:0] _U1058_in;
wire _U1058_clk;
wire [15:0] _U1058_out;
wire [15:0] _U1059_in;
wire _U1059_clk;
wire [15:0] _U1059_out;
wire [15:0] _U1060_in;
wire _U1060_clk;
wire [15:0] _U1060_out;
wire [15:0] _U1061_in;
wire _U1061_clk;
wire [15:0] _U1061_out;
wire [15:0] _U1062_in;
wire _U1062_clk;
wire [15:0] _U1062_out;
wire [15:0] _U1063_in;
wire _U1063_clk;
wire [15:0] _U1063_out;
wire [15:0] _U1064_in;
wire _U1064_clk;
wire [15:0] _U1064_out;
wire [15:0] _U1065_in;
wire _U1065_clk;
wire [15:0] _U1065_out;
wire [15:0] _U1066_in;
wire _U1066_clk;
wire [15:0] _U1066_out;
wire [15:0] _U1067_in;
wire [15:0] _U1067_out;
wire [15:0] _U1069_in;
wire _U1069_clk;
wire [15:0] _U1069_out;
wire [15:0] _U1070_in;
wire _U1070_clk;
wire [15:0] _U1070_out;
wire [15:0] _U1071_in;
wire _U1071_clk;
wire [15:0] _U1071_out;
wire [15:0] _U1072_in;
wire _U1072_clk;
wire [15:0] _U1072_out;
wire [15:0] _U1073_in;
wire _U1073_clk;
wire [15:0] _U1073_out;
wire [15:0] _U1074_in;
wire [15:0] _U1074_out;
wire [15:0] _U1076_in;
wire _U1076_clk;
wire [15:0] _U1076_out;
wire [15:0] _U1077_in;
wire _U1077_clk;
wire [15:0] _U1077_out;
wire [15:0] _U1078_in;
wire _U1078_clk;
wire [15:0] _U1078_out;
wire [15:0] _U1079_in;
wire _U1079_clk;
wire [15:0] _U1079_out;
wire [15:0] _U1080_in;
wire _U1080_clk;
wire [15:0] _U1080_out;
wire [15:0] _U1081_in;
wire _U1081_clk;
wire [15:0] _U1081_out;
wire [15:0] _U1082_in;
wire _U1082_clk;
wire [15:0] _U1082_out;
wire [15:0] _U1083_in;
wire _U1083_clk;
wire [15:0] _U1083_out;
wire [15:0] _U1084_in;
wire _U1084_clk;
wire [15:0] _U1084_out;
wire [15:0] _U1085_in;
wire _U1085_clk;
wire [15:0] _U1085_out;
wire [15:0] _U1086_in;
wire _U1086_clk;
wire [15:0] _U1086_out;
wire [15:0] _U1087_in;
wire _U1087_clk;
wire [15:0] _U1087_out;
wire [15:0] _U1088_in;
wire _U1088_clk;
wire [15:0] _U1088_out;
wire [15:0] _U1089_in;
wire _U1089_clk;
wire [15:0] _U1089_out;
wire [15:0] _U1090_in;
wire [15:0] _U1090_out;
wire [15:0] _U1092_in;
wire _U1092_clk;
wire [15:0] _U1092_out;
wire [15:0] _U1093_in;
wire _U1093_clk;
wire [15:0] _U1093_out;
wire [15:0] _U1094_in;
wire _U1094_clk;
wire [15:0] _U1094_out;
wire [15:0] _U1095_in;
wire _U1095_clk;
wire [15:0] _U1095_out;
wire [15:0] _U1096_in;
wire [15:0] _U1096_out;
wire [15:0] _U1098_in;
wire _U1098_clk;
wire [15:0] _U1098_out;
wire [15:0] _U1099_in;
wire _U1099_clk;
wire [15:0] _U1099_out;
wire [15:0] _U1100_in;
wire _U1100_clk;
wire [15:0] _U1100_out;
wire [15:0] _U1101_in;
wire _U1101_clk;
wire [15:0] _U1101_out;
wire [15:0] _U1102_in;
wire [15:0] _U1102_out;
wire [15:0] _U1104_in;
wire _U1104_clk;
wire [15:0] _U1104_out;
wire [15:0] _U1105_in;
wire _U1105_clk;
wire [15:0] _U1105_out;
wire [15:0] _U1106_in;
wire _U1106_clk;
wire [15:0] _U1106_out;
wire [15:0] _U1107_in;
wire _U1107_clk;
wire [15:0] _U1107_out;
wire [15:0] _U1108_in;
wire _U1108_clk;
wire [15:0] _U1108_out;
wire [15:0] _U1109_in;
wire [15:0] _U1109_out;
wire [15:0] _U1111_in;
wire _U1111_clk;
wire [15:0] _U1111_out;
wire [15:0] _U1112_in;
wire [15:0] _U1112_out;
wire [15:0] _U1114_in;
wire _U1114_clk;
wire [15:0] _U1114_out;
wire [15:0] _U1115_in;
wire [15:0] _U1115_out;
wire [15:0] _U1117_in;
wire _U1117_clk;
wire [15:0] _U1117_out;
wire [15:0] _U1118_in;
wire _U1118_clk;
wire [15:0] _U1118_out;
wire [15:0] _U1119_in;
wire _U1119_clk;
wire [15:0] _U1119_out;
wire [15:0] _U1120_in;
wire _U1120_clk;
wire [15:0] _U1120_out;
wire [15:0] _U1121_in;
wire _U1121_clk;
wire [15:0] _U1121_out;
wire [15:0] _U1122_in;
wire _U1122_clk;
wire [15:0] _U1122_out;
wire [15:0] _U1123_in;
wire [15:0] _U1123_out;
wire [15:0] _U1125_in;
wire _U1125_clk;
wire [15:0] _U1125_out;
wire [15:0] _U1126_in;
wire [15:0] _U1126_out;
wire [15:0] _U1128_in;
wire _U1128_clk;
wire [15:0] _U1128_out;
wire [15:0] _U1129_in;
wire _U1129_clk;
wire [15:0] _U1129_out;
wire [15:0] _U1130_in;
wire _U1130_clk;
wire [15:0] _U1130_out;
wire [15:0] _U1131_in;
wire _U1131_clk;
wire [15:0] _U1131_out;
wire [15:0] _U1132_in;
wire [15:0] _U1132_out;
wire [15:0] _U1134_in;
wire _U1134_clk;
wire [15:0] _U1134_out;
wire [15:0] _U1135_in;
wire [15:0] _U1135_out;
wire [15:0] _U1137_in;
wire _U1137_clk;
wire [15:0] _U1137_out;
wire [15:0] _U1138_in;
wire [15:0] _U1140_in;
wire [15:0] _U1140_out;
wire [15:0] _U1142_in;
wire _U1142_clk;
wire [15:0] _U1142_out;
wire [15:0] _U1143_in;
wire _U1143_clk;
wire [15:0] _U1143_out;
wire [15:0] _U1144_in;
wire _U1144_clk;
wire [15:0] _U1144_out;
wire [15:0] _U1145_in;
wire _U1145_clk;
wire [15:0] _U1145_out;
wire [15:0] _U1146_in;
wire _U1146_clk;
wire [15:0] _U1146_out;
wire [15:0] _U1147_in;
wire [15:0] _U1147_out;
wire [15:0] _U1149_in;
wire _U1149_clk;
wire [15:0] _U1149_out;
wire [15:0] _U1150_in;
wire _U1150_clk;
wire [15:0] _U1150_out;
wire [15:0] _U1151_in;
wire _U1151_clk;
wire [15:0] _U1151_out;
wire [15:0] _U1152_in;
wire _U1152_clk;
wire [15:0] _U1152_out;
wire [15:0] _U1153_in;
wire _U1153_clk;
wire [15:0] _U1153_out;
wire [15:0] _U1154_in;
wire _U1154_clk;
wire [15:0] _U1154_out;
wire [15:0] _U1155_in;
wire [15:0] _U1155_out;
wire [15:0] _U1157_in;
wire _U1157_clk;
wire [15:0] _U1157_out;
wire [15:0] _U1158_in;
wire _U1158_clk;
wire [15:0] _U1158_out;
wire [15:0] _U1159_in;
wire _U1159_clk;
wire [15:0] _U1159_out;
wire [15:0] _U1160_in;
wire _U1160_clk;
wire [15:0] _U1160_out;
wire [15:0] _U1161_in;
wire _U1161_clk;
wire [15:0] _U1161_out;
wire [15:0] _U1162_in;
wire _U1162_clk;
wire [15:0] _U1162_out;
wire [15:0] _U1163_in;
wire [15:0] _U1163_out;
wire [15:0] _U1165_in;
wire _U1165_clk;
wire [15:0] _U1165_out;
wire [15:0] _U1166_in;
wire _U1166_clk;
wire [15:0] _U1166_out;
wire [15:0] _U1167_in;
wire _U1167_clk;
wire [15:0] _U1167_out;
wire [15:0] _U1168_in;
wire _U1168_clk;
wire [15:0] _U1168_out;
wire [15:0] _U1169_in;
wire _U1169_clk;
wire [15:0] _U1169_out;
wire [15:0] _U1170_in;
wire _U1170_clk;
wire [15:0] _U1170_out;
wire [15:0] _U1171_in;
wire _U1171_clk;
wire [15:0] _U1171_out;
wire [15:0] _U1172_in;
wire [15:0] _U1172_out;
wire [15:0] _U1174_in;
wire _U1174_clk;
wire [15:0] _U1174_out;
wire [15:0] _U1175_in;
wire _U1175_clk;
wire [15:0] _U1175_out;
wire [15:0] _U1176_in;
wire _U1176_clk;
wire [15:0] _U1176_out;
wire [15:0] _U1177_in;
wire _U1177_clk;
wire [15:0] _U1177_out;
wire [15:0] _U1178_in;
wire _U1178_clk;
wire [15:0] _U1178_out;
wire [15:0] _U1179_in;
wire _U1179_clk;
wire [15:0] _U1179_out;
wire [15:0] _U1180_in;
wire _U1180_clk;
wire [15:0] _U1180_out;
wire [15:0] _U1181_in;
wire [15:0] _U1181_out;
wire [15:0] _U1183_in;
wire [15:0] _U1183_out;
wire [15:0] _U1185_in;
wire [15:0] _U1185_out;
wire [15:0] _U1187_in;
wire _U1187_clk;
wire [15:0] _U1187_out;
wire [15:0] _U1188_in;
wire [15:0] _U1188_out;
wire [15:0] _U1190_in;
wire _U1190_clk;
wire [15:0] _U1190_out;
wire [15:0] _U1191_in;
wire [15:0] _U1191_out;
wire [15:0] _U1193_in;
wire _U1193_clk;
wire [15:0] _U1193_out;
wire [15:0] _U1194_in;
wire _U1194_clk;
wire [15:0] _U1194_out;
wire [15:0] _U1195_in;
wire [15:0] _U1195_out;
wire [15:0] _U1197_in;
wire _U1197_clk;
wire [15:0] _U1197_out;
wire [15:0] _U1198_in;
wire _U1198_clk;
wire [15:0] _U1198_out;
wire [15:0] _U1199_in;
wire [15:0] _U1199_out;
wire [15:0] _U1201_in;
wire _U1201_clk;
wire [15:0] _U1201_out;
wire [15:0] _U1202_in;
wire _U1202_clk;
wire [15:0] _U1202_out;
wire [15:0] _U1203_in;
wire _U1203_clk;
wire [15:0] _U1203_out;
wire [15:0] _U1204_in;
wire [15:0] _U1204_out;
wire [15:0] _U1206_in;
wire _U1206_clk;
wire [15:0] _U1206_out;
wire [15:0] _U1207_in;
wire _U1207_clk;
wire [15:0] _U1207_out;
wire [15:0] _U1208_in;
wire _U1208_clk;
wire [15:0] _U1208_out;
wire [15:0] _U1209_in;
wire _U1209_clk;
wire [15:0] _U1209_out;
wire [15:0] _U1210_in;
wire _U1210_clk;
wire [15:0] _U1210_out;
wire [15:0] _U1211_in;
wire _U1211_clk;
wire [15:0] _U1211_out;
wire [15:0] _U1212_in;
wire _U1212_clk;
wire [15:0] _U1212_out;
wire [15:0] _U1213_in;
wire _U1213_clk;
wire [15:0] _U1213_out;
wire [15:0] _U1214_in;
wire _U1214_clk;
wire [15:0] _U1214_out;
wire [15:0] _U1215_in;
wire _U1215_clk;
wire [15:0] _U1215_out;
wire [15:0] _U1216_in;
wire [15:0] _U1216_out;
wire [15:0] _U1218_in;
wire _U1218_clk;
wire [15:0] _U1218_out;
wire [15:0] _U1219_in;
wire [15:0] _U1219_out;
wire [15:0] _U1221_in;
wire _U1221_clk;
wire [15:0] _U1221_out;
wire [15:0] _U1222_in;
wire _U1222_clk;
wire [15:0] _U1222_out;
wire [15:0] _U1223_in;
wire _U1223_clk;
wire [15:0] _U1223_out;
wire [15:0] _U1224_in;
wire _U1224_clk;
wire [15:0] _U1224_out;
wire [15:0] _U1225_in;
wire _U1225_clk;
wire [15:0] _U1225_out;
wire [15:0] _U1226_in;
wire _U1226_clk;
wire [15:0] _U1226_out;
wire [15:0] _U1227_in;
wire _U1227_clk;
wire [15:0] _U1227_out;
wire [15:0] _U1228_in;
wire _U1228_clk;
wire [15:0] _U1228_out;
wire [15:0] _U1229_in;
wire [15:0] _U1229_out;
wire [15:0] _U1231_in;
wire _U1231_clk;
wire [15:0] _U1231_out;
wire [15:0] _U1232_in;
wire [15:0] _U1232_out;
wire [15:0] _U1234_in;
wire _U1234_clk;
wire [15:0] _U1234_out;
wire [15:0] _U1235_in;
wire _U1235_clk;
wire [15:0] _U1235_out;
wire [15:0] _U1236_in;
wire _U1236_clk;
wire [15:0] _U1236_out;
wire [15:0] _U1237_in;
wire _U1237_clk;
wire [15:0] _U1237_out;
wire [15:0] _U1238_in;
wire _U1238_clk;
wire [15:0] _U1238_out;
wire [15:0] _U1239_in;
wire _U1239_clk;
wire [15:0] _U1239_out;
assign _U1039_in = _U1048_out;
_U1039_pt__U1040 _U1039 (
    .in(_U1039_in),
    .out(_U1039_out)
);
assign _U1041_in = 16'(_U1102_out * _U1140_out);
assign _U1041_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1041 (
    .in(_U1041_in),
    .clk(_U1041_clk),
    .out(_U1041_out)
);
assign _U1042_in = _U1041_out;
assign _U1042_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1042 (
    .in(_U1042_in),
    .clk(_U1042_clk),
    .out(_U1042_out)
);
assign _U1043_in = _U1042_out;
assign _U1043_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1043 (
    .in(_U1043_in),
    .clk(_U1043_clk),
    .out(_U1043_out)
);
assign _U1044_in = _U1043_out;
assign _U1044_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1044 (
    .in(_U1044_in),
    .clk(_U1044_clk),
    .out(_U1044_out)
);
assign _U1045_in = _U1044_out;
assign _U1045_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1045 (
    .in(_U1045_in),
    .clk(_U1045_clk),
    .out(_U1045_out)
);
assign _U1046_in = _U1045_out;
assign _U1046_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1046 (
    .in(_U1046_in),
    .clk(_U1046_clk),
    .out(_U1046_out)
);
assign _U1047_in = _U1046_out;
assign _U1047_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1047 (
    .in(_U1047_in),
    .clk(_U1047_clk),
    .out(_U1047_out)
);
assign _U1048_in = _U1047_out;
assign _U1048_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1048 (
    .in(_U1048_in),
    .clk(_U1048_clk),
    .out(_U1048_out)
);
assign _U1049_in = _U1053_out;
_U1049_pt__U1050 _U1049 (
    .in(_U1049_in),
    .out(_U1049_out)
);
assign _U1051_in = in1_hw_input_global_wrapper_stencil[7];
assign _U1051_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1051 (
    .in(_U1051_in),
    .clk(_U1051_clk),
    .out(_U1051_out)
);
assign _U1052_in = _U1051_out;
assign _U1052_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1052 (
    .in(_U1052_in),
    .clk(_U1052_clk),
    .out(_U1052_out)
);
assign _U1053_in = _U1052_out;
assign _U1053_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1053 (
    .in(_U1053_in),
    .clk(_U1053_clk),
    .out(_U1053_out)
);
assign _U1054_in = _U1066_out;
_U1054_pt__U1055 _U1054 (
    .in(_U1054_in),
    .out(_U1054_out)
);
assign _U1056_in = 16'(_U1090_out * _U1096_out);
assign _U1056_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1056 (
    .in(_U1056_in),
    .clk(_U1056_clk),
    .out(_U1056_out)
);
assign _U1057_in = _U1056_out;
assign _U1057_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1057 (
    .in(_U1057_in),
    .clk(_U1057_clk),
    .out(_U1057_out)
);
assign _U1058_in = _U1057_out;
assign _U1058_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1058 (
    .in(_U1058_in),
    .clk(_U1058_clk),
    .out(_U1058_out)
);
assign _U1059_in = _U1058_out;
assign _U1059_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1059 (
    .in(_U1059_in),
    .clk(_U1059_clk),
    .out(_U1059_out)
);
assign _U1060_in = _U1059_out;
assign _U1060_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1060 (
    .in(_U1060_in),
    .clk(_U1060_clk),
    .out(_U1060_out)
);
assign _U1061_in = _U1060_out;
assign _U1061_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1061 (
    .in(_U1061_in),
    .clk(_U1061_clk),
    .out(_U1061_out)
);
assign _U1062_in = _U1061_out;
assign _U1062_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1062 (
    .in(_U1062_in),
    .clk(_U1062_clk),
    .out(_U1062_out)
);
assign _U1063_in = _U1062_out;
assign _U1063_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1063 (
    .in(_U1063_in),
    .clk(_U1063_clk),
    .out(_U1063_out)
);
assign _U1064_in = _U1063_out;
assign _U1064_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1064 (
    .in(_U1064_in),
    .clk(_U1064_clk),
    .out(_U1064_out)
);
assign _U1065_in = _U1064_out;
assign _U1065_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1065 (
    .in(_U1065_in),
    .clk(_U1065_clk),
    .out(_U1065_out)
);
assign _U1066_in = _U1065_out;
assign _U1066_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1066 (
    .in(_U1066_in),
    .clk(_U1066_clk),
    .out(_U1066_out)
);
assign _U1067_in = _U1073_out;
_U1067_pt__U1068 _U1067 (
    .in(_U1067_in),
    .out(_U1067_out)
);
assign _U1069_in = 16'(_U1199_out * _U1049_out);
assign _U1069_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1069 (
    .in(_U1069_in),
    .clk(_U1069_clk),
    .out(_U1069_out)
);
assign _U1070_in = _U1069_out;
assign _U1070_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1070 (
    .in(_U1070_in),
    .clk(_U1070_clk),
    .out(_U1070_out)
);
assign _U1071_in = _U1070_out;
assign _U1071_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1071 (
    .in(_U1071_in),
    .clk(_U1071_clk),
    .out(_U1071_out)
);
assign _U1072_in = _U1071_out;
assign _U1072_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1072 (
    .in(_U1072_in),
    .clk(_U1072_clk),
    .out(_U1072_out)
);
assign _U1073_in = _U1072_out;
assign _U1073_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1073 (
    .in(_U1073_in),
    .clk(_U1073_clk),
    .out(_U1073_out)
);
assign _U1074_in = _U1089_out;
_U1074_pt__U1075 _U1074 (
    .in(_U1074_in),
    .out(_U1074_out)
);
assign _U1076_in = in0_conv_stencil[0];
assign _U1076_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1076 (
    .in(_U1076_in),
    .clk(_U1076_clk),
    .out(_U1076_out)
);
assign _U1077_in = _U1076_out;
assign _U1077_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1077 (
    .in(_U1077_in),
    .clk(_U1077_clk),
    .out(_U1077_out)
);
assign _U1078_in = _U1077_out;
assign _U1078_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1078 (
    .in(_U1078_in),
    .clk(_U1078_clk),
    .out(_U1078_out)
);
assign _U1079_in = _U1078_out;
assign _U1079_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1079 (
    .in(_U1079_in),
    .clk(_U1079_clk),
    .out(_U1079_out)
);
assign _U1080_in = _U1079_out;
assign _U1080_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1080 (
    .in(_U1080_in),
    .clk(_U1080_clk),
    .out(_U1080_out)
);
assign _U1081_in = _U1080_out;
assign _U1081_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1081 (
    .in(_U1081_in),
    .clk(_U1081_clk),
    .out(_U1081_out)
);
assign _U1082_in = _U1081_out;
assign _U1082_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1082 (
    .in(_U1082_in),
    .clk(_U1082_clk),
    .out(_U1082_out)
);
assign _U1083_in = _U1082_out;
assign _U1083_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1083 (
    .in(_U1083_in),
    .clk(_U1083_clk),
    .out(_U1083_out)
);
assign _U1084_in = _U1083_out;
assign _U1084_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1084 (
    .in(_U1084_in),
    .clk(_U1084_clk),
    .out(_U1084_out)
);
assign _U1085_in = _U1084_out;
assign _U1085_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1085 (
    .in(_U1085_in),
    .clk(_U1085_clk),
    .out(_U1085_out)
);
assign _U1086_in = _U1085_out;
assign _U1086_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1086 (
    .in(_U1086_in),
    .clk(_U1086_clk),
    .out(_U1086_out)
);
assign _U1087_in = _U1086_out;
assign _U1087_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1087 (
    .in(_U1087_in),
    .clk(_U1087_clk),
    .out(_U1087_out)
);
assign _U1088_in = _U1087_out;
assign _U1088_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1088 (
    .in(_U1088_in),
    .clk(_U1088_clk),
    .out(_U1088_out)
);
assign _U1089_in = _U1088_out;
assign _U1089_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1089 (
    .in(_U1089_in),
    .clk(_U1089_clk),
    .out(_U1089_out)
);
assign _U1090_in = _U1095_out;
_U1090_pt__U1091 _U1090 (
    .in(_U1090_in),
    .out(_U1090_out)
);
assign _U1092_in = in2_hw_kernel_global_wrapper_stencil[0];
assign _U1092_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1092 (
    .in(_U1092_in),
    .clk(_U1092_clk),
    .out(_U1092_out)
);
assign _U1093_in = _U1092_out;
assign _U1093_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1093 (
    .in(_U1093_in),
    .clk(_U1093_clk),
    .out(_U1093_out)
);
assign _U1094_in = _U1093_out;
assign _U1094_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1094 (
    .in(_U1094_in),
    .clk(_U1094_clk),
    .out(_U1094_out)
);
assign _U1095_in = _U1094_out;
assign _U1095_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1095 (
    .in(_U1095_in),
    .clk(_U1095_clk),
    .out(_U1095_out)
);
assign _U1096_in = _U1101_out;
_U1096_pt__U1097 _U1096 (
    .in(_U1096_in),
    .out(_U1096_out)
);
assign _U1098_in = in1_hw_input_global_wrapper_stencil[0];
assign _U1098_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1098 (
    .in(_U1098_in),
    .clk(_U1098_clk),
    .out(_U1098_out)
);
assign _U1099_in = _U1098_out;
assign _U1099_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1099 (
    .in(_U1099_in),
    .clk(_U1099_clk),
    .out(_U1099_out)
);
assign _U1100_in = _U1099_out;
assign _U1100_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1100 (
    .in(_U1100_in),
    .clk(_U1100_clk),
    .out(_U1100_out)
);
assign _U1101_in = _U1100_out;
assign _U1101_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1101 (
    .in(_U1101_in),
    .clk(_U1101_clk),
    .out(_U1101_out)
);
assign _U1102_in = _U1108_out;
_U1102_pt__U1103 _U1102 (
    .in(_U1102_in),
    .out(_U1102_out)
);
assign _U1104_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U1104_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1104 (
    .in(_U1104_in),
    .clk(_U1104_clk),
    .out(_U1104_out)
);
assign _U1105_in = _U1104_out;
assign _U1105_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1105 (
    .in(_U1105_in),
    .clk(_U1105_clk),
    .out(_U1105_out)
);
assign _U1106_in = _U1105_out;
assign _U1106_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1106 (
    .in(_U1106_in),
    .clk(_U1106_clk),
    .out(_U1106_out)
);
assign _U1107_in = _U1106_out;
assign _U1107_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1107 (
    .in(_U1107_in),
    .clk(_U1107_clk),
    .out(_U1107_out)
);
assign _U1108_in = _U1107_out;
assign _U1108_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1108 (
    .in(_U1108_in),
    .clk(_U1108_clk),
    .out(_U1108_out)
);
assign _U1109_in = _U1111_out;
_U1109_pt__U1110 _U1109 (
    .in(_U1109_in),
    .out(_U1109_out)
);
assign _U1111_in = 16'(_U1115_out + _U1123_out);
assign _U1111_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1111 (
    .in(_U1111_in),
    .clk(_U1111_clk),
    .out(_U1111_out)
);
assign _U1112_in = _U1114_out;
_U1112_pt__U1113 _U1112 (
    .in(_U1112_in),
    .out(_U1112_out)
);
assign _U1114_in = 16'(_U1039_out + _U1109_out);
assign _U1114_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1114 (
    .in(_U1114_in),
    .clk(_U1114_clk),
    .out(_U1114_out)
);
assign _U1115_in = _U1122_out;
_U1115_pt__U1116 _U1115 (
    .in(_U1115_in),
    .out(_U1115_out)
);
assign _U1117_in = 16'(_U1147_out * _U1155_out);
assign _U1117_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1117 (
    .in(_U1117_in),
    .clk(_U1117_clk),
    .out(_U1117_out)
);
assign _U1118_in = _U1117_out;
assign _U1118_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1118 (
    .in(_U1118_in),
    .clk(_U1118_clk),
    .out(_U1118_out)
);
assign _U1119_in = _U1118_out;
assign _U1119_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1119 (
    .in(_U1119_in),
    .clk(_U1119_clk),
    .out(_U1119_out)
);
assign _U1120_in = _U1119_out;
assign _U1120_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1120 (
    .in(_U1120_in),
    .clk(_U1120_clk),
    .out(_U1120_out)
);
assign _U1121_in = _U1120_out;
assign _U1121_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1121 (
    .in(_U1121_in),
    .clk(_U1121_clk),
    .out(_U1121_out)
);
assign _U1122_in = _U1121_out;
assign _U1122_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1122 (
    .in(_U1122_in),
    .clk(_U1122_clk),
    .out(_U1122_out)
);
assign _U1123_in = _U1125_out;
_U1123_pt__U1124 _U1123 (
    .in(_U1123_in),
    .out(_U1123_out)
);
assign _U1125_in = 16'(_U1126_out + _U1132_out);
assign _U1125_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1125 (
    .in(_U1125_in),
    .clk(_U1125_clk),
    .out(_U1125_out)
);
assign _U1126_in = _U1131_out;
_U1126_pt__U1127 _U1126 (
    .in(_U1126_in),
    .out(_U1126_out)
);
assign _U1128_in = 16'(_U1163_out * _U1172_out);
assign _U1128_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1128 (
    .in(_U1128_in),
    .clk(_U1128_clk),
    .out(_U1128_out)
);
assign _U1129_in = _U1128_out;
assign _U1129_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1129 (
    .in(_U1129_in),
    .clk(_U1129_clk),
    .out(_U1129_out)
);
assign _U1130_in = _U1129_out;
assign _U1130_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1130 (
    .in(_U1130_in),
    .clk(_U1130_clk),
    .out(_U1130_out)
);
assign _U1131_in = _U1130_out;
assign _U1131_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1131 (
    .in(_U1131_in),
    .clk(_U1131_clk),
    .out(_U1131_out)
);
assign _U1132_in = _U1134_out;
_U1132_pt__U1133 _U1132 (
    .in(_U1132_in),
    .out(_U1132_out)
);
assign _U1134_in = 16'(_U1204_out + _U1216_out);
assign _U1134_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1134 (
    .in(_U1134_in),
    .clk(_U1134_clk),
    .out(_U1134_out)
);
assign _U1135_in = _U1137_out;
_U1135_pt__U1136 _U1135 (
    .in(_U1135_in),
    .out(_U1135_out)
);
assign _U1137_in = 16'(_U1074_out + _U1112_out);
assign _U1137_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1137 (
    .in(_U1137_in),
    .clk(_U1137_clk),
    .out(_U1137_out)
);
assign _U1138_in = 16'(_U1054_out + _U1135_out);
_U1138_pt__U1139 _U1138 (
    .in(_U1138_in),
    .out(out_conv_stencil)
);
assign _U1140_in = _U1146_out;
_U1140_pt__U1141 _U1140 (
    .in(_U1140_in),
    .out(_U1140_out)
);
assign _U1142_in = in1_hw_input_global_wrapper_stencil[1];
assign _U1142_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1142 (
    .in(_U1142_in),
    .clk(_U1142_clk),
    .out(_U1142_out)
);
assign _U1143_in = _U1142_out;
assign _U1143_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1143 (
    .in(_U1143_in),
    .clk(_U1143_clk),
    .out(_U1143_out)
);
assign _U1144_in = _U1143_out;
assign _U1144_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1144 (
    .in(_U1144_in),
    .clk(_U1144_clk),
    .out(_U1144_out)
);
assign _U1145_in = _U1144_out;
assign _U1145_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1145 (
    .in(_U1145_in),
    .clk(_U1145_clk),
    .out(_U1145_out)
);
assign _U1146_in = _U1145_out;
assign _U1146_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1146 (
    .in(_U1146_in),
    .clk(_U1146_clk),
    .out(_U1146_out)
);
assign _U1147_in = _U1154_out;
_U1147_pt__U1148 _U1147 (
    .in(_U1147_in),
    .out(_U1147_out)
);
assign _U1149_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U1149_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1149 (
    .in(_U1149_in),
    .clk(_U1149_clk),
    .out(_U1149_out)
);
assign _U1150_in = _U1149_out;
assign _U1150_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1150 (
    .in(_U1150_in),
    .clk(_U1150_clk),
    .out(_U1150_out)
);
assign _U1151_in = _U1150_out;
assign _U1151_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1151 (
    .in(_U1151_in),
    .clk(_U1151_clk),
    .out(_U1151_out)
);
assign _U1152_in = _U1151_out;
assign _U1152_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1152 (
    .in(_U1152_in),
    .clk(_U1152_clk),
    .out(_U1152_out)
);
assign _U1153_in = _U1152_out;
assign _U1153_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1153 (
    .in(_U1153_in),
    .clk(_U1153_clk),
    .out(_U1153_out)
);
assign _U1154_in = _U1153_out;
assign _U1154_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1154 (
    .in(_U1154_in),
    .clk(_U1154_clk),
    .out(_U1154_out)
);
assign _U1155_in = _U1162_out;
_U1155_pt__U1156 _U1155 (
    .in(_U1155_in),
    .out(_U1155_out)
);
assign _U1157_in = in1_hw_input_global_wrapper_stencil[2];
assign _U1157_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1157 (
    .in(_U1157_in),
    .clk(_U1157_clk),
    .out(_U1157_out)
);
assign _U1158_in = _U1157_out;
assign _U1158_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1158 (
    .in(_U1158_in),
    .clk(_U1158_clk),
    .out(_U1158_out)
);
assign _U1159_in = _U1158_out;
assign _U1159_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1159 (
    .in(_U1159_in),
    .clk(_U1159_clk),
    .out(_U1159_out)
);
assign _U1160_in = _U1159_out;
assign _U1160_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1160 (
    .in(_U1160_in),
    .clk(_U1160_clk),
    .out(_U1160_out)
);
assign _U1161_in = _U1160_out;
assign _U1161_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1161 (
    .in(_U1161_in),
    .clk(_U1161_clk),
    .out(_U1161_out)
);
assign _U1162_in = _U1161_out;
assign _U1162_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1162 (
    .in(_U1162_in),
    .clk(_U1162_clk),
    .out(_U1162_out)
);
assign _U1163_in = _U1171_out;
_U1163_pt__U1164 _U1163 (
    .in(_U1163_in),
    .out(_U1163_out)
);
assign _U1165_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U1165_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1165 (
    .in(_U1165_in),
    .clk(_U1165_clk),
    .out(_U1165_out)
);
assign _U1166_in = _U1165_out;
assign _U1166_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1166 (
    .in(_U1166_in),
    .clk(_U1166_clk),
    .out(_U1166_out)
);
assign _U1167_in = _U1166_out;
assign _U1167_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1167 (
    .in(_U1167_in),
    .clk(_U1167_clk),
    .out(_U1167_out)
);
assign _U1168_in = _U1167_out;
assign _U1168_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1168 (
    .in(_U1168_in),
    .clk(_U1168_clk),
    .out(_U1168_out)
);
assign _U1169_in = _U1168_out;
assign _U1169_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1169 (
    .in(_U1169_in),
    .clk(_U1169_clk),
    .out(_U1169_out)
);
assign _U1170_in = _U1169_out;
assign _U1170_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1170 (
    .in(_U1170_in),
    .clk(_U1170_clk),
    .out(_U1170_out)
);
assign _U1171_in = _U1170_out;
assign _U1171_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1171 (
    .in(_U1171_in),
    .clk(_U1171_clk),
    .out(_U1171_out)
);
assign _U1172_in = _U1180_out;
_U1172_pt__U1173 _U1172 (
    .in(_U1172_in),
    .out(_U1172_out)
);
assign _U1174_in = in1_hw_input_global_wrapper_stencil[3];
assign _U1174_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1174 (
    .in(_U1174_in),
    .clk(_U1174_clk),
    .out(_U1174_out)
);
assign _U1175_in = _U1174_out;
assign _U1175_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1175 (
    .in(_U1175_in),
    .clk(_U1175_clk),
    .out(_U1175_out)
);
assign _U1176_in = _U1175_out;
assign _U1176_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1176 (
    .in(_U1176_in),
    .clk(_U1176_clk),
    .out(_U1176_out)
);
assign _U1177_in = _U1176_out;
assign _U1177_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1177 (
    .in(_U1177_in),
    .clk(_U1177_clk),
    .out(_U1177_out)
);
assign _U1178_in = _U1177_out;
assign _U1178_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1178 (
    .in(_U1178_in),
    .clk(_U1178_clk),
    .out(_U1178_out)
);
assign _U1179_in = _U1178_out;
assign _U1179_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1179 (
    .in(_U1179_in),
    .clk(_U1179_clk),
    .out(_U1179_out)
);
assign _U1180_in = _U1179_out;
assign _U1180_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1180 (
    .in(_U1180_in),
    .clk(_U1180_clk),
    .out(_U1180_out)
);
assign _U1181_in = in2_hw_kernel_global_wrapper_stencil[4];
_U1181_pt__U1182 _U1181 (
    .in(_U1181_in),
    .out(_U1181_out)
);
assign _U1183_in = in1_hw_input_global_wrapper_stencil[4];
_U1183_pt__U1184 _U1183 (
    .in(_U1183_in),
    .out(_U1183_out)
);
assign _U1185_in = _U1187_out;
_U1185_pt__U1186 _U1185 (
    .in(_U1185_in),
    .out(_U1185_out)
);
assign _U1187_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U1187_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1187 (
    .in(_U1187_in),
    .clk(_U1187_clk),
    .out(_U1187_out)
);
assign _U1188_in = _U1190_out;
_U1188_pt__U1189 _U1188 (
    .in(_U1188_in),
    .out(_U1188_out)
);
assign _U1190_in = in1_hw_input_global_wrapper_stencil[5];
assign _U1190_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1190 (
    .in(_U1190_in),
    .clk(_U1190_clk),
    .out(_U1190_out)
);
assign _U1191_in = _U1194_out;
_U1191_pt__U1192 _U1191 (
    .in(_U1191_in),
    .out(_U1191_out)
);
assign _U1193_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U1193_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1193 (
    .in(_U1193_in),
    .clk(_U1193_clk),
    .out(_U1193_out)
);
assign _U1194_in = _U1193_out;
assign _U1194_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1194 (
    .in(_U1194_in),
    .clk(_U1194_clk),
    .out(_U1194_out)
);
assign _U1195_in = _U1198_out;
_U1195_pt__U1196 _U1195 (
    .in(_U1195_in),
    .out(_U1195_out)
);
assign _U1197_in = in1_hw_input_global_wrapper_stencil[6];
assign _U1197_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1197 (
    .in(_U1197_in),
    .clk(_U1197_clk),
    .out(_U1197_out)
);
assign _U1198_in = _U1197_out;
assign _U1198_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1198 (
    .in(_U1198_in),
    .clk(_U1198_clk),
    .out(_U1198_out)
);
assign _U1199_in = _U1203_out;
_U1199_pt__U1200 _U1199 (
    .in(_U1199_in),
    .out(_U1199_out)
);
assign _U1201_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U1201_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1201 (
    .in(_U1201_in),
    .clk(_U1201_clk),
    .out(_U1201_out)
);
assign _U1202_in = _U1201_out;
assign _U1202_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1202 (
    .in(_U1202_in),
    .clk(_U1202_clk),
    .out(_U1202_out)
);
assign _U1203_in = _U1202_out;
assign _U1203_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1203 (
    .in(_U1203_in),
    .clk(_U1203_clk),
    .out(_U1203_out)
);
assign _U1204_in = _U1215_out;
_U1204_pt__U1205 _U1204 (
    .in(_U1204_in),
    .out(_U1204_out)
);
assign _U1206_in = 16'(_U1181_out * _U1183_out);
assign _U1206_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1206 (
    .in(_U1206_in),
    .clk(_U1206_clk),
    .out(_U1206_out)
);
assign _U1207_in = _U1206_out;
assign _U1207_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1207 (
    .in(_U1207_in),
    .clk(_U1207_clk),
    .out(_U1207_out)
);
assign _U1208_in = _U1207_out;
assign _U1208_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1208 (
    .in(_U1208_in),
    .clk(_U1208_clk),
    .out(_U1208_out)
);
assign _U1209_in = _U1208_out;
assign _U1209_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1209 (
    .in(_U1209_in),
    .clk(_U1209_clk),
    .out(_U1209_out)
);
assign _U1210_in = _U1209_out;
assign _U1210_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1210 (
    .in(_U1210_in),
    .clk(_U1210_clk),
    .out(_U1210_out)
);
assign _U1211_in = _U1210_out;
assign _U1211_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1211 (
    .in(_U1211_in),
    .clk(_U1211_clk),
    .out(_U1211_out)
);
assign _U1212_in = _U1211_out;
assign _U1212_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1212 (
    .in(_U1212_in),
    .clk(_U1212_clk),
    .out(_U1212_out)
);
assign _U1213_in = _U1212_out;
assign _U1213_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1213 (
    .in(_U1213_in),
    .clk(_U1213_clk),
    .out(_U1213_out)
);
assign _U1214_in = _U1213_out;
assign _U1214_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1214 (
    .in(_U1214_in),
    .clk(_U1214_clk),
    .out(_U1214_out)
);
assign _U1215_in = _U1214_out;
assign _U1215_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1215 (
    .in(_U1215_in),
    .clk(_U1215_clk),
    .out(_U1215_out)
);
assign _U1216_in = _U1218_out;
_U1216_pt__U1217 _U1216 (
    .in(_U1216_in),
    .out(_U1216_out)
);
assign _U1218_in = 16'(_U1219_out + _U1229_out);
assign _U1218_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1218 (
    .in(_U1218_in),
    .clk(_U1218_clk),
    .out(_U1218_out)
);
assign _U1219_in = _U1228_out;
_U1219_pt__U1220 _U1219 (
    .in(_U1219_in),
    .out(_U1219_out)
);
assign _U1221_in = 16'(_U1185_out * _U1188_out);
assign _U1221_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1221 (
    .in(_U1221_in),
    .clk(_U1221_clk),
    .out(_U1221_out)
);
assign _U1222_in = _U1221_out;
assign _U1222_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1222 (
    .in(_U1222_in),
    .clk(_U1222_clk),
    .out(_U1222_out)
);
assign _U1223_in = _U1222_out;
assign _U1223_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1223 (
    .in(_U1223_in),
    .clk(_U1223_clk),
    .out(_U1223_out)
);
assign _U1224_in = _U1223_out;
assign _U1224_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1224 (
    .in(_U1224_in),
    .clk(_U1224_clk),
    .out(_U1224_out)
);
assign _U1225_in = _U1224_out;
assign _U1225_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1225 (
    .in(_U1225_in),
    .clk(_U1225_clk),
    .out(_U1225_out)
);
assign _U1226_in = _U1225_out;
assign _U1226_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1226 (
    .in(_U1226_in),
    .clk(_U1226_clk),
    .out(_U1226_out)
);
assign _U1227_in = _U1226_out;
assign _U1227_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1227 (
    .in(_U1227_in),
    .clk(_U1227_clk),
    .out(_U1227_out)
);
assign _U1228_in = _U1227_out;
assign _U1228_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1228 (
    .in(_U1228_in),
    .clk(_U1228_clk),
    .out(_U1228_out)
);
assign _U1229_in = _U1231_out;
_U1229_pt__U1230 _U1229 (
    .in(_U1229_in),
    .out(_U1229_out)
);
assign _U1231_in = 16'(_U1232_out + _U1067_out);
assign _U1231_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1231 (
    .in(_U1231_in),
    .clk(_U1231_clk),
    .out(_U1231_out)
);
assign _U1232_in = _U1239_out;
_U1232_pt__U1233 _U1232 (
    .in(_U1232_in),
    .out(_U1232_out)
);
assign _U1234_in = 16'(_U1191_out * _U1195_out);
assign _U1234_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1234 (
    .in(_U1234_in),
    .clk(_U1234_clk),
    .out(_U1234_out)
);
assign _U1235_in = _U1234_out;
assign _U1235_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1235 (
    .in(_U1235_in),
    .clk(_U1235_clk),
    .out(_U1235_out)
);
assign _U1236_in = _U1235_out;
assign _U1236_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1236 (
    .in(_U1236_in),
    .clk(_U1236_clk),
    .out(_U1236_out)
);
assign _U1237_in = _U1236_out;
assign _U1237_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1237 (
    .in(_U1237_in),
    .clk(_U1237_clk),
    .out(_U1237_out)
);
assign _U1238_in = _U1237_out;
assign _U1238_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1238 (
    .in(_U1238_in),
    .clk(_U1238_clk),
    .out(_U1238_out)
);
assign _U1239_in = _U1238_out;
assign _U1239_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1239 (
    .in(_U1239_in),
    .clk(_U1239_clk),
    .out(_U1239_out)
);
endmodule

module cu_op_hcompute_conv_stencil_13 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_13_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_13_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_13_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[0];
hcompute_conv_stencil_13_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_13_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U1030_pt__U1031 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1026_pt__U1027 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1018_pt__U1019 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1010_pt__U1011 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1007_pt__U1008 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1004_pt__U1005 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U1002_pt__U1003 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_12_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U1000_in;
wire _U1000_clk;
wire [15:0] _U1000_out;
wire [15:0] _U1001_in;
wire _U1001_clk;
wire [15:0] _U1001_out;
wire [15:0] _U1002_in;
wire [15:0] _U1004_in;
wire [15:0] _U1004_out;
wire [15:0] _U1006_in;
wire _U1006_clk;
wire [15:0] _U1006_out;
wire [15:0] _U1007_in;
wire [15:0] _U1007_out;
wire [15:0] _U1009_in;
wire _U1009_clk;
wire [15:0] _U1009_out;
wire [15:0] _U1010_in;
wire [15:0] _U1010_out;
wire [15:0] _U1012_in;
wire _U1012_clk;
wire [15:0] _U1012_out;
wire [15:0] _U1013_in;
wire _U1013_clk;
wire [15:0] _U1013_out;
wire [15:0] _U1014_in;
wire _U1014_clk;
wire [15:0] _U1014_out;
wire [15:0] _U1015_in;
wire _U1015_clk;
wire [15:0] _U1015_out;
wire [15:0] _U1016_in;
wire _U1016_clk;
wire [15:0] _U1016_out;
wire [15:0] _U1017_in;
wire _U1017_clk;
wire [15:0] _U1017_out;
wire [15:0] _U1018_in;
wire [15:0] _U1018_out;
wire [15:0] _U1020_in;
wire _U1020_clk;
wire [15:0] _U1020_out;
wire [15:0] _U1021_in;
wire _U1021_clk;
wire [15:0] _U1021_out;
wire [15:0] _U1022_in;
wire _U1022_clk;
wire [15:0] _U1022_out;
wire [15:0] _U1023_in;
wire _U1023_clk;
wire [15:0] _U1023_out;
wire [15:0] _U1024_in;
wire _U1024_clk;
wire [15:0] _U1024_out;
wire [15:0] _U1025_in;
wire _U1025_clk;
wire [15:0] _U1025_out;
wire [15:0] _U1026_in;
wire [15:0] _U1026_out;
wire [15:0] _U1028_in;
wire _U1028_clk;
wire [15:0] _U1028_out;
wire [15:0] _U1029_in;
wire _U1029_clk;
wire [15:0] _U1029_out;
wire [15:0] _U1030_in;
wire [15:0] _U1030_out;
wire [15:0] _U1032_in;
wire _U1032_clk;
wire [15:0] _U1032_out;
wire [15:0] _U1033_in;
wire _U1033_clk;
wire [15:0] _U1033_out;
wire [15:0] _U1034_in;
wire _U1034_clk;
wire [15:0] _U1034_out;
wire [15:0] _U1035_in;
wire _U1035_clk;
wire [15:0] _U1035_out;
wire [15:0] _U1036_in;
wire _U1036_clk;
wire [15:0] _U1036_out;
wire [15:0] _U1037_in;
wire _U1037_clk;
wire [15:0] _U1037_out;
wire [15:0] _U1038_in;
wire _U1038_clk;
wire [15:0] _U1038_out;
wire [15:0] _U838_in;
wire [15:0] _U838_out;
wire [15:0] _U840_in;
wire _U840_clk;
wire [15:0] _U840_out;
wire [15:0] _U841_in;
wire _U841_clk;
wire [15:0] _U841_out;
wire [15:0] _U842_in;
wire _U842_clk;
wire [15:0] _U842_out;
wire [15:0] _U843_in;
wire _U843_clk;
wire [15:0] _U843_out;
wire [15:0] _U844_in;
wire _U844_clk;
wire [15:0] _U844_out;
wire [15:0] _U845_in;
wire _U845_clk;
wire [15:0] _U845_out;
wire [15:0] _U846_in;
wire _U846_clk;
wire [15:0] _U846_out;
wire [15:0] _U847_in;
wire _U847_clk;
wire [15:0] _U847_out;
wire [15:0] _U848_in;
wire _U848_clk;
wire [15:0] _U848_out;
wire [15:0] _U849_in;
wire _U849_clk;
wire [15:0] _U849_out;
wire [15:0] _U850_in;
wire _U850_clk;
wire [15:0] _U850_out;
wire [15:0] _U851_in;
wire _U851_clk;
wire [15:0] _U851_out;
wire [15:0] _U852_in;
wire _U852_clk;
wire [15:0] _U852_out;
wire [15:0] _U853_in;
wire _U853_clk;
wire [15:0] _U853_out;
wire [15:0] _U854_in;
wire [15:0] _U854_out;
wire [15:0] _U856_in;
wire _U856_clk;
wire [15:0] _U856_out;
wire [15:0] _U857_in;
wire _U857_clk;
wire [15:0] _U857_out;
wire [15:0] _U858_in;
wire _U858_clk;
wire [15:0] _U858_out;
wire [15:0] _U859_in;
wire _U859_clk;
wire [15:0] _U859_out;
wire [15:0] _U860_in;
wire _U860_clk;
wire [15:0] _U860_out;
wire [15:0] _U861_in;
wire _U861_clk;
wire [15:0] _U861_out;
wire [15:0] _U862_in;
wire _U862_clk;
wire [15:0] _U862_out;
wire [15:0] _U863_in;
wire _U863_clk;
wire [15:0] _U863_out;
wire [15:0] _U864_in;
wire _U864_clk;
wire [15:0] _U864_out;
wire [15:0] _U865_in;
wire _U865_clk;
wire [15:0] _U865_out;
wire [15:0] _U866_in;
wire _U866_clk;
wire [15:0] _U866_out;
wire [15:0] _U867_in;
wire _U867_clk;
wire [15:0] _U867_out;
wire [15:0] _U868_in;
wire _U868_clk;
wire [15:0] _U868_out;
wire [15:0] _U869_in;
wire _U869_clk;
wire [15:0] _U869_out;
wire [15:0] _U870_in;
wire [15:0] _U870_out;
wire [15:0] _U872_in;
wire _U872_clk;
wire [15:0] _U872_out;
wire [15:0] _U873_in;
wire [15:0] _U873_out;
wire [15:0] _U875_in;
wire _U875_clk;
wire [15:0] _U875_out;
wire [15:0] _U876_in;
wire _U876_clk;
wire [15:0] _U876_out;
wire [15:0] _U877_in;
wire _U877_clk;
wire [15:0] _U877_out;
wire [15:0] _U878_in;
wire _U878_clk;
wire [15:0] _U878_out;
wire [15:0] _U879_in;
wire _U879_clk;
wire [15:0] _U879_out;
wire [15:0] _U880_in;
wire _U880_clk;
wire [15:0] _U880_out;
wire [15:0] _U881_in;
wire [15:0] _U881_out;
wire [15:0] _U883_in;
wire _U883_clk;
wire [15:0] _U883_out;
wire [15:0] _U884_in;
wire _U884_clk;
wire [15:0] _U884_out;
wire [15:0] _U885_in;
wire _U885_clk;
wire [15:0] _U885_out;
wire [15:0] _U886_in;
wire _U886_clk;
wire [15:0] _U886_out;
wire [15:0] _U887_in;
wire _U887_clk;
wire [15:0] _U887_out;
wire [15:0] _U888_in;
wire [15:0] _U888_out;
wire [15:0] _U890_in;
wire _U890_clk;
wire [15:0] _U890_out;
wire [15:0] _U891_in;
wire _U891_clk;
wire [15:0] _U891_out;
wire [15:0] _U892_in;
wire _U892_clk;
wire [15:0] _U892_out;
wire [15:0] _U893_in;
wire _U893_clk;
wire [15:0] _U893_out;
wire [15:0] _U894_in;
wire _U894_clk;
wire [15:0] _U894_out;
wire [15:0] _U895_in;
wire _U895_clk;
wire [15:0] _U895_out;
wire [15:0] _U896_in;
wire _U896_clk;
wire [15:0] _U896_out;
wire [15:0] _U897_in;
wire _U897_clk;
wire [15:0] _U897_out;
wire [15:0] _U898_in;
wire [15:0] _U898_out;
wire [15:0] _U900_in;
wire _U900_clk;
wire [15:0] _U900_out;
wire [15:0] _U901_in;
wire [15:0] _U901_out;
wire [15:0] _U903_in;
wire _U903_clk;
wire [15:0] _U903_out;
wire [15:0] _U904_in;
wire [15:0] _U904_out;
wire [15:0] _U906_in;
wire _U906_clk;
wire [15:0] _U906_out;
wire [15:0] _U907_in;
wire _U907_clk;
wire [15:0] _U907_out;
wire [15:0] _U908_in;
wire [15:0] _U908_out;
wire [15:0] _U910_in;
wire [15:0] _U910_out;
wire [15:0] _U912_in;
wire [15:0] _U912_out;
wire [15:0] _U914_in;
wire _U914_clk;
wire [15:0] _U914_out;
wire [15:0] _U915_in;
wire _U915_clk;
wire [15:0] _U915_out;
wire [15:0] _U916_in;
wire _U916_clk;
wire [15:0] _U916_out;
wire [15:0] _U917_in;
wire _U917_clk;
wire [15:0] _U917_out;
wire [15:0] _U918_in;
wire [15:0] _U918_out;
wire [15:0] _U920_in;
wire _U920_clk;
wire [15:0] _U920_out;
wire [15:0] _U921_in;
wire _U921_clk;
wire [15:0] _U921_out;
wire [15:0] _U922_in;
wire _U922_clk;
wire [15:0] _U922_out;
wire [15:0] _U923_in;
wire _U923_clk;
wire [15:0] _U923_out;
wire [15:0] _U924_in;
wire [15:0] _U924_out;
wire [15:0] _U926_in;
wire _U926_clk;
wire [15:0] _U926_out;
wire [15:0] _U927_in;
wire [15:0] _U927_out;
wire [15:0] _U929_in;
wire _U929_clk;
wire [15:0] _U929_out;
wire [15:0] _U930_in;
wire _U930_clk;
wire [15:0] _U930_out;
wire [15:0] _U931_in;
wire _U931_clk;
wire [15:0] _U931_out;
wire [15:0] _U932_in;
wire _U932_clk;
wire [15:0] _U932_out;
wire [15:0] _U933_in;
wire _U933_clk;
wire [15:0] _U933_out;
wire [15:0] _U934_in;
wire [15:0] _U934_out;
wire [15:0] _U936_in;
wire _U936_clk;
wire [15:0] _U936_out;
wire [15:0] _U937_in;
wire _U937_clk;
wire [15:0] _U937_out;
wire [15:0] _U938_in;
wire _U938_clk;
wire [15:0] _U938_out;
wire [15:0] _U939_in;
wire _U939_clk;
wire [15:0] _U939_out;
wire [15:0] _U940_in;
wire _U940_clk;
wire [15:0] _U940_out;
wire [15:0] _U941_in;
wire [15:0] _U941_out;
wire [15:0] _U943_in;
wire _U943_clk;
wire [15:0] _U943_out;
wire [15:0] _U944_in;
wire _U944_clk;
wire [15:0] _U944_out;
wire [15:0] _U945_in;
wire _U945_clk;
wire [15:0] _U945_out;
wire [15:0] _U946_in;
wire [15:0] _U946_out;
wire [15:0] _U948_in;
wire _U948_clk;
wire [15:0] _U948_out;
wire [15:0] _U949_in;
wire _U949_clk;
wire [15:0] _U949_out;
wire [15:0] _U950_in;
wire _U950_clk;
wire [15:0] _U950_out;
wire [15:0] _U951_in;
wire [15:0] _U951_out;
wire [15:0] _U953_in;
wire _U953_clk;
wire [15:0] _U953_out;
wire [15:0] _U954_in;
wire _U954_clk;
wire [15:0] _U954_out;
wire [15:0] _U955_in;
wire _U955_clk;
wire [15:0] _U955_out;
wire [15:0] _U956_in;
wire _U956_clk;
wire [15:0] _U956_out;
wire [15:0] _U957_in;
wire _U957_clk;
wire [15:0] _U957_out;
wire [15:0] _U958_in;
wire _U958_clk;
wire [15:0] _U958_out;
wire [15:0] _U959_in;
wire _U959_clk;
wire [15:0] _U959_out;
wire [15:0] _U960_in;
wire _U960_clk;
wire [15:0] _U960_out;
wire [15:0] _U961_in;
wire _U961_clk;
wire [15:0] _U961_out;
wire [15:0] _U962_in;
wire _U962_clk;
wire [15:0] _U962_out;
wire [15:0] _U963_in;
wire [15:0] _U963_out;
wire [15:0] _U965_in;
wire _U965_clk;
wire [15:0] _U965_out;
wire [15:0] _U966_in;
wire [15:0] _U966_out;
wire [15:0] _U968_in;
wire _U968_clk;
wire [15:0] _U968_out;
wire [15:0] _U969_in;
wire [15:0] _U969_out;
wire [15:0] _U971_in;
wire _U971_clk;
wire [15:0] _U971_out;
wire [15:0] _U972_in;
wire _U972_clk;
wire [15:0] _U972_out;
wire [15:0] _U973_in;
wire _U973_clk;
wire [15:0] _U973_out;
wire [15:0] _U974_in;
wire _U974_clk;
wire [15:0] _U974_out;
wire [15:0] _U975_in;
wire _U975_clk;
wire [15:0] _U975_out;
wire [15:0] _U976_in;
wire _U976_clk;
wire [15:0] _U976_out;
wire [15:0] _U977_in;
wire _U977_clk;
wire [15:0] _U977_out;
wire [15:0] _U978_in;
wire [15:0] _U978_out;
wire [15:0] _U980_in;
wire _U980_clk;
wire [15:0] _U980_out;
wire [15:0] _U981_in;
wire [15:0] _U981_out;
wire [15:0] _U983_in;
wire _U983_clk;
wire [15:0] _U983_out;
wire [15:0] _U984_in;
wire _U984_clk;
wire [15:0] _U984_out;
wire [15:0] _U985_in;
wire _U985_clk;
wire [15:0] _U985_out;
wire [15:0] _U986_in;
wire _U986_clk;
wire [15:0] _U986_out;
wire [15:0] _U987_in;
wire _U987_clk;
wire [15:0] _U987_out;
wire [15:0] _U988_in;
wire _U988_clk;
wire [15:0] _U988_out;
wire [15:0] _U989_in;
wire _U989_clk;
wire [15:0] _U989_out;
wire [15:0] _U990_in;
wire [15:0] _U990_out;
wire [15:0] _U992_in;
wire _U992_clk;
wire [15:0] _U992_out;
wire [15:0] _U993_in;
wire _U993_clk;
wire [15:0] _U993_out;
wire [15:0] _U994_in;
wire _U994_clk;
wire [15:0] _U994_out;
wire [15:0] _U995_in;
wire _U995_clk;
wire [15:0] _U995_out;
wire [15:0] _U996_in;
wire [15:0] _U996_out;
wire [15:0] _U998_in;
wire _U998_clk;
wire [15:0] _U998_out;
wire [15:0] _U999_in;
wire _U999_clk;
wire [15:0] _U999_out;
assign _U1000_in = _U999_out;
assign _U1000_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1000 (
    .in(_U1000_in),
    .clk(_U1000_clk),
    .out(_U1000_out)
);
assign _U1001_in = _U1000_out;
assign _U1001_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1001 (
    .in(_U1001_in),
    .clk(_U1001_clk),
    .out(_U1001_out)
);
assign _U1002_in = 16'(_U854_out + _U1004_out);
_U1002_pt__U1003 _U1002 (
    .in(_U1002_in),
    .out(out_conv_stencil)
);
assign _U1004_in = _U1006_out;
_U1004_pt__U1005 _U1004 (
    .in(_U1004_in),
    .out(_U1004_out)
);
assign _U1006_in = 16'(_U838_out + _U1007_out);
assign _U1006_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1006 (
    .in(_U1006_in),
    .clk(_U1006_clk),
    .out(_U1006_out)
);
assign _U1007_in = _U1009_out;
_U1007_pt__U1008 _U1007 (
    .in(_U1007_in),
    .out(_U1007_out)
);
assign _U1009_in = 16'(_U969_out + _U978_out);
assign _U1009_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1009 (
    .in(_U1009_in),
    .clk(_U1009_clk),
    .out(_U1009_out)
);
assign _U1010_in = _U1017_out;
_U1010_pt__U1011 _U1010 (
    .in(_U1010_in),
    .out(_U1010_out)
);
assign _U1012_in = 16'(_U990_out * _U918_out);
assign _U1012_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1012 (
    .in(_U1012_in),
    .clk(_U1012_clk),
    .out(_U1012_out)
);
assign _U1013_in = _U1012_out;
assign _U1013_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1013 (
    .in(_U1013_in),
    .clk(_U1013_clk),
    .out(_U1013_out)
);
assign _U1014_in = _U1013_out;
assign _U1014_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1014 (
    .in(_U1014_in),
    .clk(_U1014_clk),
    .out(_U1014_out)
);
assign _U1015_in = _U1014_out;
assign _U1015_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1015 (
    .in(_U1015_in),
    .clk(_U1015_clk),
    .out(_U1015_out)
);
assign _U1016_in = _U1015_out;
assign _U1016_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1016 (
    .in(_U1016_in),
    .clk(_U1016_clk),
    .out(_U1016_out)
);
assign _U1017_in = _U1016_out;
assign _U1017_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1017 (
    .in(_U1017_in),
    .clk(_U1017_clk),
    .out(_U1017_out)
);
assign _U1018_in = _U1025_out;
_U1018_pt__U1019 _U1018 (
    .in(_U1018_in),
    .out(_U1018_out)
);
assign _U1020_in = in1_hw_input_global_wrapper_stencil[1];
assign _U1020_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1020 (
    .in(_U1020_in),
    .clk(_U1020_clk),
    .out(_U1020_out)
);
assign _U1021_in = _U1020_out;
assign _U1021_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1021 (
    .in(_U1021_in),
    .clk(_U1021_clk),
    .out(_U1021_out)
);
assign _U1022_in = _U1021_out;
assign _U1022_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1022 (
    .in(_U1022_in),
    .clk(_U1022_clk),
    .out(_U1022_out)
);
assign _U1023_in = _U1022_out;
assign _U1023_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1023 (
    .in(_U1023_in),
    .clk(_U1023_clk),
    .out(_U1023_out)
);
assign _U1024_in = _U1023_out;
assign _U1024_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1024 (
    .in(_U1024_in),
    .clk(_U1024_clk),
    .out(_U1024_out)
);
assign _U1025_in = _U1024_out;
assign _U1025_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1025 (
    .in(_U1025_in),
    .clk(_U1025_clk),
    .out(_U1025_out)
);
assign _U1026_in = _U1029_out;
_U1026_pt__U1027 _U1026 (
    .in(_U1026_in),
    .out(_U1026_out)
);
assign _U1028_in = in1_hw_input_global_wrapper_stencil[2];
assign _U1028_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1028 (
    .in(_U1028_in),
    .clk(_U1028_clk),
    .out(_U1028_out)
);
assign _U1029_in = _U1028_out;
assign _U1029_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1029 (
    .in(_U1029_in),
    .clk(_U1029_clk),
    .out(_U1029_out)
);
assign _U1030_in = _U1038_out;
_U1030_pt__U1031 _U1030 (
    .in(_U1030_in),
    .out(_U1030_out)
);
assign _U1032_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U1032_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1032 (
    .in(_U1032_in),
    .clk(_U1032_clk),
    .out(_U1032_out)
);
assign _U1033_in = _U1032_out;
assign _U1033_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1033 (
    .in(_U1033_in),
    .clk(_U1033_clk),
    .out(_U1033_out)
);
assign _U1034_in = _U1033_out;
assign _U1034_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1034 (
    .in(_U1034_in),
    .clk(_U1034_clk),
    .out(_U1034_out)
);
assign _U1035_in = _U1034_out;
assign _U1035_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1035 (
    .in(_U1035_in),
    .clk(_U1035_clk),
    .out(_U1035_out)
);
assign _U1036_in = _U1035_out;
assign _U1036_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1036 (
    .in(_U1036_in),
    .clk(_U1036_clk),
    .out(_U1036_out)
);
assign _U1037_in = _U1036_out;
assign _U1037_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1037 (
    .in(_U1037_in),
    .clk(_U1037_clk),
    .out(_U1037_out)
);
assign _U1038_in = _U1037_out;
assign _U1038_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U1038 (
    .in(_U1038_in),
    .clk(_U1038_clk),
    .out(_U1038_out)
);
assign _U838_in = _U853_out;
_U838_pt__U839 _U838 (
    .in(_U838_in),
    .out(_U838_out)
);
assign _U840_in = in0_conv_stencil[0];
assign _U840_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U840 (
    .in(_U840_in),
    .clk(_U840_clk),
    .out(_U840_out)
);
assign _U841_in = _U840_out;
assign _U841_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U841 (
    .in(_U841_in),
    .clk(_U841_clk),
    .out(_U841_out)
);
assign _U842_in = _U841_out;
assign _U842_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U842 (
    .in(_U842_in),
    .clk(_U842_clk),
    .out(_U842_out)
);
assign _U843_in = _U842_out;
assign _U843_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U843 (
    .in(_U843_in),
    .clk(_U843_clk),
    .out(_U843_out)
);
assign _U844_in = _U843_out;
assign _U844_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U844 (
    .in(_U844_in),
    .clk(_U844_clk),
    .out(_U844_out)
);
assign _U845_in = _U844_out;
assign _U845_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U845 (
    .in(_U845_in),
    .clk(_U845_clk),
    .out(_U845_out)
);
assign _U846_in = _U845_out;
assign _U846_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U846 (
    .in(_U846_in),
    .clk(_U846_clk),
    .out(_U846_out)
);
assign _U847_in = _U846_out;
assign _U847_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U847 (
    .in(_U847_in),
    .clk(_U847_clk),
    .out(_U847_out)
);
assign _U848_in = _U847_out;
assign _U848_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U848 (
    .in(_U848_in),
    .clk(_U848_clk),
    .out(_U848_out)
);
assign _U849_in = _U848_out;
assign _U849_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U849 (
    .in(_U849_in),
    .clk(_U849_clk),
    .out(_U849_out)
);
assign _U850_in = _U849_out;
assign _U850_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U850 (
    .in(_U850_in),
    .clk(_U850_clk),
    .out(_U850_out)
);
assign _U851_in = _U850_out;
assign _U851_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U851 (
    .in(_U851_in),
    .clk(_U851_clk),
    .out(_U851_out)
);
assign _U852_in = _U851_out;
assign _U852_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U852 (
    .in(_U852_in),
    .clk(_U852_clk),
    .out(_U852_out)
);
assign _U853_in = _U852_out;
assign _U853_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U853 (
    .in(_U853_in),
    .clk(_U853_clk),
    .out(_U853_out)
);
assign _U854_in = _U869_out;
_U854_pt__U855 _U854 (
    .in(_U854_in),
    .out(_U854_out)
);
assign _U856_in = 16'(_U901_out * _U870_out);
assign _U856_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U856 (
    .in(_U856_in),
    .clk(_U856_clk),
    .out(_U856_out)
);
assign _U857_in = _U856_out;
assign _U857_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U857 (
    .in(_U857_in),
    .clk(_U857_clk),
    .out(_U857_out)
);
assign _U858_in = _U857_out;
assign _U858_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U858 (
    .in(_U858_in),
    .clk(_U858_clk),
    .out(_U858_out)
);
assign _U859_in = _U858_out;
assign _U859_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U859 (
    .in(_U859_in),
    .clk(_U859_clk),
    .out(_U859_out)
);
assign _U860_in = _U859_out;
assign _U860_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U860 (
    .in(_U860_in),
    .clk(_U860_clk),
    .out(_U860_out)
);
assign _U861_in = _U860_out;
assign _U861_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U861 (
    .in(_U861_in),
    .clk(_U861_clk),
    .out(_U861_out)
);
assign _U862_in = _U861_out;
assign _U862_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U862 (
    .in(_U862_in),
    .clk(_U862_clk),
    .out(_U862_out)
);
assign _U863_in = _U862_out;
assign _U863_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U863 (
    .in(_U863_in),
    .clk(_U863_clk),
    .out(_U863_out)
);
assign _U864_in = _U863_out;
assign _U864_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U864 (
    .in(_U864_in),
    .clk(_U864_clk),
    .out(_U864_out)
);
assign _U865_in = _U864_out;
assign _U865_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U865 (
    .in(_U865_in),
    .clk(_U865_clk),
    .out(_U865_out)
);
assign _U866_in = _U865_out;
assign _U866_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U866 (
    .in(_U866_in),
    .clk(_U866_clk),
    .out(_U866_out)
);
assign _U867_in = _U866_out;
assign _U867_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U867 (
    .in(_U867_in),
    .clk(_U867_clk),
    .out(_U867_out)
);
assign _U868_in = _U867_out;
assign _U868_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U868 (
    .in(_U868_in),
    .clk(_U868_clk),
    .out(_U868_out)
);
assign _U869_in = _U868_out;
assign _U869_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U869 (
    .in(_U869_in),
    .clk(_U869_clk),
    .out(_U869_out)
);
assign _U870_in = _U872_out;
_U870_pt__U871 _U870 (
    .in(_U870_in),
    .out(_U870_out)
);
assign _U872_in = in1_hw_input_global_wrapper_stencil[0];
assign _U872_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U872 (
    .in(_U872_in),
    .clk(_U872_clk),
    .out(_U872_out)
);
assign _U873_in = _U880_out;
_U873_pt__U874 _U873 (
    .in(_U873_in),
    .out(_U873_out)
);
assign _U875_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U875_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U875 (
    .in(_U875_in),
    .clk(_U875_clk),
    .out(_U875_out)
);
assign _U876_in = _U875_out;
assign _U876_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U876 (
    .in(_U876_in),
    .clk(_U876_clk),
    .out(_U876_out)
);
assign _U877_in = _U876_out;
assign _U877_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U877 (
    .in(_U877_in),
    .clk(_U877_clk),
    .out(_U877_out)
);
assign _U878_in = _U877_out;
assign _U878_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U878 (
    .in(_U878_in),
    .clk(_U878_clk),
    .out(_U878_out)
);
assign _U879_in = _U878_out;
assign _U879_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U879 (
    .in(_U879_in),
    .clk(_U879_clk),
    .out(_U879_out)
);
assign _U880_in = _U879_out;
assign _U880_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U880 (
    .in(_U880_in),
    .clk(_U880_clk),
    .out(_U880_out)
);
assign _U881_in = _U887_out;
_U881_pt__U882 _U881 (
    .in(_U881_in),
    .out(_U881_out)
);
assign _U883_in = 16'(_U941_out * _U946_out);
assign _U883_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U883 (
    .in(_U883_in),
    .clk(_U883_clk),
    .out(_U883_out)
);
assign _U884_in = _U883_out;
assign _U884_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U884 (
    .in(_U884_in),
    .clk(_U884_clk),
    .out(_U884_out)
);
assign _U885_in = _U884_out;
assign _U885_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U885 (
    .in(_U885_in),
    .clk(_U885_clk),
    .out(_U885_out)
);
assign _U886_in = _U885_out;
assign _U886_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U886 (
    .in(_U886_in),
    .clk(_U886_clk),
    .out(_U886_out)
);
assign _U887_in = _U886_out;
assign _U887_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U887 (
    .in(_U887_in),
    .clk(_U887_clk),
    .out(_U887_out)
);
assign _U888_in = _U897_out;
_U888_pt__U889 _U888 (
    .in(_U888_in),
    .out(_U888_out)
);
assign _U890_in = 16'(_U908_out * _U910_out);
assign _U890_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U890 (
    .in(_U890_in),
    .clk(_U890_clk),
    .out(_U890_out)
);
assign _U891_in = _U890_out;
assign _U891_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U891 (
    .in(_U891_in),
    .clk(_U891_clk),
    .out(_U891_out)
);
assign _U892_in = _U891_out;
assign _U892_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U892 (
    .in(_U892_in),
    .clk(_U892_clk),
    .out(_U892_out)
);
assign _U893_in = _U892_out;
assign _U893_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U893 (
    .in(_U893_in),
    .clk(_U893_clk),
    .out(_U893_out)
);
assign _U894_in = _U893_out;
assign _U894_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U894 (
    .in(_U894_in),
    .clk(_U894_clk),
    .out(_U894_out)
);
assign _U895_in = _U894_out;
assign _U895_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U895 (
    .in(_U895_in),
    .clk(_U895_clk),
    .out(_U895_out)
);
assign _U896_in = _U895_out;
assign _U896_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U896 (
    .in(_U896_in),
    .clk(_U896_clk),
    .out(_U896_out)
);
assign _U897_in = _U896_out;
assign _U897_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U897 (
    .in(_U897_in),
    .clk(_U897_clk),
    .out(_U897_out)
);
assign _U898_in = _U900_out;
_U898_pt__U899 _U898 (
    .in(_U898_in),
    .out(_U898_out)
);
assign _U900_in = 16'(_U881_out + _U888_out);
assign _U900_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U900 (
    .in(_U900_in),
    .clk(_U900_clk),
    .out(_U900_out)
);
assign _U901_in = _U903_out;
_U901_pt__U902 _U901 (
    .in(_U901_in),
    .out(_U901_out)
);
assign _U903_in = in2_hw_kernel_global_wrapper_stencil[0];
assign _U903_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U903 (
    .in(_U903_in),
    .clk(_U903_clk),
    .out(_U903_out)
);
assign _U904_in = _U907_out;
_U904_pt__U905 _U904 (
    .in(_U904_in),
    .out(_U904_out)
);
assign _U906_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U906_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U906 (
    .in(_U906_in),
    .clk(_U906_clk),
    .out(_U906_out)
);
assign _U907_in = _U906_out;
assign _U907_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U907 (
    .in(_U907_in),
    .clk(_U907_clk),
    .out(_U907_out)
);
assign _U908_in = in2_hw_kernel_global_wrapper_stencil[7];
_U908_pt__U909 _U908 (
    .in(_U908_in),
    .out(_U908_out)
);
assign _U910_in = in1_hw_input_global_wrapper_stencil[7];
_U910_pt__U911 _U910 (
    .in(_U910_in),
    .out(_U910_out)
);
assign _U912_in = _U917_out;
_U912_pt__U913 _U912 (
    .in(_U912_in),
    .out(_U912_out)
);
assign _U914_in = 16'(_U927_out * _U934_out);
assign _U914_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U914 (
    .in(_U914_in),
    .clk(_U914_clk),
    .out(_U914_out)
);
assign _U915_in = _U914_out;
assign _U915_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U915 (
    .in(_U915_in),
    .clk(_U915_clk),
    .out(_U915_out)
);
assign _U916_in = _U915_out;
assign _U916_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U916 (
    .in(_U916_in),
    .clk(_U916_clk),
    .out(_U916_out)
);
assign _U917_in = _U916_out;
assign _U917_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U917 (
    .in(_U917_in),
    .clk(_U917_clk),
    .out(_U917_out)
);
assign _U918_in = _U923_out;
_U918_pt__U919 _U918 (
    .in(_U918_in),
    .out(_U918_out)
);
assign _U920_in = in1_hw_input_global_wrapper_stencil[4];
assign _U920_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U920 (
    .in(_U920_in),
    .clk(_U920_clk),
    .out(_U920_out)
);
assign _U921_in = _U920_out;
assign _U921_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U921 (
    .in(_U921_in),
    .clk(_U921_clk),
    .out(_U921_out)
);
assign _U922_in = _U921_out;
assign _U922_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U922 (
    .in(_U922_in),
    .clk(_U922_clk),
    .out(_U922_out)
);
assign _U923_in = _U922_out;
assign _U923_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U923 (
    .in(_U923_in),
    .clk(_U923_clk),
    .out(_U923_out)
);
assign _U924_in = _U926_out;
_U924_pt__U925 _U924 (
    .in(_U924_in),
    .out(_U924_out)
);
assign _U926_in = 16'(_U1010_out + _U966_out);
assign _U926_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U926 (
    .in(_U926_in),
    .clk(_U926_clk),
    .out(_U926_out)
);
assign _U927_in = _U933_out;
_U927_pt__U928 _U927 (
    .in(_U927_in),
    .out(_U927_out)
);
assign _U929_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U929_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U929 (
    .in(_U929_in),
    .clk(_U929_clk),
    .out(_U929_out)
);
assign _U930_in = _U929_out;
assign _U930_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U930 (
    .in(_U930_in),
    .clk(_U930_clk),
    .out(_U930_out)
);
assign _U931_in = _U930_out;
assign _U931_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U931 (
    .in(_U931_in),
    .clk(_U931_clk),
    .out(_U931_out)
);
assign _U932_in = _U931_out;
assign _U932_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U932 (
    .in(_U932_in),
    .clk(_U932_clk),
    .out(_U932_out)
);
assign _U933_in = _U932_out;
assign _U933_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U933 (
    .in(_U933_in),
    .clk(_U933_clk),
    .out(_U933_out)
);
assign _U934_in = _U940_out;
_U934_pt__U935 _U934 (
    .in(_U934_in),
    .out(_U934_out)
);
assign _U936_in = in1_hw_input_global_wrapper_stencil[5];
assign _U936_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U936 (
    .in(_U936_in),
    .clk(_U936_clk),
    .out(_U936_out)
);
assign _U937_in = _U936_out;
assign _U937_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U937 (
    .in(_U937_in),
    .clk(_U937_clk),
    .out(_U937_out)
);
assign _U938_in = _U937_out;
assign _U938_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U938 (
    .in(_U938_in),
    .clk(_U938_clk),
    .out(_U938_out)
);
assign _U939_in = _U938_out;
assign _U939_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U939 (
    .in(_U939_in),
    .clk(_U939_clk),
    .out(_U939_out)
);
assign _U940_in = _U939_out;
assign _U940_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U940 (
    .in(_U940_in),
    .clk(_U940_clk),
    .out(_U940_out)
);
assign _U941_in = _U945_out;
_U941_pt__U942 _U941 (
    .in(_U941_in),
    .out(_U941_out)
);
assign _U943_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U943_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U943 (
    .in(_U943_in),
    .clk(_U943_clk),
    .out(_U943_out)
);
assign _U944_in = _U943_out;
assign _U944_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U944 (
    .in(_U944_in),
    .clk(_U944_clk),
    .out(_U944_out)
);
assign _U945_in = _U944_out;
assign _U945_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U945 (
    .in(_U945_in),
    .clk(_U945_clk),
    .out(_U945_out)
);
assign _U946_in = _U950_out;
_U946_pt__U947 _U946 (
    .in(_U946_in),
    .out(_U946_out)
);
assign _U948_in = in1_hw_input_global_wrapper_stencil[6];
assign _U948_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U948 (
    .in(_U948_in),
    .clk(_U948_clk),
    .out(_U948_out)
);
assign _U949_in = _U948_out;
assign _U949_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U949 (
    .in(_U949_in),
    .clk(_U949_clk),
    .out(_U949_out)
);
assign _U950_in = _U949_out;
assign _U950_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U950 (
    .in(_U950_in),
    .clk(_U950_clk),
    .out(_U950_out)
);
assign _U951_in = _U962_out;
_U951_pt__U952 _U951 (
    .in(_U951_in),
    .out(_U951_out)
);
assign _U953_in = 16'(_U904_out * _U1026_out);
assign _U953_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U953 (
    .in(_U953_in),
    .clk(_U953_clk),
    .out(_U953_out)
);
assign _U954_in = _U953_out;
assign _U954_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U954 (
    .in(_U954_in),
    .clk(_U954_clk),
    .out(_U954_out)
);
assign _U955_in = _U954_out;
assign _U955_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U955 (
    .in(_U955_in),
    .clk(_U955_clk),
    .out(_U955_out)
);
assign _U956_in = _U955_out;
assign _U956_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U956 (
    .in(_U956_in),
    .clk(_U956_clk),
    .out(_U956_out)
);
assign _U957_in = _U956_out;
assign _U957_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U957 (
    .in(_U957_in),
    .clk(_U957_clk),
    .out(_U957_out)
);
assign _U958_in = _U957_out;
assign _U958_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U958 (
    .in(_U958_in),
    .clk(_U958_clk),
    .out(_U958_out)
);
assign _U959_in = _U958_out;
assign _U959_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U959 (
    .in(_U959_in),
    .clk(_U959_clk),
    .out(_U959_out)
);
assign _U960_in = _U959_out;
assign _U960_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U960 (
    .in(_U960_in),
    .clk(_U960_clk),
    .out(_U960_out)
);
assign _U961_in = _U960_out;
assign _U961_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U961 (
    .in(_U961_in),
    .clk(_U961_clk),
    .out(_U961_out)
);
assign _U962_in = _U961_out;
assign _U962_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U962 (
    .in(_U962_in),
    .clk(_U962_clk),
    .out(_U962_out)
);
assign _U963_in = _U965_out;
_U963_pt__U964 _U963 (
    .in(_U963_in),
    .out(_U963_out)
);
assign _U965_in = 16'(_U996_out + _U924_out);
assign _U965_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U965 (
    .in(_U965_in),
    .clk(_U965_clk),
    .out(_U965_out)
);
assign _U966_in = _U968_out;
_U966_pt__U967 _U966 (
    .in(_U966_in),
    .out(_U966_out)
);
assign _U968_in = 16'(_U912_out + _U898_out);
assign _U968_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U968 (
    .in(_U968_in),
    .clk(_U968_clk),
    .out(_U968_out)
);
assign _U969_in = _U977_out;
_U969_pt__U970 _U969 (
    .in(_U969_in),
    .out(_U969_out)
);
assign _U971_in = 16'(_U873_out * _U1018_out);
assign _U971_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U971 (
    .in(_U971_in),
    .clk(_U971_clk),
    .out(_U971_out)
);
assign _U972_in = _U971_out;
assign _U972_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U972 (
    .in(_U972_in),
    .clk(_U972_clk),
    .out(_U972_out)
);
assign _U973_in = _U972_out;
assign _U973_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U973 (
    .in(_U973_in),
    .clk(_U973_clk),
    .out(_U973_out)
);
assign _U974_in = _U973_out;
assign _U974_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U974 (
    .in(_U974_in),
    .clk(_U974_clk),
    .out(_U974_out)
);
assign _U975_in = _U974_out;
assign _U975_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U975 (
    .in(_U975_in),
    .clk(_U975_clk),
    .out(_U975_out)
);
assign _U976_in = _U975_out;
assign _U976_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U976 (
    .in(_U976_in),
    .clk(_U976_clk),
    .out(_U976_out)
);
assign _U977_in = _U976_out;
assign _U977_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U977 (
    .in(_U977_in),
    .clk(_U977_clk),
    .out(_U977_out)
);
assign _U978_in = _U980_out;
_U978_pt__U979 _U978 (
    .in(_U978_in),
    .out(_U978_out)
);
assign _U980_in = 16'(_U951_out + _U963_out);
assign _U980_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U980 (
    .in(_U980_in),
    .clk(_U980_clk),
    .out(_U980_out)
);
assign _U981_in = _U989_out;
_U981_pt__U982 _U981 (
    .in(_U981_in),
    .out(_U981_out)
);
assign _U983_in = in1_hw_input_global_wrapper_stencil[3];
assign _U983_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U983 (
    .in(_U983_in),
    .clk(_U983_clk),
    .out(_U983_out)
);
assign _U984_in = _U983_out;
assign _U984_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U984 (
    .in(_U984_in),
    .clk(_U984_clk),
    .out(_U984_out)
);
assign _U985_in = _U984_out;
assign _U985_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U985 (
    .in(_U985_in),
    .clk(_U985_clk),
    .out(_U985_out)
);
assign _U986_in = _U985_out;
assign _U986_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U986 (
    .in(_U986_in),
    .clk(_U986_clk),
    .out(_U986_out)
);
assign _U987_in = _U986_out;
assign _U987_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U987 (
    .in(_U987_in),
    .clk(_U987_clk),
    .out(_U987_out)
);
assign _U988_in = _U987_out;
assign _U988_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U988 (
    .in(_U988_in),
    .clk(_U988_clk),
    .out(_U988_out)
);
assign _U989_in = _U988_out;
assign _U989_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U989 (
    .in(_U989_in),
    .clk(_U989_clk),
    .out(_U989_out)
);
assign _U990_in = _U995_out;
_U990_pt__U991 _U990 (
    .in(_U990_in),
    .out(_U990_out)
);
assign _U992_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U992_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U992 (
    .in(_U992_in),
    .clk(_U992_clk),
    .out(_U992_out)
);
assign _U993_in = _U992_out;
assign _U993_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U993 (
    .in(_U993_in),
    .clk(_U993_clk),
    .out(_U993_out)
);
assign _U994_in = _U993_out;
assign _U994_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U994 (
    .in(_U994_in),
    .clk(_U994_clk),
    .out(_U994_out)
);
assign _U995_in = _U994_out;
assign _U995_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U995 (
    .in(_U995_in),
    .clk(_U995_clk),
    .out(_U995_out)
);
assign _U996_in = _U1001_out;
_U996_pt__U997 _U996 (
    .in(_U996_in),
    .out(_U996_out)
);
assign _U998_in = 16'(_U1030_out * _U981_out);
assign _U998_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U998 (
    .in(_U998_in),
    .clk(_U998_clk),
    .out(_U998_out)
);
assign _U999_in = _U998_out;
assign _U999_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U999 (
    .in(_U999_in),
    .clk(_U999_clk),
    .out(_U999_out)
);
endmodule

module cu_op_hcompute_conv_stencil_12 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_12_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_12_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_12_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[0];
hcompute_conv_stencil_12_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_12_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U0_pt__U1 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
wire [15:0] _U0_in;
assign _U0_in = in0_hw_input_stencil[0];
_U0_pt__U1 _U0 (
    .in(_U0_in),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil (
    input clk,
    input [15:0] hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read[0];
hcompute_hw_input_global_wrapper_stencil_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module resnet88 (
    input clk,
    input rst_n,
    input flush,
    output hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read_en,
    input [15:0] hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read_en,
    input [15:0] hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read [0:0],
    output hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read_en,
    input [15:0] hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read [0:0],
    output hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read_en,
    input [15:0] hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read [0:0],
    output hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read_en,
    input [15:0] hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read [0:0],
    output hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read_en,
    input [15:0] hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read [0:0],
    output hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read_en,
    input [15:0] hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read [0:0],
    output hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read_en,
    input [15:0] hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read [0:0],
    output hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write_valid,
    output [15:0] hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write [0:0],
    output hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write_valid,
    output [15:0] hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write [0:0],
    output hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write_valid,
    output [15:0] hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write [0:0],
    output hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write_valid,
    output [15:0] hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write [0:0],
    output hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write_valid,
    output [15:0] hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write [0:0],
    output hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write_valid,
    output [15:0] hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write [0:0],
    output hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write_valid,
    output [15:0] hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write [0:0],
    output hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write_valid,
    output [15:0] hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write [0:0]
);
wire arr__U1004_clk;
wire [15:0] arr__U1004_in [4:0];
wire [15:0] arr__U1004_out [4:0];
wire arr__U1011_clk;
wire [15:0] arr__U1011_in [4:0];
wire [15:0] arr__U1011_out [4:0];
wire arr__U1037_clk;
wire [15:0] arr__U1037_in [4:0];
wire [15:0] arr__U1037_out [4:0];
wire arr__U1044_clk;
wire [15:0] arr__U1044_in [4:0];
wire [15:0] arr__U1044_out [4:0];
wire arr__U1051_clk;
wire [15:0] arr__U1051_in [4:0];
wire [15:0] arr__U1051_out [4:0];
wire arr__U1058_clk;
wire [15:0] arr__U1058_in [4:0];
wire [15:0] arr__U1058_out [4:0];
wire arr__U1065_clk;
wire [15:0] arr__U1065_in [4:0];
wire [15:0] arr__U1065_out [4:0];
wire arr__U1072_clk;
wire [15:0] arr__U1072_in [4:0];
wire [15:0] arr__U1072_out [4:0];
wire arr__U1079_clk;
wire [15:0] arr__U1079_in [4:0];
wire [15:0] arr__U1079_out [4:0];
wire arr__U1086_clk;
wire [15:0] arr__U1086_in [4:0];
wire [15:0] arr__U1086_out [4:0];
wire arr__U1093_clk;
wire [15:0] arr__U1093_in [4:0];
wire [15:0] arr__U1093_out [4:0];
wire arr__U1100_clk;
wire [15:0] arr__U1100_in [4:0];
wire [15:0] arr__U1100_out [4:0];
wire arr__U1107_clk;
wire [15:0] arr__U1107_in [4:0];
wire [15:0] arr__U1107_out [4:0];
wire arr__U1114_clk;
wire [15:0] arr__U1114_in [4:0];
wire [15:0] arr__U1114_out [4:0];
wire arr__U1121_clk;
wire [15:0] arr__U1121_in [4:0];
wire [15:0] arr__U1121_out [4:0];
wire arr__U1128_clk;
wire [15:0] arr__U1128_in [4:0];
wire [15:0] arr__U1128_out [4:0];
wire arr__U1135_clk;
wire [15:0] arr__U1135_in [4:0];
wire [15:0] arr__U1135_out [4:0];
wire arr__U1142_clk;
wire [15:0] arr__U1142_in [4:0];
wire [15:0] arr__U1142_out [4:0];
wire arr__U1149_clk;
wire [15:0] arr__U1149_in [4:0];
wire [15:0] arr__U1149_out [4:0];
wire arr__U1192_clk;
wire [15:0] arr__U1192_in [4:0];
wire [15:0] arr__U1192_out [4:0];
wire arr__U1199_clk;
wire [15:0] arr__U1199_in [4:0];
wire [15:0] arr__U1199_out [4:0];
wire arr__U1225_clk;
wire [15:0] arr__U1225_in [4:0];
wire [15:0] arr__U1225_out [4:0];
wire arr__U1232_clk;
wire [15:0] arr__U1232_in [4:0];
wire [15:0] arr__U1232_out [4:0];
wire arr__U1239_clk;
wire [15:0] arr__U1239_in [4:0];
wire [15:0] arr__U1239_out [4:0];
wire arr__U1246_clk;
wire [15:0] arr__U1246_in [4:0];
wire [15:0] arr__U1246_out [4:0];
wire arr__U1253_clk;
wire [15:0] arr__U1253_in [4:0];
wire [15:0] arr__U1253_out [4:0];
wire arr__U1260_clk;
wire [15:0] arr__U1260_in [4:0];
wire [15:0] arr__U1260_out [4:0];
wire arr__U1267_clk;
wire [15:0] arr__U1267_in [4:0];
wire [15:0] arr__U1267_out [4:0];
wire arr__U1274_clk;
wire [15:0] arr__U1274_in [4:0];
wire [15:0] arr__U1274_out [4:0];
wire arr__U1281_clk;
wire [15:0] arr__U1281_in [4:0];
wire [15:0] arr__U1281_out [4:0];
wire arr__U1288_clk;
wire [15:0] arr__U1288_in [4:0];
wire [15:0] arr__U1288_out [4:0];
wire arr__U1295_clk;
wire [15:0] arr__U1295_in [4:0];
wire [15:0] arr__U1295_out [4:0];
wire arr__U1302_clk;
wire [15:0] arr__U1302_in [4:0];
wire [15:0] arr__U1302_out [4:0];
wire arr__U1309_clk;
wire [15:0] arr__U1309_in [4:0];
wire [15:0] arr__U1309_out [4:0];
wire arr__U1316_clk;
wire [15:0] arr__U1316_in [4:0];
wire [15:0] arr__U1316_out [4:0];
wire arr__U1323_clk;
wire [15:0] arr__U1323_in [4:0];
wire [15:0] arr__U1323_out [4:0];
wire arr__U1330_clk;
wire [15:0] arr__U1330_in [4:0];
wire [15:0] arr__U1330_out [4:0];
wire arr__U1337_clk;
wire [15:0] arr__U1337_in [4:0];
wire [15:0] arr__U1337_out [4:0];
wire arr__U1380_clk;
wire [15:0] arr__U1380_in [4:0];
wire [15:0] arr__U1380_out [4:0];
wire arr__U1387_clk;
wire [15:0] arr__U1387_in [4:0];
wire [15:0] arr__U1387_out [4:0];
wire arr__U1413_clk;
wire [15:0] arr__U1413_in [4:0];
wire [15:0] arr__U1413_out [4:0];
wire arr__U1420_clk;
wire [15:0] arr__U1420_in [4:0];
wire [15:0] arr__U1420_out [4:0];
wire arr__U1427_clk;
wire [15:0] arr__U1427_in [4:0];
wire [15:0] arr__U1427_out [4:0];
wire arr__U1434_clk;
wire [15:0] arr__U1434_in [4:0];
wire [15:0] arr__U1434_out [4:0];
wire arr__U1441_clk;
wire [15:0] arr__U1441_in [4:0];
wire [15:0] arr__U1441_out [4:0];
wire arr__U1448_clk;
wire [15:0] arr__U1448_in [4:0];
wire [15:0] arr__U1448_out [4:0];
wire arr__U1455_clk;
wire [15:0] arr__U1455_in [4:0];
wire [15:0] arr__U1455_out [4:0];
wire arr__U1462_clk;
wire [15:0] arr__U1462_in [4:0];
wire [15:0] arr__U1462_out [4:0];
wire arr__U1469_clk;
wire [15:0] arr__U1469_in [4:0];
wire [15:0] arr__U1469_out [4:0];
wire arr__U1476_clk;
wire [15:0] arr__U1476_in [4:0];
wire [15:0] arr__U1476_out [4:0];
wire arr__U1483_clk;
wire [15:0] arr__U1483_in [4:0];
wire [15:0] arr__U1483_out [4:0];
wire arr__U1490_clk;
wire [15:0] arr__U1490_in [4:0];
wire [15:0] arr__U1490_out [4:0];
wire arr__U1497_clk;
wire [15:0] arr__U1497_in [4:0];
wire [15:0] arr__U1497_out [4:0];
wire arr__U1504_clk;
wire [15:0] arr__U1504_in [4:0];
wire [15:0] arr__U1504_out [4:0];
wire arr__U1511_clk;
wire [15:0] arr__U1511_in [4:0];
wire [15:0] arr__U1511_out [4:0];
wire arr__U1518_clk;
wire [15:0] arr__U1518_in [4:0];
wire [15:0] arr__U1518_out [4:0];
wire arr__U1525_clk;
wire [15:0] arr__U1525_in [4:0];
wire [15:0] arr__U1525_out [4:0];
wire arr__U1568_clk;
wire [15:0] arr__U1568_in [4:0];
wire [15:0] arr__U1568_out [4:0];
wire arr__U1575_clk;
wire [15:0] arr__U1575_in [4:0];
wire [15:0] arr__U1575_out [4:0];
wire arr__U1601_clk;
wire [15:0] arr__U1601_in [4:0];
wire [15:0] arr__U1601_out [4:0];
wire arr__U1608_clk;
wire [15:0] arr__U1608_in [4:0];
wire [15:0] arr__U1608_out [4:0];
wire arr__U1615_clk;
wire [15:0] arr__U1615_in [4:0];
wire [15:0] arr__U1615_out [4:0];
wire arr__U1622_clk;
wire [15:0] arr__U1622_in [4:0];
wire [15:0] arr__U1622_out [4:0];
wire arr__U1629_clk;
wire [15:0] arr__U1629_in [4:0];
wire [15:0] arr__U1629_out [4:0];
wire arr__U1636_clk;
wire [15:0] arr__U1636_in [4:0];
wire [15:0] arr__U1636_out [4:0];
wire arr__U1643_clk;
wire [15:0] arr__U1643_in [4:0];
wire [15:0] arr__U1643_out [4:0];
wire arr__U1650_clk;
wire [15:0] arr__U1650_in [4:0];
wire [15:0] arr__U1650_out [4:0];
wire arr__U1657_clk;
wire [15:0] arr__U1657_in [4:0];
wire [15:0] arr__U1657_out [4:0];
wire arr__U1664_clk;
wire [15:0] arr__U1664_in [4:0];
wire [15:0] arr__U1664_out [4:0];
wire arr__U1671_clk;
wire [15:0] arr__U1671_in [4:0];
wire [15:0] arr__U1671_out [4:0];
wire arr__U1678_clk;
wire [15:0] arr__U1678_in [4:0];
wire [15:0] arr__U1678_out [4:0];
wire arr__U1685_clk;
wire [15:0] arr__U1685_in [4:0];
wire [15:0] arr__U1685_out [4:0];
wire arr__U1692_clk;
wire [15:0] arr__U1692_in [4:0];
wire [15:0] arr__U1692_out [4:0];
wire arr__U1699_clk;
wire [15:0] arr__U1699_in [4:0];
wire [15:0] arr__U1699_out [4:0];
wire arr__U1706_clk;
wire [15:0] arr__U1706_in [4:0];
wire [15:0] arr__U1706_out [4:0];
wire arr__U1713_clk;
wire [15:0] arr__U1713_in [4:0];
wire [15:0] arr__U1713_out [4:0];
wire arr__U1756_clk;
wire [15:0] arr__U1756_in [4:0];
wire [15:0] arr__U1756_out [4:0];
wire arr__U1763_clk;
wire [15:0] arr__U1763_in [4:0];
wire [15:0] arr__U1763_out [4:0];
wire arr__U1789_clk;
wire [15:0] arr__U1789_in [4:0];
wire [15:0] arr__U1789_out [4:0];
wire arr__U1796_clk;
wire [15:0] arr__U1796_in [4:0];
wire [15:0] arr__U1796_out [4:0];
wire arr__U1803_clk;
wire [15:0] arr__U1803_in [4:0];
wire [15:0] arr__U1803_out [4:0];
wire arr__U1810_clk;
wire [15:0] arr__U1810_in [4:0];
wire [15:0] arr__U1810_out [4:0];
wire arr__U1817_clk;
wire [15:0] arr__U1817_in [4:0];
wire [15:0] arr__U1817_out [4:0];
wire arr__U1824_clk;
wire [15:0] arr__U1824_in [4:0];
wire [15:0] arr__U1824_out [4:0];
wire arr__U1831_clk;
wire [15:0] arr__U1831_in [4:0];
wire [15:0] arr__U1831_out [4:0];
wire arr__U1838_clk;
wire [15:0] arr__U1838_in [4:0];
wire [15:0] arr__U1838_out [4:0];
wire arr__U1845_clk;
wire [15:0] arr__U1845_in [4:0];
wire [15:0] arr__U1845_out [4:0];
wire arr__U1852_clk;
wire [15:0] arr__U1852_in [4:0];
wire [15:0] arr__U1852_out [4:0];
wire arr__U1859_clk;
wire [15:0] arr__U1859_in [4:0];
wire [15:0] arr__U1859_out [4:0];
wire arr__U1866_clk;
wire [15:0] arr__U1866_in [4:0];
wire [15:0] arr__U1866_out [4:0];
wire arr__U1873_clk;
wire [15:0] arr__U1873_in [4:0];
wire [15:0] arr__U1873_out [4:0];
wire arr__U1880_clk;
wire [15:0] arr__U1880_in [4:0];
wire [15:0] arr__U1880_out [4:0];
wire arr__U1887_clk;
wire [15:0] arr__U1887_in [4:0];
wire [15:0] arr__U1887_out [4:0];
wire arr__U1894_clk;
wire [15:0] arr__U1894_in [4:0];
wire [15:0] arr__U1894_out [4:0];
wire arr__U1901_clk;
wire [15:0] arr__U1901_in [4:0];
wire [15:0] arr__U1901_out [4:0];
wire arr__U1931_clk;
wire [15:0] arr__U1931_in [2:0];
wire [15:0] arr__U1931_out [2:0];
wire arr__U1936_clk;
wire [15:0] arr__U1936_in [2:0];
wire [15:0] arr__U1936_out [2:0];
wire arr__U1945_clk;
wire [15:0] arr__U1945_in [2:0];
wire [15:0] arr__U1945_out [2:0];
wire arr__U1950_clk;
wire [15:0] arr__U1950_in [2:0];
wire [15:0] arr__U1950_out [2:0];
wire arr__U1978_clk;
wire [15:0] arr__U1978_in [2:0];
wire [15:0] arr__U1978_out [2:0];
wire arr__U1983_clk;
wire [15:0] arr__U1983_in [2:0];
wire [15:0] arr__U1983_out [2:0];
wire arr__U1992_clk;
wire [15:0] arr__U1992_in [2:0];
wire [15:0] arr__U1992_out [2:0];
wire arr__U1997_clk;
wire [15:0] arr__U1997_in [2:0];
wire [15:0] arr__U1997_out [2:0];
wire arr__U2025_clk;
wire [15:0] arr__U2025_in [2:0];
wire [15:0] arr__U2025_out [2:0];
wire arr__U2030_clk;
wire [15:0] arr__U2030_in [2:0];
wire [15:0] arr__U2030_out [2:0];
wire arr__U2039_clk;
wire [15:0] arr__U2039_in [2:0];
wire [15:0] arr__U2039_out [2:0];
wire arr__U2044_clk;
wire [15:0] arr__U2044_in [2:0];
wire [15:0] arr__U2044_out [2:0];
wire arr__U2072_clk;
wire [15:0] arr__U2072_in [2:0];
wire [15:0] arr__U2072_out [2:0];
wire arr__U2077_clk;
wire [15:0] arr__U2077_in [2:0];
wire [15:0] arr__U2077_out [2:0];
wire arr__U2086_clk;
wire [15:0] arr__U2086_in [2:0];
wire [15:0] arr__U2086_out [2:0];
wire arr__U2091_clk;
wire [15:0] arr__U2091_in [2:0];
wire [15:0] arr__U2091_out [2:0];
wire arr__U2119_clk;
wire [15:0] arr__U2119_in [2:0];
wire [15:0] arr__U2119_out [2:0];
wire arr__U2124_clk;
wire [15:0] arr__U2124_in [2:0];
wire [15:0] arr__U2124_out [2:0];
wire arr__U2133_clk;
wire [15:0] arr__U2133_in [2:0];
wire [15:0] arr__U2133_out [2:0];
wire arr__U2138_clk;
wire [15:0] arr__U2138_in [2:0];
wire [15:0] arr__U2138_out [2:0];
wire arr__U2166_clk;
wire [15:0] arr__U2166_in [2:0];
wire [15:0] arr__U2166_out [2:0];
wire arr__U2171_clk;
wire [15:0] arr__U2171_in [2:0];
wire [15:0] arr__U2171_out [2:0];
wire arr__U2180_clk;
wire [15:0] arr__U2180_in [2:0];
wire [15:0] arr__U2180_out [2:0];
wire arr__U2185_clk;
wire [15:0] arr__U2185_in [2:0];
wire [15:0] arr__U2185_out [2:0];
wire arr__U2213_clk;
wire [15:0] arr__U2213_in [2:0];
wire [15:0] arr__U2213_out [2:0];
wire arr__U2218_clk;
wire [15:0] arr__U2218_in [2:0];
wire [15:0] arr__U2218_out [2:0];
wire arr__U2227_clk;
wire [15:0] arr__U2227_in [2:0];
wire [15:0] arr__U2227_out [2:0];
wire arr__U2232_clk;
wire [15:0] arr__U2232_in [2:0];
wire [15:0] arr__U2232_out [2:0];
wire arr__U2260_clk;
wire [15:0] arr__U2260_in [2:0];
wire [15:0] arr__U2260_out [2:0];
wire arr__U2265_clk;
wire [15:0] arr__U2265_in [2:0];
wire [15:0] arr__U2265_out [2:0];
wire arr__U2274_clk;
wire [15:0] arr__U2274_in [2:0];
wire [15:0] arr__U2274_out [2:0];
wire arr__U2279_clk;
wire [15:0] arr__U2279_in [2:0];
wire [15:0] arr__U2279_out [2:0];
wire arr__U440_clk;
wire [15:0] arr__U440_in [4:0];
wire [15:0] arr__U440_out [4:0];
wire arr__U447_clk;
wire [15:0] arr__U447_in [4:0];
wire [15:0] arr__U447_out [4:0];
wire arr__U473_clk;
wire [15:0] arr__U473_in [4:0];
wire [15:0] arr__U473_out [4:0];
wire arr__U480_clk;
wire [15:0] arr__U480_in [4:0];
wire [15:0] arr__U480_out [4:0];
wire arr__U487_clk;
wire [15:0] arr__U487_in [4:0];
wire [15:0] arr__U487_out [4:0];
wire arr__U494_clk;
wire [15:0] arr__U494_in [4:0];
wire [15:0] arr__U494_out [4:0];
wire arr__U501_clk;
wire [15:0] arr__U501_in [4:0];
wire [15:0] arr__U501_out [4:0];
wire arr__U508_clk;
wire [15:0] arr__U508_in [4:0];
wire [15:0] arr__U508_out [4:0];
wire arr__U515_clk;
wire [15:0] arr__U515_in [4:0];
wire [15:0] arr__U515_out [4:0];
wire arr__U522_clk;
wire [15:0] arr__U522_in [4:0];
wire [15:0] arr__U522_out [4:0];
wire arr__U529_clk;
wire [15:0] arr__U529_in [4:0];
wire [15:0] arr__U529_out [4:0];
wire arr__U536_clk;
wire [15:0] arr__U536_in [4:0];
wire [15:0] arr__U536_out [4:0];
wire arr__U543_clk;
wire [15:0] arr__U543_in [4:0];
wire [15:0] arr__U543_out [4:0];
wire arr__U550_clk;
wire [15:0] arr__U550_in [4:0];
wire [15:0] arr__U550_out [4:0];
wire arr__U557_clk;
wire [15:0] arr__U557_in [4:0];
wire [15:0] arr__U557_out [4:0];
wire arr__U564_clk;
wire [15:0] arr__U564_in [4:0];
wire [15:0] arr__U564_out [4:0];
wire arr__U571_clk;
wire [15:0] arr__U571_in [4:0];
wire [15:0] arr__U571_out [4:0];
wire arr__U578_clk;
wire [15:0] arr__U578_in [4:0];
wire [15:0] arr__U578_out [4:0];
wire arr__U585_clk;
wire [15:0] arr__U585_in [4:0];
wire [15:0] arr__U585_out [4:0];
wire arr__U628_clk;
wire [15:0] arr__U628_in [4:0];
wire [15:0] arr__U628_out [4:0];
wire arr__U635_clk;
wire [15:0] arr__U635_in [4:0];
wire [15:0] arr__U635_out [4:0];
wire arr__U661_clk;
wire [15:0] arr__U661_in [4:0];
wire [15:0] arr__U661_out [4:0];
wire arr__U668_clk;
wire [15:0] arr__U668_in [4:0];
wire [15:0] arr__U668_out [4:0];
wire arr__U675_clk;
wire [15:0] arr__U675_in [4:0];
wire [15:0] arr__U675_out [4:0];
wire arr__U682_clk;
wire [15:0] arr__U682_in [4:0];
wire [15:0] arr__U682_out [4:0];
wire arr__U689_clk;
wire [15:0] arr__U689_in [4:0];
wire [15:0] arr__U689_out [4:0];
wire arr__U696_clk;
wire [15:0] arr__U696_in [4:0];
wire [15:0] arr__U696_out [4:0];
wire arr__U703_clk;
wire [15:0] arr__U703_in [4:0];
wire [15:0] arr__U703_out [4:0];
wire arr__U710_clk;
wire [15:0] arr__U710_in [4:0];
wire [15:0] arr__U710_out [4:0];
wire arr__U717_clk;
wire [15:0] arr__U717_in [4:0];
wire [15:0] arr__U717_out [4:0];
wire arr__U724_clk;
wire [15:0] arr__U724_in [4:0];
wire [15:0] arr__U724_out [4:0];
wire arr__U731_clk;
wire [15:0] arr__U731_in [4:0];
wire [15:0] arr__U731_out [4:0];
wire arr__U738_clk;
wire [15:0] arr__U738_in [4:0];
wire [15:0] arr__U738_out [4:0];
wire arr__U745_clk;
wire [15:0] arr__U745_in [4:0];
wire [15:0] arr__U745_out [4:0];
wire arr__U752_clk;
wire [15:0] arr__U752_in [4:0];
wire [15:0] arr__U752_out [4:0];
wire arr__U759_clk;
wire [15:0] arr__U759_in [4:0];
wire [15:0] arr__U759_out [4:0];
wire arr__U766_clk;
wire [15:0] arr__U766_in [4:0];
wire [15:0] arr__U766_out [4:0];
wire arr__U773_clk;
wire [15:0] arr__U773_in [4:0];
wire [15:0] arr__U773_out [4:0];
wire arr__U816_clk;
wire [15:0] arr__U816_in [4:0];
wire [15:0] arr__U816_out [4:0];
wire arr__U823_clk;
wire [15:0] arr__U823_in [4:0];
wire [15:0] arr__U823_out [4:0];
wire arr__U849_clk;
wire [15:0] arr__U849_in [4:0];
wire [15:0] arr__U849_out [4:0];
wire arr__U856_clk;
wire [15:0] arr__U856_in [4:0];
wire [15:0] arr__U856_out [4:0];
wire arr__U863_clk;
wire [15:0] arr__U863_in [4:0];
wire [15:0] arr__U863_out [4:0];
wire arr__U870_clk;
wire [15:0] arr__U870_in [4:0];
wire [15:0] arr__U870_out [4:0];
wire arr__U877_clk;
wire [15:0] arr__U877_in [4:0];
wire [15:0] arr__U877_out [4:0];
wire arr__U884_clk;
wire [15:0] arr__U884_in [4:0];
wire [15:0] arr__U884_out [4:0];
wire arr__U891_clk;
wire [15:0] arr__U891_in [4:0];
wire [15:0] arr__U891_out [4:0];
wire arr__U898_clk;
wire [15:0] arr__U898_in [4:0];
wire [15:0] arr__U898_out [4:0];
wire arr__U905_clk;
wire [15:0] arr__U905_in [4:0];
wire [15:0] arr__U905_out [4:0];
wire arr__U912_clk;
wire [15:0] arr__U912_in [4:0];
wire [15:0] arr__U912_out [4:0];
wire arr__U919_clk;
wire [15:0] arr__U919_in [4:0];
wire [15:0] arr__U919_out [4:0];
wire arr__U926_clk;
wire [15:0] arr__U926_in [4:0];
wire [15:0] arr__U926_out [4:0];
wire arr__U933_clk;
wire [15:0] arr__U933_in [4:0];
wire [15:0] arr__U933_out [4:0];
wire arr__U940_clk;
wire [15:0] arr__U940_in [4:0];
wire [15:0] arr__U940_out [4:0];
wire arr__U947_clk;
wire [15:0] arr__U947_in [4:0];
wire [15:0] arr__U947_out [4:0];
wire arr__U954_clk;
wire [15:0] arr__U954_in [4:0];
wire [15:0] arr__U954_out [4:0];
wire arr__U961_clk;
wire [15:0] arr__U961_in [4:0];
wire [15:0] arr__U961_out [4:0];
wire conv_stencil_clk;
wire conv_stencil_flush;
wire conv_stencil_rst_n;
wire conv_stencil_op_hcompute_conv_stencil_10_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_10_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_10_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_10_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_10_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_11_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_11_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_11_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_11_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_11_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_12_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_12_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_12_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_12_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_12_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_13_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_13_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_13_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_13_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_13_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_14_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_14_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_14_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_14_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_14_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_15_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_15_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_15_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_15_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_15_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_1_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_2_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_3_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_4_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_5_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_6_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_6_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_6_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_7_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_7_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_7_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_8_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_8_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_8_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_8_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_8_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_9_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_9_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_9_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_9_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_9_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire conv_stencil_op_hcompute_hw_output_stencil_1_read_ren;
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_1_read_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_1_read [0:0];
wire conv_stencil_op_hcompute_hw_output_stencil_2_read_ren;
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_2_read_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_2_read [0:0];
wire conv_stencil_op_hcompute_hw_output_stencil_3_read_ren;
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_3_read_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_3_read [0:0];
wire conv_stencil_op_hcompute_hw_output_stencil_4_read_ren;
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_4_read_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_4_read [0:0];
wire conv_stencil_op_hcompute_hw_output_stencil_5_read_ren;
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_5_read_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_5_read [0:0];
wire conv_stencil_op_hcompute_hw_output_stencil_6_read_ren;
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_6_read_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_6_read [0:0];
wire conv_stencil_op_hcompute_hw_output_stencil_7_read_ren;
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_7_read_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_7_read [0:0];
wire conv_stencil_op_hcompute_hw_output_stencil_read_ren;
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire delay_reg__U1001_clk;
wire delay_reg__U1001_in;
wire delay_reg__U1001_out;
wire delay_reg__U1002_clk;
wire delay_reg__U1002_in;
wire delay_reg__U1002_out;
wire delay_reg__U1019_clk;
wire delay_reg__U1019_in;
wire delay_reg__U1019_out;
wire delay_reg__U1020_clk;
wire delay_reg__U1020_in;
wire delay_reg__U1020_out;
wire delay_reg__U1021_clk;
wire delay_reg__U1021_in;
wire delay_reg__U1021_out;
wire delay_reg__U1022_clk;
wire delay_reg__U1022_in;
wire delay_reg__U1022_out;
wire delay_reg__U1023_clk;
wire delay_reg__U1023_in;
wire delay_reg__U1023_out;
wire delay_reg__U1024_clk;
wire delay_reg__U1024_in;
wire delay_reg__U1024_out;
wire delay_reg__U1025_clk;
wire delay_reg__U1025_in;
wire delay_reg__U1025_out;
wire delay_reg__U1026_clk;
wire delay_reg__U1026_in;
wire delay_reg__U1026_out;
wire delay_reg__U1027_clk;
wire delay_reg__U1027_in;
wire delay_reg__U1027_out;
wire delay_reg__U1028_clk;
wire delay_reg__U1028_in;
wire delay_reg__U1028_out;
wire delay_reg__U1029_clk;
wire delay_reg__U1029_in;
wire delay_reg__U1029_out;
wire delay_reg__U1030_clk;
wire delay_reg__U1030_in;
wire delay_reg__U1030_out;
wire delay_reg__U1031_clk;
wire delay_reg__U1031_in;
wire delay_reg__U1031_out;
wire delay_reg__U1032_clk;
wire delay_reg__U1032_in;
wire delay_reg__U1032_out;
wire delay_reg__U1033_clk;
wire delay_reg__U1033_in;
wire delay_reg__U1033_out;
wire delay_reg__U1034_clk;
wire delay_reg__U1034_in;
wire delay_reg__U1034_out;
wire delay_reg__U1035_clk;
wire delay_reg__U1035_in;
wire delay_reg__U1035_out;
wire delay_reg__U1189_clk;
wire delay_reg__U1189_in;
wire delay_reg__U1189_out;
wire delay_reg__U1190_clk;
wire delay_reg__U1190_in;
wire delay_reg__U1190_out;
wire delay_reg__U1207_clk;
wire delay_reg__U1207_in;
wire delay_reg__U1207_out;
wire delay_reg__U1208_clk;
wire delay_reg__U1208_in;
wire delay_reg__U1208_out;
wire delay_reg__U1209_clk;
wire delay_reg__U1209_in;
wire delay_reg__U1209_out;
wire delay_reg__U1210_clk;
wire delay_reg__U1210_in;
wire delay_reg__U1210_out;
wire delay_reg__U1211_clk;
wire delay_reg__U1211_in;
wire delay_reg__U1211_out;
wire delay_reg__U1212_clk;
wire delay_reg__U1212_in;
wire delay_reg__U1212_out;
wire delay_reg__U1213_clk;
wire delay_reg__U1213_in;
wire delay_reg__U1213_out;
wire delay_reg__U1214_clk;
wire delay_reg__U1214_in;
wire delay_reg__U1214_out;
wire delay_reg__U1215_clk;
wire delay_reg__U1215_in;
wire delay_reg__U1215_out;
wire delay_reg__U1216_clk;
wire delay_reg__U1216_in;
wire delay_reg__U1216_out;
wire delay_reg__U1217_clk;
wire delay_reg__U1217_in;
wire delay_reg__U1217_out;
wire delay_reg__U1218_clk;
wire delay_reg__U1218_in;
wire delay_reg__U1218_out;
wire delay_reg__U1219_clk;
wire delay_reg__U1219_in;
wire delay_reg__U1219_out;
wire delay_reg__U1220_clk;
wire delay_reg__U1220_in;
wire delay_reg__U1220_out;
wire delay_reg__U1221_clk;
wire delay_reg__U1221_in;
wire delay_reg__U1221_out;
wire delay_reg__U1222_clk;
wire delay_reg__U1222_in;
wire delay_reg__U1222_out;
wire delay_reg__U1223_clk;
wire delay_reg__U1223_in;
wire delay_reg__U1223_out;
wire delay_reg__U1377_clk;
wire delay_reg__U1377_in;
wire delay_reg__U1377_out;
wire delay_reg__U1378_clk;
wire delay_reg__U1378_in;
wire delay_reg__U1378_out;
wire delay_reg__U1395_clk;
wire delay_reg__U1395_in;
wire delay_reg__U1395_out;
wire delay_reg__U1396_clk;
wire delay_reg__U1396_in;
wire delay_reg__U1396_out;
wire delay_reg__U1397_clk;
wire delay_reg__U1397_in;
wire delay_reg__U1397_out;
wire delay_reg__U1398_clk;
wire delay_reg__U1398_in;
wire delay_reg__U1398_out;
wire delay_reg__U1399_clk;
wire delay_reg__U1399_in;
wire delay_reg__U1399_out;
wire delay_reg__U1400_clk;
wire delay_reg__U1400_in;
wire delay_reg__U1400_out;
wire delay_reg__U1401_clk;
wire delay_reg__U1401_in;
wire delay_reg__U1401_out;
wire delay_reg__U1402_clk;
wire delay_reg__U1402_in;
wire delay_reg__U1402_out;
wire delay_reg__U1403_clk;
wire delay_reg__U1403_in;
wire delay_reg__U1403_out;
wire delay_reg__U1404_clk;
wire delay_reg__U1404_in;
wire delay_reg__U1404_out;
wire delay_reg__U1405_clk;
wire delay_reg__U1405_in;
wire delay_reg__U1405_out;
wire delay_reg__U1406_clk;
wire delay_reg__U1406_in;
wire delay_reg__U1406_out;
wire delay_reg__U1407_clk;
wire delay_reg__U1407_in;
wire delay_reg__U1407_out;
wire delay_reg__U1408_clk;
wire delay_reg__U1408_in;
wire delay_reg__U1408_out;
wire delay_reg__U1409_clk;
wire delay_reg__U1409_in;
wire delay_reg__U1409_out;
wire delay_reg__U1410_clk;
wire delay_reg__U1410_in;
wire delay_reg__U1410_out;
wire delay_reg__U1411_clk;
wire delay_reg__U1411_in;
wire delay_reg__U1411_out;
wire delay_reg__U1565_clk;
wire delay_reg__U1565_in;
wire delay_reg__U1565_out;
wire delay_reg__U1566_clk;
wire delay_reg__U1566_in;
wire delay_reg__U1566_out;
wire delay_reg__U1583_clk;
wire delay_reg__U1583_in;
wire delay_reg__U1583_out;
wire delay_reg__U1584_clk;
wire delay_reg__U1584_in;
wire delay_reg__U1584_out;
wire delay_reg__U1585_clk;
wire delay_reg__U1585_in;
wire delay_reg__U1585_out;
wire delay_reg__U1586_clk;
wire delay_reg__U1586_in;
wire delay_reg__U1586_out;
wire delay_reg__U1587_clk;
wire delay_reg__U1587_in;
wire delay_reg__U1587_out;
wire delay_reg__U1588_clk;
wire delay_reg__U1588_in;
wire delay_reg__U1588_out;
wire delay_reg__U1589_clk;
wire delay_reg__U1589_in;
wire delay_reg__U1589_out;
wire delay_reg__U1590_clk;
wire delay_reg__U1590_in;
wire delay_reg__U1590_out;
wire delay_reg__U1591_clk;
wire delay_reg__U1591_in;
wire delay_reg__U1591_out;
wire delay_reg__U1592_clk;
wire delay_reg__U1592_in;
wire delay_reg__U1592_out;
wire delay_reg__U1593_clk;
wire delay_reg__U1593_in;
wire delay_reg__U1593_out;
wire delay_reg__U1594_clk;
wire delay_reg__U1594_in;
wire delay_reg__U1594_out;
wire delay_reg__U1595_clk;
wire delay_reg__U1595_in;
wire delay_reg__U1595_out;
wire delay_reg__U1596_clk;
wire delay_reg__U1596_in;
wire delay_reg__U1596_out;
wire delay_reg__U1597_clk;
wire delay_reg__U1597_in;
wire delay_reg__U1597_out;
wire delay_reg__U1598_clk;
wire delay_reg__U1598_in;
wire delay_reg__U1598_out;
wire delay_reg__U1599_clk;
wire delay_reg__U1599_in;
wire delay_reg__U1599_out;
wire delay_reg__U1753_clk;
wire delay_reg__U1753_in;
wire delay_reg__U1753_out;
wire delay_reg__U1754_clk;
wire delay_reg__U1754_in;
wire delay_reg__U1754_out;
wire delay_reg__U1771_clk;
wire delay_reg__U1771_in;
wire delay_reg__U1771_out;
wire delay_reg__U1772_clk;
wire delay_reg__U1772_in;
wire delay_reg__U1772_out;
wire delay_reg__U1773_clk;
wire delay_reg__U1773_in;
wire delay_reg__U1773_out;
wire delay_reg__U1774_clk;
wire delay_reg__U1774_in;
wire delay_reg__U1774_out;
wire delay_reg__U1775_clk;
wire delay_reg__U1775_in;
wire delay_reg__U1775_out;
wire delay_reg__U1776_clk;
wire delay_reg__U1776_in;
wire delay_reg__U1776_out;
wire delay_reg__U1777_clk;
wire delay_reg__U1777_in;
wire delay_reg__U1777_out;
wire delay_reg__U1778_clk;
wire delay_reg__U1778_in;
wire delay_reg__U1778_out;
wire delay_reg__U1779_clk;
wire delay_reg__U1779_in;
wire delay_reg__U1779_out;
wire delay_reg__U1780_clk;
wire delay_reg__U1780_in;
wire delay_reg__U1780_out;
wire delay_reg__U1781_clk;
wire delay_reg__U1781_in;
wire delay_reg__U1781_out;
wire delay_reg__U1782_clk;
wire delay_reg__U1782_in;
wire delay_reg__U1782_out;
wire delay_reg__U1783_clk;
wire delay_reg__U1783_in;
wire delay_reg__U1783_out;
wire delay_reg__U1784_clk;
wire delay_reg__U1784_in;
wire delay_reg__U1784_out;
wire delay_reg__U1785_clk;
wire delay_reg__U1785_in;
wire delay_reg__U1785_out;
wire delay_reg__U1786_clk;
wire delay_reg__U1786_in;
wire delay_reg__U1786_out;
wire delay_reg__U1787_clk;
wire delay_reg__U1787_in;
wire delay_reg__U1787_out;
wire delay_reg__U1928_clk;
wire delay_reg__U1928_in;
wire delay_reg__U1928_out;
wire delay_reg__U1929_clk;
wire delay_reg__U1929_in;
wire delay_reg__U1929_out;
wire delay_reg__U1942_clk;
wire delay_reg__U1942_in;
wire delay_reg__U1942_out;
wire delay_reg__U1943_clk;
wire delay_reg__U1943_in;
wire delay_reg__U1943_out;
wire delay_reg__U1975_clk;
wire delay_reg__U1975_in;
wire delay_reg__U1975_out;
wire delay_reg__U1976_clk;
wire delay_reg__U1976_in;
wire delay_reg__U1976_out;
wire delay_reg__U1989_clk;
wire delay_reg__U1989_in;
wire delay_reg__U1989_out;
wire delay_reg__U1990_clk;
wire delay_reg__U1990_in;
wire delay_reg__U1990_out;
wire delay_reg__U2022_clk;
wire delay_reg__U2022_in;
wire delay_reg__U2022_out;
wire delay_reg__U2023_clk;
wire delay_reg__U2023_in;
wire delay_reg__U2023_out;
wire delay_reg__U2036_clk;
wire delay_reg__U2036_in;
wire delay_reg__U2036_out;
wire delay_reg__U2037_clk;
wire delay_reg__U2037_in;
wire delay_reg__U2037_out;
wire delay_reg__U2069_clk;
wire delay_reg__U2069_in;
wire delay_reg__U2069_out;
wire delay_reg__U2070_clk;
wire delay_reg__U2070_in;
wire delay_reg__U2070_out;
wire delay_reg__U2083_clk;
wire delay_reg__U2083_in;
wire delay_reg__U2083_out;
wire delay_reg__U2084_clk;
wire delay_reg__U2084_in;
wire delay_reg__U2084_out;
wire delay_reg__U2116_clk;
wire delay_reg__U2116_in;
wire delay_reg__U2116_out;
wire delay_reg__U2117_clk;
wire delay_reg__U2117_in;
wire delay_reg__U2117_out;
wire delay_reg__U2130_clk;
wire delay_reg__U2130_in;
wire delay_reg__U2130_out;
wire delay_reg__U2131_clk;
wire delay_reg__U2131_in;
wire delay_reg__U2131_out;
wire delay_reg__U2163_clk;
wire delay_reg__U2163_in;
wire delay_reg__U2163_out;
wire delay_reg__U2164_clk;
wire delay_reg__U2164_in;
wire delay_reg__U2164_out;
wire delay_reg__U2177_clk;
wire delay_reg__U2177_in;
wire delay_reg__U2177_out;
wire delay_reg__U2178_clk;
wire delay_reg__U2178_in;
wire delay_reg__U2178_out;
wire delay_reg__U2210_clk;
wire delay_reg__U2210_in;
wire delay_reg__U2210_out;
wire delay_reg__U2211_clk;
wire delay_reg__U2211_in;
wire delay_reg__U2211_out;
wire delay_reg__U2224_clk;
wire delay_reg__U2224_in;
wire delay_reg__U2224_out;
wire delay_reg__U2225_clk;
wire delay_reg__U2225_in;
wire delay_reg__U2225_out;
wire delay_reg__U2257_clk;
wire delay_reg__U2257_in;
wire delay_reg__U2257_out;
wire delay_reg__U2258_clk;
wire delay_reg__U2258_in;
wire delay_reg__U2258_out;
wire delay_reg__U2271_clk;
wire delay_reg__U2271_in;
wire delay_reg__U2271_out;
wire delay_reg__U2272_clk;
wire delay_reg__U2272_in;
wire delay_reg__U2272_out;
wire delay_reg__U437_clk;
wire delay_reg__U437_in;
wire delay_reg__U437_out;
wire delay_reg__U438_clk;
wire delay_reg__U438_in;
wire delay_reg__U438_out;
wire delay_reg__U455_clk;
wire delay_reg__U455_in;
wire delay_reg__U455_out;
wire delay_reg__U456_clk;
wire delay_reg__U456_in;
wire delay_reg__U456_out;
wire delay_reg__U457_clk;
wire delay_reg__U457_in;
wire delay_reg__U457_out;
wire delay_reg__U458_clk;
wire delay_reg__U458_in;
wire delay_reg__U458_out;
wire delay_reg__U459_clk;
wire delay_reg__U459_in;
wire delay_reg__U459_out;
wire delay_reg__U460_clk;
wire delay_reg__U460_in;
wire delay_reg__U460_out;
wire delay_reg__U461_clk;
wire delay_reg__U461_in;
wire delay_reg__U461_out;
wire delay_reg__U462_clk;
wire delay_reg__U462_in;
wire delay_reg__U462_out;
wire delay_reg__U463_clk;
wire delay_reg__U463_in;
wire delay_reg__U463_out;
wire delay_reg__U464_clk;
wire delay_reg__U464_in;
wire delay_reg__U464_out;
wire delay_reg__U465_clk;
wire delay_reg__U465_in;
wire delay_reg__U465_out;
wire delay_reg__U466_clk;
wire delay_reg__U466_in;
wire delay_reg__U466_out;
wire delay_reg__U467_clk;
wire delay_reg__U467_in;
wire delay_reg__U467_out;
wire delay_reg__U468_clk;
wire delay_reg__U468_in;
wire delay_reg__U468_out;
wire delay_reg__U469_clk;
wire delay_reg__U469_in;
wire delay_reg__U469_out;
wire delay_reg__U470_clk;
wire delay_reg__U470_in;
wire delay_reg__U470_out;
wire delay_reg__U471_clk;
wire delay_reg__U471_in;
wire delay_reg__U471_out;
wire delay_reg__U625_clk;
wire delay_reg__U625_in;
wire delay_reg__U625_out;
wire delay_reg__U626_clk;
wire delay_reg__U626_in;
wire delay_reg__U626_out;
wire delay_reg__U643_clk;
wire delay_reg__U643_in;
wire delay_reg__U643_out;
wire delay_reg__U644_clk;
wire delay_reg__U644_in;
wire delay_reg__U644_out;
wire delay_reg__U645_clk;
wire delay_reg__U645_in;
wire delay_reg__U645_out;
wire delay_reg__U646_clk;
wire delay_reg__U646_in;
wire delay_reg__U646_out;
wire delay_reg__U647_clk;
wire delay_reg__U647_in;
wire delay_reg__U647_out;
wire delay_reg__U648_clk;
wire delay_reg__U648_in;
wire delay_reg__U648_out;
wire delay_reg__U649_clk;
wire delay_reg__U649_in;
wire delay_reg__U649_out;
wire delay_reg__U650_clk;
wire delay_reg__U650_in;
wire delay_reg__U650_out;
wire delay_reg__U651_clk;
wire delay_reg__U651_in;
wire delay_reg__U651_out;
wire delay_reg__U652_clk;
wire delay_reg__U652_in;
wire delay_reg__U652_out;
wire delay_reg__U653_clk;
wire delay_reg__U653_in;
wire delay_reg__U653_out;
wire delay_reg__U654_clk;
wire delay_reg__U654_in;
wire delay_reg__U654_out;
wire delay_reg__U655_clk;
wire delay_reg__U655_in;
wire delay_reg__U655_out;
wire delay_reg__U656_clk;
wire delay_reg__U656_in;
wire delay_reg__U656_out;
wire delay_reg__U657_clk;
wire delay_reg__U657_in;
wire delay_reg__U657_out;
wire delay_reg__U658_clk;
wire delay_reg__U658_in;
wire delay_reg__U658_out;
wire delay_reg__U659_clk;
wire delay_reg__U659_in;
wire delay_reg__U659_out;
wire delay_reg__U813_clk;
wire delay_reg__U813_in;
wire delay_reg__U813_out;
wire delay_reg__U814_clk;
wire delay_reg__U814_in;
wire delay_reg__U814_out;
wire delay_reg__U831_clk;
wire delay_reg__U831_in;
wire delay_reg__U831_out;
wire delay_reg__U832_clk;
wire delay_reg__U832_in;
wire delay_reg__U832_out;
wire delay_reg__U833_clk;
wire delay_reg__U833_in;
wire delay_reg__U833_out;
wire delay_reg__U834_clk;
wire delay_reg__U834_in;
wire delay_reg__U834_out;
wire delay_reg__U835_clk;
wire delay_reg__U835_in;
wire delay_reg__U835_out;
wire delay_reg__U836_clk;
wire delay_reg__U836_in;
wire delay_reg__U836_out;
wire delay_reg__U837_clk;
wire delay_reg__U837_in;
wire delay_reg__U837_out;
wire delay_reg__U838_clk;
wire delay_reg__U838_in;
wire delay_reg__U838_out;
wire delay_reg__U839_clk;
wire delay_reg__U839_in;
wire delay_reg__U839_out;
wire delay_reg__U840_clk;
wire delay_reg__U840_in;
wire delay_reg__U840_out;
wire delay_reg__U841_clk;
wire delay_reg__U841_in;
wire delay_reg__U841_out;
wire delay_reg__U842_clk;
wire delay_reg__U842_in;
wire delay_reg__U842_out;
wire delay_reg__U843_clk;
wire delay_reg__U843_in;
wire delay_reg__U843_out;
wire delay_reg__U844_clk;
wire delay_reg__U844_in;
wire delay_reg__U844_out;
wire delay_reg__U845_clk;
wire delay_reg__U845_in;
wire delay_reg__U845_out;
wire delay_reg__U846_clk;
wire delay_reg__U846_in;
wire delay_reg__U846_out;
wire delay_reg__U847_clk;
wire delay_reg__U847_in;
wire delay_reg__U847_out;
wire hw_input_global_wrapper_stencil_clk;
wire hw_input_global_wrapper_stencil_flush;
wire hw_input_global_wrapper_stencil_rst_n;
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write_wen;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write_ctrl_vars [2:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write [0:0];
wire hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write_wen;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write_ctrl_vars [2:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write [0:0];
wire hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write_wen;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write_ctrl_vars [2:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write [0:0];
wire hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write_wen;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write_ctrl_vars [2:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write [0:0];
wire hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write_wen;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write_ctrl_vars [2:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write [0:0];
wire hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write_wen;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write_ctrl_vars [2:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write [0:0];
wire hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write_wen;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write_ctrl_vars [2:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write [0:0];
wire hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars [2:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire hw_kernel_global_wrapper_stencil_clk;
wire hw_kernel_global_wrapper_stencil_flush;
wire hw_kernel_global_wrapper_stencil_rst_n;
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_conv_stencil_clk;
wire [15:0] op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire op_hcompute_conv_stencil_1_clk;
wire [15:0] op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire op_hcompute_conv_stencil_10_clk;
wire [15:0] op_hcompute_conv_stencil_10_conv_stencil_op_hcompute_conv_stencil_10_read [0:0];
wire [15:0] op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read [7:0];
wire [15:0] op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read [7:0];
wire [15:0] op_hcompute_conv_stencil_10_conv_stencil_op_hcompute_conv_stencil_10_write [0:0];
wire op_hcompute_conv_stencil_10_exe_start_in;
wire op_hcompute_conv_stencil_10_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_10_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_10_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_10_port_controller_clk;
wire op_hcompute_conv_stencil_10_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_10_port_controller_d [4:0];
wire op_hcompute_conv_stencil_10_read_start_in;
wire op_hcompute_conv_stencil_10_read_start_out;
wire [15:0] op_hcompute_conv_stencil_10_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_10_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_10_write_start_in;
wire op_hcompute_conv_stencil_10_write_start_out;
wire [15:0] op_hcompute_conv_stencil_10_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_10_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_11_clk;
wire [15:0] op_hcompute_conv_stencil_11_conv_stencil_op_hcompute_conv_stencil_11_read [0:0];
wire [15:0] op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read [7:0];
wire [15:0] op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read [7:0];
wire [15:0] op_hcompute_conv_stencil_11_conv_stencil_op_hcompute_conv_stencil_11_write [0:0];
wire op_hcompute_conv_stencil_11_exe_start_in;
wire op_hcompute_conv_stencil_11_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_11_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_11_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_11_port_controller_clk;
wire op_hcompute_conv_stencil_11_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_11_port_controller_d [4:0];
wire op_hcompute_conv_stencil_11_read_start_in;
wire op_hcompute_conv_stencil_11_read_start_out;
wire [15:0] op_hcompute_conv_stencil_11_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_11_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_11_write_start_in;
wire op_hcompute_conv_stencil_11_write_start_out;
wire [15:0] op_hcompute_conv_stencil_11_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_11_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_12_clk;
wire [15:0] op_hcompute_conv_stencil_12_conv_stencil_op_hcompute_conv_stencil_12_read [0:0];
wire [15:0] op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read [7:0];
wire [15:0] op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read [7:0];
wire [15:0] op_hcompute_conv_stencil_12_conv_stencil_op_hcompute_conv_stencil_12_write [0:0];
wire op_hcompute_conv_stencil_12_exe_start_in;
wire op_hcompute_conv_stencil_12_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_12_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_12_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_12_port_controller_clk;
wire op_hcompute_conv_stencil_12_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_12_port_controller_d [4:0];
wire op_hcompute_conv_stencil_12_read_start_in;
wire op_hcompute_conv_stencil_12_read_start_out;
wire [15:0] op_hcompute_conv_stencil_12_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_12_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_12_write_start_in;
wire op_hcompute_conv_stencil_12_write_start_out;
wire [15:0] op_hcompute_conv_stencil_12_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_12_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_13_clk;
wire [15:0] op_hcompute_conv_stencil_13_conv_stencil_op_hcompute_conv_stencil_13_read [0:0];
wire [15:0] op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read [7:0];
wire [15:0] op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read [7:0];
wire [15:0] op_hcompute_conv_stencil_13_conv_stencil_op_hcompute_conv_stencil_13_write [0:0];
wire op_hcompute_conv_stencil_13_exe_start_in;
wire op_hcompute_conv_stencil_13_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_13_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_13_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_13_port_controller_clk;
wire op_hcompute_conv_stencil_13_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_13_port_controller_d [4:0];
wire op_hcompute_conv_stencil_13_read_start_in;
wire op_hcompute_conv_stencil_13_read_start_out;
wire [15:0] op_hcompute_conv_stencil_13_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_13_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_13_write_start_in;
wire op_hcompute_conv_stencil_13_write_start_out;
wire [15:0] op_hcompute_conv_stencil_13_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_13_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_14_clk;
wire [15:0] op_hcompute_conv_stencil_14_conv_stencil_op_hcompute_conv_stencil_14_read [0:0];
wire [15:0] op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read [7:0];
wire [15:0] op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read [7:0];
wire [15:0] op_hcompute_conv_stencil_14_conv_stencil_op_hcompute_conv_stencil_14_write [0:0];
wire op_hcompute_conv_stencil_14_exe_start_in;
wire op_hcompute_conv_stencil_14_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_14_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_14_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_14_port_controller_clk;
wire op_hcompute_conv_stencil_14_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_14_port_controller_d [4:0];
wire op_hcompute_conv_stencil_14_read_start_in;
wire op_hcompute_conv_stencil_14_read_start_out;
wire [15:0] op_hcompute_conv_stencil_14_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_14_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_14_write_start_in;
wire op_hcompute_conv_stencil_14_write_start_out;
wire [15:0] op_hcompute_conv_stencil_14_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_14_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_15_clk;
wire [15:0] op_hcompute_conv_stencil_15_conv_stencil_op_hcompute_conv_stencil_15_read [0:0];
wire [15:0] op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read [7:0];
wire [15:0] op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read [7:0];
wire [15:0] op_hcompute_conv_stencil_15_conv_stencil_op_hcompute_conv_stencil_15_write [0:0];
wire op_hcompute_conv_stencil_15_exe_start_in;
wire op_hcompute_conv_stencil_15_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_15_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_15_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_15_port_controller_clk;
wire op_hcompute_conv_stencil_15_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_15_port_controller_d [4:0];
wire op_hcompute_conv_stencil_15_read_start_in;
wire op_hcompute_conv_stencil_15_read_start_out;
wire [15:0] op_hcompute_conv_stencil_15_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_15_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_15_write_start_in;
wire op_hcompute_conv_stencil_15_write_start_out;
wire [15:0] op_hcompute_conv_stencil_15_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_15_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_1_exe_start_in;
wire op_hcompute_conv_stencil_1_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_port_controller_clk;
wire op_hcompute_conv_stencil_1_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_1_port_controller_d [2:0];
wire op_hcompute_conv_stencil_1_read_start_in;
wire op_hcompute_conv_stencil_1_read_start_out;
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_write_start_in;
wire op_hcompute_conv_stencil_1_write_start_out;
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_clk;
wire [15:0] op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire op_hcompute_conv_stencil_2_exe_start_in;
wire op_hcompute_conv_stencil_2_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_port_controller_clk;
wire op_hcompute_conv_stencil_2_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_2_port_controller_d [2:0];
wire op_hcompute_conv_stencil_2_read_start_in;
wire op_hcompute_conv_stencil_2_read_start_out;
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_write_start_in;
wire op_hcompute_conv_stencil_2_write_start_out;
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_3_clk;
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire op_hcompute_conv_stencil_3_exe_start_in;
wire op_hcompute_conv_stencil_3_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_3_port_controller_clk;
wire op_hcompute_conv_stencil_3_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_3_port_controller_d [2:0];
wire op_hcompute_conv_stencil_3_read_start_in;
wire op_hcompute_conv_stencil_3_read_start_out;
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_3_write_start_in;
wire op_hcompute_conv_stencil_3_write_start_out;
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_4_clk;
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire op_hcompute_conv_stencil_4_exe_start_in;
wire op_hcompute_conv_stencil_4_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_4_port_controller_clk;
wire op_hcompute_conv_stencil_4_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_4_port_controller_d [2:0];
wire op_hcompute_conv_stencil_4_read_start_in;
wire op_hcompute_conv_stencil_4_read_start_out;
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_4_write_start_in;
wire op_hcompute_conv_stencil_4_write_start_out;
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_5_clk;
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire op_hcompute_conv_stencil_5_exe_start_in;
wire op_hcompute_conv_stencil_5_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_5_port_controller_clk;
wire op_hcompute_conv_stencil_5_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_5_port_controller_d [2:0];
wire op_hcompute_conv_stencil_5_read_start_in;
wire op_hcompute_conv_stencil_5_read_start_out;
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_5_write_start_in;
wire op_hcompute_conv_stencil_5_write_start_out;
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_6_clk;
wire [15:0] op_hcompute_conv_stencil_6_conv_stencil_op_hcompute_conv_stencil_6_write [0:0];
wire op_hcompute_conv_stencil_6_exe_start_in;
wire op_hcompute_conv_stencil_6_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_6_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_6_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_6_port_controller_clk;
wire op_hcompute_conv_stencil_6_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_6_port_controller_d [2:0];
wire op_hcompute_conv_stencil_6_read_start_in;
wire op_hcompute_conv_stencil_6_read_start_out;
wire [15:0] op_hcompute_conv_stencil_6_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_6_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_6_write_start_in;
wire op_hcompute_conv_stencil_6_write_start_out;
wire [15:0] op_hcompute_conv_stencil_6_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_6_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_7_clk;
wire [15:0] op_hcompute_conv_stencil_7_conv_stencil_op_hcompute_conv_stencil_7_write [0:0];
wire op_hcompute_conv_stencil_7_exe_start_in;
wire op_hcompute_conv_stencil_7_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_7_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_7_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_7_port_controller_clk;
wire op_hcompute_conv_stencil_7_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_7_port_controller_d [2:0];
wire op_hcompute_conv_stencil_7_read_start_in;
wire op_hcompute_conv_stencil_7_read_start_out;
wire [15:0] op_hcompute_conv_stencil_7_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_7_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_7_write_start_in;
wire op_hcompute_conv_stencil_7_write_start_out;
wire [15:0] op_hcompute_conv_stencil_7_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_7_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_8_clk;
wire [15:0] op_hcompute_conv_stencil_8_conv_stencil_op_hcompute_conv_stencil_8_read [0:0];
wire [15:0] op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read [7:0];
wire [15:0] op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read [7:0];
wire [15:0] op_hcompute_conv_stencil_8_conv_stencil_op_hcompute_conv_stencil_8_write [0:0];
wire op_hcompute_conv_stencil_8_exe_start_in;
wire op_hcompute_conv_stencil_8_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_8_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_8_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_8_port_controller_clk;
wire op_hcompute_conv_stencil_8_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_8_port_controller_d [4:0];
wire op_hcompute_conv_stencil_8_read_start_in;
wire op_hcompute_conv_stencil_8_read_start_out;
wire [15:0] op_hcompute_conv_stencil_8_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_8_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_8_write_start_in;
wire op_hcompute_conv_stencil_8_write_start_out;
wire [15:0] op_hcompute_conv_stencil_8_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_8_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_9_clk;
wire [15:0] op_hcompute_conv_stencil_9_conv_stencil_op_hcompute_conv_stencil_9_read [0:0];
wire [15:0] op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read [7:0];
wire [15:0] op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read [7:0];
wire [15:0] op_hcompute_conv_stencil_9_conv_stencil_op_hcompute_conv_stencil_9_write [0:0];
wire op_hcompute_conv_stencil_9_exe_start_in;
wire op_hcompute_conv_stencil_9_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_9_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_9_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_9_port_controller_clk;
wire op_hcompute_conv_stencil_9_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_9_port_controller_d [4:0];
wire op_hcompute_conv_stencil_9_read_start_in;
wire op_hcompute_conv_stencil_9_read_start_out;
wire [15:0] op_hcompute_conv_stencil_9_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_9_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_9_write_start_in;
wire op_hcompute_conv_stencil_9_write_start_out;
wire [15:0] op_hcompute_conv_stencil_9_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_9_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_exe_start_in;
wire op_hcompute_conv_stencil_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_port_controller_clk;
wire op_hcompute_conv_stencil_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_port_controller_d [2:0];
wire op_hcompute_conv_stencil_read_start_in;
wire op_hcompute_conv_stencil_read_start_out;
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_write_start_in;
wire op_hcompute_conv_stencil_write_start_out;
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_clk;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_1_clk;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_clk;
wire op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_1_read_start_in;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_1_write_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_1_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_2_clk;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_clk;
wire op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_2_read_start_in;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_2_write_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_2_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_3_clk;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_clk;
wire op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_3_read_start_in;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_3_write_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_3_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_4_clk;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_clk;
wire op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_4_read_start_in;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_4_write_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_4_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_5_clk;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_clk;
wire op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_5_read_start_in;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_5_write_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_5_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_6_clk;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_clk;
wire op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_6_read_start_in;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_6_write_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_6_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_7_clk;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_clk;
wire op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_7_read_start_in;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_7_write_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_7_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk;
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_port_controller_d [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_read_start_in;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out [2:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_clk;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in;
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk;
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in;
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out [4:0];
wire op_hcompute_hw_output_stencil_clk;
wire [15:0] op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire [15:0] op_hcompute_hw_output_stencil_hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write [0:0];
wire op_hcompute_hw_output_stencil_1_clk;
wire [15:0] op_hcompute_hw_output_stencil_1_conv_stencil_op_hcompute_hw_output_stencil_1_read [0:0];
wire [15:0] op_hcompute_hw_output_stencil_1_hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write [0:0];
wire op_hcompute_hw_output_stencil_1_exe_start_in;
wire op_hcompute_hw_output_stencil_1_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_1_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_1_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_1_port_controller_clk;
wire op_hcompute_hw_output_stencil_1_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_1_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_1_read_start_in;
wire op_hcompute_hw_output_stencil_1_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_1_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_1_read_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_1_write_start_in;
wire [15:0] op_hcompute_hw_output_stencil_1_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_1_write_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_2_clk;
wire [15:0] op_hcompute_hw_output_stencil_2_conv_stencil_op_hcompute_hw_output_stencil_2_read [0:0];
wire [15:0] op_hcompute_hw_output_stencil_2_hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write [0:0];
wire op_hcompute_hw_output_stencil_2_exe_start_in;
wire op_hcompute_hw_output_stencil_2_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_2_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_2_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_2_port_controller_clk;
wire op_hcompute_hw_output_stencil_2_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_2_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_2_read_start_in;
wire op_hcompute_hw_output_stencil_2_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_2_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_2_read_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_2_write_start_in;
wire [15:0] op_hcompute_hw_output_stencil_2_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_2_write_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_3_clk;
wire [15:0] op_hcompute_hw_output_stencil_3_conv_stencil_op_hcompute_hw_output_stencil_3_read [0:0];
wire [15:0] op_hcompute_hw_output_stencil_3_hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write [0:0];
wire op_hcompute_hw_output_stencil_3_exe_start_in;
wire op_hcompute_hw_output_stencil_3_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_3_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_3_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_3_port_controller_clk;
wire op_hcompute_hw_output_stencil_3_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_3_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_3_read_start_in;
wire op_hcompute_hw_output_stencil_3_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_3_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_3_read_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_3_write_start_in;
wire [15:0] op_hcompute_hw_output_stencil_3_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_3_write_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_4_clk;
wire [15:0] op_hcompute_hw_output_stencil_4_conv_stencil_op_hcompute_hw_output_stencil_4_read [0:0];
wire [15:0] op_hcompute_hw_output_stencil_4_hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write [0:0];
wire op_hcompute_hw_output_stencil_4_exe_start_in;
wire op_hcompute_hw_output_stencil_4_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_4_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_4_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_4_port_controller_clk;
wire op_hcompute_hw_output_stencil_4_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_4_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_4_read_start_in;
wire op_hcompute_hw_output_stencil_4_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_4_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_4_read_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_4_write_start_in;
wire [15:0] op_hcompute_hw_output_stencil_4_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_4_write_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_5_clk;
wire [15:0] op_hcompute_hw_output_stencil_5_conv_stencil_op_hcompute_hw_output_stencil_5_read [0:0];
wire [15:0] op_hcompute_hw_output_stencil_5_hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write [0:0];
wire op_hcompute_hw_output_stencil_5_exe_start_in;
wire op_hcompute_hw_output_stencil_5_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_5_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_5_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_5_port_controller_clk;
wire op_hcompute_hw_output_stencil_5_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_5_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_5_read_start_in;
wire op_hcompute_hw_output_stencil_5_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_5_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_5_read_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_5_write_start_in;
wire [15:0] op_hcompute_hw_output_stencil_5_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_5_write_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_6_clk;
wire [15:0] op_hcompute_hw_output_stencil_6_conv_stencil_op_hcompute_hw_output_stencil_6_read [0:0];
wire [15:0] op_hcompute_hw_output_stencil_6_hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write [0:0];
wire op_hcompute_hw_output_stencil_6_exe_start_in;
wire op_hcompute_hw_output_stencil_6_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_6_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_6_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_6_port_controller_clk;
wire op_hcompute_hw_output_stencil_6_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_6_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_6_read_start_in;
wire op_hcompute_hw_output_stencil_6_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_6_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_6_read_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_6_write_start_in;
wire [15:0] op_hcompute_hw_output_stencil_6_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_6_write_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_7_clk;
wire [15:0] op_hcompute_hw_output_stencil_7_conv_stencil_op_hcompute_hw_output_stencil_7_read [0:0];
wire [15:0] op_hcompute_hw_output_stencil_7_hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write [0:0];
wire op_hcompute_hw_output_stencil_7_exe_start_in;
wire op_hcompute_hw_output_stencil_7_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_7_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_7_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_7_port_controller_clk;
wire op_hcompute_hw_output_stencil_7_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_7_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_7_read_start_in;
wire op_hcompute_hw_output_stencil_7_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_7_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_7_read_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_7_write_start_in;
wire [15:0] op_hcompute_hw_output_stencil_7_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_7_write_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_exe_start_in;
wire op_hcompute_hw_output_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_port_controller_clk;
wire op_hcompute_hw_output_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_port_controller_d [2:0];
wire op_hcompute_hw_output_stencil_read_start_in;
wire op_hcompute_hw_output_stencil_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_out [2:0];
wire op_hcompute_hw_output_stencil_write_start_in;
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_out [2:0];
assign arr__U1004_clk = clk;
assign arr__U1004_in[4] = op_hcompute_conv_stencil_11_port_controller_d[4];
assign arr__U1004_in[3] = op_hcompute_conv_stencil_11_port_controller_d[3];
assign arr__U1004_in[2] = op_hcompute_conv_stencil_11_port_controller_d[2];
assign arr__U1004_in[1] = op_hcompute_conv_stencil_11_port_controller_d[1];
assign arr__U1004_in[0] = op_hcompute_conv_stencil_11_port_controller_d[0];
array_delay_U1005 arr__U1004 (
    .clk(arr__U1004_clk),
    .in(arr__U1004_in),
    .out(arr__U1004_out)
);
assign arr__U1011_clk = clk;
assign arr__U1011_in[4] = arr__U1004_out[4];
assign arr__U1011_in[3] = arr__U1004_out[3];
assign arr__U1011_in[2] = arr__U1004_out[2];
assign arr__U1011_in[1] = arr__U1004_out[1];
assign arr__U1011_in[0] = arr__U1004_out[0];
array_delay_U1012 arr__U1011 (
    .clk(arr__U1011_clk),
    .in(arr__U1011_in),
    .out(arr__U1011_out)
);
assign arr__U1037_clk = clk;
assign arr__U1037_in[4] = op_hcompute_conv_stencil_11_port_controller_d[4];
assign arr__U1037_in[3] = op_hcompute_conv_stencil_11_port_controller_d[3];
assign arr__U1037_in[2] = op_hcompute_conv_stencil_11_port_controller_d[2];
assign arr__U1037_in[1] = op_hcompute_conv_stencil_11_port_controller_d[1];
assign arr__U1037_in[0] = op_hcompute_conv_stencil_11_port_controller_d[0];
array_delay_U1038 arr__U1037 (
    .clk(arr__U1037_clk),
    .in(arr__U1037_in),
    .out(arr__U1037_out)
);
assign arr__U1044_clk = clk;
assign arr__U1044_in[4] = arr__U1037_out[4];
assign arr__U1044_in[3] = arr__U1037_out[3];
assign arr__U1044_in[2] = arr__U1037_out[2];
assign arr__U1044_in[1] = arr__U1037_out[1];
assign arr__U1044_in[0] = arr__U1037_out[0];
array_delay_U1045 arr__U1044 (
    .clk(arr__U1044_clk),
    .in(arr__U1044_in),
    .out(arr__U1044_out)
);
assign arr__U1051_clk = clk;
assign arr__U1051_in[4] = arr__U1044_out[4];
assign arr__U1051_in[3] = arr__U1044_out[3];
assign arr__U1051_in[2] = arr__U1044_out[2];
assign arr__U1051_in[1] = arr__U1044_out[1];
assign arr__U1051_in[0] = arr__U1044_out[0];
array_delay_U1052 arr__U1051 (
    .clk(arr__U1051_clk),
    .in(arr__U1051_in),
    .out(arr__U1051_out)
);
assign arr__U1058_clk = clk;
assign arr__U1058_in[4] = arr__U1051_out[4];
assign arr__U1058_in[3] = arr__U1051_out[3];
assign arr__U1058_in[2] = arr__U1051_out[2];
assign arr__U1058_in[1] = arr__U1051_out[1];
assign arr__U1058_in[0] = arr__U1051_out[0];
array_delay_U1059 arr__U1058 (
    .clk(arr__U1058_clk),
    .in(arr__U1058_in),
    .out(arr__U1058_out)
);
assign arr__U1065_clk = clk;
assign arr__U1065_in[4] = arr__U1058_out[4];
assign arr__U1065_in[3] = arr__U1058_out[3];
assign arr__U1065_in[2] = arr__U1058_out[2];
assign arr__U1065_in[1] = arr__U1058_out[1];
assign arr__U1065_in[0] = arr__U1058_out[0];
array_delay_U1066 arr__U1065 (
    .clk(arr__U1065_clk),
    .in(arr__U1065_in),
    .out(arr__U1065_out)
);
assign arr__U1072_clk = clk;
assign arr__U1072_in[4] = arr__U1065_out[4];
assign arr__U1072_in[3] = arr__U1065_out[3];
assign arr__U1072_in[2] = arr__U1065_out[2];
assign arr__U1072_in[1] = arr__U1065_out[1];
assign arr__U1072_in[0] = arr__U1065_out[0];
array_delay_U1073 arr__U1072 (
    .clk(arr__U1072_clk),
    .in(arr__U1072_in),
    .out(arr__U1072_out)
);
assign arr__U1079_clk = clk;
assign arr__U1079_in[4] = arr__U1072_out[4];
assign arr__U1079_in[3] = arr__U1072_out[3];
assign arr__U1079_in[2] = arr__U1072_out[2];
assign arr__U1079_in[1] = arr__U1072_out[1];
assign arr__U1079_in[0] = arr__U1072_out[0];
array_delay_U1080 arr__U1079 (
    .clk(arr__U1079_clk),
    .in(arr__U1079_in),
    .out(arr__U1079_out)
);
assign arr__U1086_clk = clk;
assign arr__U1086_in[4] = arr__U1079_out[4];
assign arr__U1086_in[3] = arr__U1079_out[3];
assign arr__U1086_in[2] = arr__U1079_out[2];
assign arr__U1086_in[1] = arr__U1079_out[1];
assign arr__U1086_in[0] = arr__U1079_out[0];
array_delay_U1087 arr__U1086 (
    .clk(arr__U1086_clk),
    .in(arr__U1086_in),
    .out(arr__U1086_out)
);
assign arr__U1093_clk = clk;
assign arr__U1093_in[4] = arr__U1086_out[4];
assign arr__U1093_in[3] = arr__U1086_out[3];
assign arr__U1093_in[2] = arr__U1086_out[2];
assign arr__U1093_in[1] = arr__U1086_out[1];
assign arr__U1093_in[0] = arr__U1086_out[0];
array_delay_U1094 arr__U1093 (
    .clk(arr__U1093_clk),
    .in(arr__U1093_in),
    .out(arr__U1093_out)
);
assign arr__U1100_clk = clk;
assign arr__U1100_in[4] = arr__U1093_out[4];
assign arr__U1100_in[3] = arr__U1093_out[3];
assign arr__U1100_in[2] = arr__U1093_out[2];
assign arr__U1100_in[1] = arr__U1093_out[1];
assign arr__U1100_in[0] = arr__U1093_out[0];
array_delay_U1101 arr__U1100 (
    .clk(arr__U1100_clk),
    .in(arr__U1100_in),
    .out(arr__U1100_out)
);
assign arr__U1107_clk = clk;
assign arr__U1107_in[4] = arr__U1100_out[4];
assign arr__U1107_in[3] = arr__U1100_out[3];
assign arr__U1107_in[2] = arr__U1100_out[2];
assign arr__U1107_in[1] = arr__U1100_out[1];
assign arr__U1107_in[0] = arr__U1100_out[0];
array_delay_U1108 arr__U1107 (
    .clk(arr__U1107_clk),
    .in(arr__U1107_in),
    .out(arr__U1107_out)
);
assign arr__U1114_clk = clk;
assign arr__U1114_in[4] = arr__U1107_out[4];
assign arr__U1114_in[3] = arr__U1107_out[3];
assign arr__U1114_in[2] = arr__U1107_out[2];
assign arr__U1114_in[1] = arr__U1107_out[1];
assign arr__U1114_in[0] = arr__U1107_out[0];
array_delay_U1115 arr__U1114 (
    .clk(arr__U1114_clk),
    .in(arr__U1114_in),
    .out(arr__U1114_out)
);
assign arr__U1121_clk = clk;
assign arr__U1121_in[4] = arr__U1114_out[4];
assign arr__U1121_in[3] = arr__U1114_out[3];
assign arr__U1121_in[2] = arr__U1114_out[2];
assign arr__U1121_in[1] = arr__U1114_out[1];
assign arr__U1121_in[0] = arr__U1114_out[0];
array_delay_U1122 arr__U1121 (
    .clk(arr__U1121_clk),
    .in(arr__U1121_in),
    .out(arr__U1121_out)
);
assign arr__U1128_clk = clk;
assign arr__U1128_in[4] = arr__U1121_out[4];
assign arr__U1128_in[3] = arr__U1121_out[3];
assign arr__U1128_in[2] = arr__U1121_out[2];
assign arr__U1128_in[1] = arr__U1121_out[1];
assign arr__U1128_in[0] = arr__U1121_out[0];
array_delay_U1129 arr__U1128 (
    .clk(arr__U1128_clk),
    .in(arr__U1128_in),
    .out(arr__U1128_out)
);
assign arr__U1135_clk = clk;
assign arr__U1135_in[4] = arr__U1128_out[4];
assign arr__U1135_in[3] = arr__U1128_out[3];
assign arr__U1135_in[2] = arr__U1128_out[2];
assign arr__U1135_in[1] = arr__U1128_out[1];
assign arr__U1135_in[0] = arr__U1128_out[0];
array_delay_U1136 arr__U1135 (
    .clk(arr__U1135_clk),
    .in(arr__U1135_in),
    .out(arr__U1135_out)
);
assign arr__U1142_clk = clk;
assign arr__U1142_in[4] = arr__U1135_out[4];
assign arr__U1142_in[3] = arr__U1135_out[3];
assign arr__U1142_in[2] = arr__U1135_out[2];
assign arr__U1142_in[1] = arr__U1135_out[1];
assign arr__U1142_in[0] = arr__U1135_out[0];
array_delay_U1143 arr__U1142 (
    .clk(arr__U1142_clk),
    .in(arr__U1142_in),
    .out(arr__U1142_out)
);
assign arr__U1149_clk = clk;
assign arr__U1149_in[4] = arr__U1142_out[4];
assign arr__U1149_in[3] = arr__U1142_out[3];
assign arr__U1149_in[2] = arr__U1142_out[2];
assign arr__U1149_in[1] = arr__U1142_out[1];
assign arr__U1149_in[0] = arr__U1142_out[0];
array_delay_U1150 arr__U1149 (
    .clk(arr__U1149_clk),
    .in(arr__U1149_in),
    .out(arr__U1149_out)
);
assign arr__U1192_clk = clk;
assign arr__U1192_in[4] = op_hcompute_conv_stencil_12_port_controller_d[4];
assign arr__U1192_in[3] = op_hcompute_conv_stencil_12_port_controller_d[3];
assign arr__U1192_in[2] = op_hcompute_conv_stencil_12_port_controller_d[2];
assign arr__U1192_in[1] = op_hcompute_conv_stencil_12_port_controller_d[1];
assign arr__U1192_in[0] = op_hcompute_conv_stencil_12_port_controller_d[0];
array_delay_U1193 arr__U1192 (
    .clk(arr__U1192_clk),
    .in(arr__U1192_in),
    .out(arr__U1192_out)
);
assign arr__U1199_clk = clk;
assign arr__U1199_in[4] = arr__U1192_out[4];
assign arr__U1199_in[3] = arr__U1192_out[3];
assign arr__U1199_in[2] = arr__U1192_out[2];
assign arr__U1199_in[1] = arr__U1192_out[1];
assign arr__U1199_in[0] = arr__U1192_out[0];
array_delay_U1200 arr__U1199 (
    .clk(arr__U1199_clk),
    .in(arr__U1199_in),
    .out(arr__U1199_out)
);
assign arr__U1225_clk = clk;
assign arr__U1225_in[4] = op_hcompute_conv_stencil_12_port_controller_d[4];
assign arr__U1225_in[3] = op_hcompute_conv_stencil_12_port_controller_d[3];
assign arr__U1225_in[2] = op_hcompute_conv_stencil_12_port_controller_d[2];
assign arr__U1225_in[1] = op_hcompute_conv_stencil_12_port_controller_d[1];
assign arr__U1225_in[0] = op_hcompute_conv_stencil_12_port_controller_d[0];
array_delay_U1226 arr__U1225 (
    .clk(arr__U1225_clk),
    .in(arr__U1225_in),
    .out(arr__U1225_out)
);
assign arr__U1232_clk = clk;
assign arr__U1232_in[4] = arr__U1225_out[4];
assign arr__U1232_in[3] = arr__U1225_out[3];
assign arr__U1232_in[2] = arr__U1225_out[2];
assign arr__U1232_in[1] = arr__U1225_out[1];
assign arr__U1232_in[0] = arr__U1225_out[0];
array_delay_U1233 arr__U1232 (
    .clk(arr__U1232_clk),
    .in(arr__U1232_in),
    .out(arr__U1232_out)
);
assign arr__U1239_clk = clk;
assign arr__U1239_in[4] = arr__U1232_out[4];
assign arr__U1239_in[3] = arr__U1232_out[3];
assign arr__U1239_in[2] = arr__U1232_out[2];
assign arr__U1239_in[1] = arr__U1232_out[1];
assign arr__U1239_in[0] = arr__U1232_out[0];
array_delay_U1240 arr__U1239 (
    .clk(arr__U1239_clk),
    .in(arr__U1239_in),
    .out(arr__U1239_out)
);
assign arr__U1246_clk = clk;
assign arr__U1246_in[4] = arr__U1239_out[4];
assign arr__U1246_in[3] = arr__U1239_out[3];
assign arr__U1246_in[2] = arr__U1239_out[2];
assign arr__U1246_in[1] = arr__U1239_out[1];
assign arr__U1246_in[0] = arr__U1239_out[0];
array_delay_U1247 arr__U1246 (
    .clk(arr__U1246_clk),
    .in(arr__U1246_in),
    .out(arr__U1246_out)
);
assign arr__U1253_clk = clk;
assign arr__U1253_in[4] = arr__U1246_out[4];
assign arr__U1253_in[3] = arr__U1246_out[3];
assign arr__U1253_in[2] = arr__U1246_out[2];
assign arr__U1253_in[1] = arr__U1246_out[1];
assign arr__U1253_in[0] = arr__U1246_out[0];
array_delay_U1254 arr__U1253 (
    .clk(arr__U1253_clk),
    .in(arr__U1253_in),
    .out(arr__U1253_out)
);
assign arr__U1260_clk = clk;
assign arr__U1260_in[4] = arr__U1253_out[4];
assign arr__U1260_in[3] = arr__U1253_out[3];
assign arr__U1260_in[2] = arr__U1253_out[2];
assign arr__U1260_in[1] = arr__U1253_out[1];
assign arr__U1260_in[0] = arr__U1253_out[0];
array_delay_U1261 arr__U1260 (
    .clk(arr__U1260_clk),
    .in(arr__U1260_in),
    .out(arr__U1260_out)
);
assign arr__U1267_clk = clk;
assign arr__U1267_in[4] = arr__U1260_out[4];
assign arr__U1267_in[3] = arr__U1260_out[3];
assign arr__U1267_in[2] = arr__U1260_out[2];
assign arr__U1267_in[1] = arr__U1260_out[1];
assign arr__U1267_in[0] = arr__U1260_out[0];
array_delay_U1268 arr__U1267 (
    .clk(arr__U1267_clk),
    .in(arr__U1267_in),
    .out(arr__U1267_out)
);
assign arr__U1274_clk = clk;
assign arr__U1274_in[4] = arr__U1267_out[4];
assign arr__U1274_in[3] = arr__U1267_out[3];
assign arr__U1274_in[2] = arr__U1267_out[2];
assign arr__U1274_in[1] = arr__U1267_out[1];
assign arr__U1274_in[0] = arr__U1267_out[0];
array_delay_U1275 arr__U1274 (
    .clk(arr__U1274_clk),
    .in(arr__U1274_in),
    .out(arr__U1274_out)
);
assign arr__U1281_clk = clk;
assign arr__U1281_in[4] = arr__U1274_out[4];
assign arr__U1281_in[3] = arr__U1274_out[3];
assign arr__U1281_in[2] = arr__U1274_out[2];
assign arr__U1281_in[1] = arr__U1274_out[1];
assign arr__U1281_in[0] = arr__U1274_out[0];
array_delay_U1282 arr__U1281 (
    .clk(arr__U1281_clk),
    .in(arr__U1281_in),
    .out(arr__U1281_out)
);
assign arr__U1288_clk = clk;
assign arr__U1288_in[4] = arr__U1281_out[4];
assign arr__U1288_in[3] = arr__U1281_out[3];
assign arr__U1288_in[2] = arr__U1281_out[2];
assign arr__U1288_in[1] = arr__U1281_out[1];
assign arr__U1288_in[0] = arr__U1281_out[0];
array_delay_U1289 arr__U1288 (
    .clk(arr__U1288_clk),
    .in(arr__U1288_in),
    .out(arr__U1288_out)
);
assign arr__U1295_clk = clk;
assign arr__U1295_in[4] = arr__U1288_out[4];
assign arr__U1295_in[3] = arr__U1288_out[3];
assign arr__U1295_in[2] = arr__U1288_out[2];
assign arr__U1295_in[1] = arr__U1288_out[1];
assign arr__U1295_in[0] = arr__U1288_out[0];
array_delay_U1296 arr__U1295 (
    .clk(arr__U1295_clk),
    .in(arr__U1295_in),
    .out(arr__U1295_out)
);
assign arr__U1302_clk = clk;
assign arr__U1302_in[4] = arr__U1295_out[4];
assign arr__U1302_in[3] = arr__U1295_out[3];
assign arr__U1302_in[2] = arr__U1295_out[2];
assign arr__U1302_in[1] = arr__U1295_out[1];
assign arr__U1302_in[0] = arr__U1295_out[0];
array_delay_U1303 arr__U1302 (
    .clk(arr__U1302_clk),
    .in(arr__U1302_in),
    .out(arr__U1302_out)
);
assign arr__U1309_clk = clk;
assign arr__U1309_in[4] = arr__U1302_out[4];
assign arr__U1309_in[3] = arr__U1302_out[3];
assign arr__U1309_in[2] = arr__U1302_out[2];
assign arr__U1309_in[1] = arr__U1302_out[1];
assign arr__U1309_in[0] = arr__U1302_out[0];
array_delay_U1310 arr__U1309 (
    .clk(arr__U1309_clk),
    .in(arr__U1309_in),
    .out(arr__U1309_out)
);
assign arr__U1316_clk = clk;
assign arr__U1316_in[4] = arr__U1309_out[4];
assign arr__U1316_in[3] = arr__U1309_out[3];
assign arr__U1316_in[2] = arr__U1309_out[2];
assign arr__U1316_in[1] = arr__U1309_out[1];
assign arr__U1316_in[0] = arr__U1309_out[0];
array_delay_U1317 arr__U1316 (
    .clk(arr__U1316_clk),
    .in(arr__U1316_in),
    .out(arr__U1316_out)
);
assign arr__U1323_clk = clk;
assign arr__U1323_in[4] = arr__U1316_out[4];
assign arr__U1323_in[3] = arr__U1316_out[3];
assign arr__U1323_in[2] = arr__U1316_out[2];
assign arr__U1323_in[1] = arr__U1316_out[1];
assign arr__U1323_in[0] = arr__U1316_out[0];
array_delay_U1324 arr__U1323 (
    .clk(arr__U1323_clk),
    .in(arr__U1323_in),
    .out(arr__U1323_out)
);
assign arr__U1330_clk = clk;
assign arr__U1330_in[4] = arr__U1323_out[4];
assign arr__U1330_in[3] = arr__U1323_out[3];
assign arr__U1330_in[2] = arr__U1323_out[2];
assign arr__U1330_in[1] = arr__U1323_out[1];
assign arr__U1330_in[0] = arr__U1323_out[0];
array_delay_U1331 arr__U1330 (
    .clk(arr__U1330_clk),
    .in(arr__U1330_in),
    .out(arr__U1330_out)
);
assign arr__U1337_clk = clk;
assign arr__U1337_in[4] = arr__U1330_out[4];
assign arr__U1337_in[3] = arr__U1330_out[3];
assign arr__U1337_in[2] = arr__U1330_out[2];
assign arr__U1337_in[1] = arr__U1330_out[1];
assign arr__U1337_in[0] = arr__U1330_out[0];
array_delay_U1338 arr__U1337 (
    .clk(arr__U1337_clk),
    .in(arr__U1337_in),
    .out(arr__U1337_out)
);
assign arr__U1380_clk = clk;
assign arr__U1380_in[4] = op_hcompute_conv_stencil_13_port_controller_d[4];
assign arr__U1380_in[3] = op_hcompute_conv_stencil_13_port_controller_d[3];
assign arr__U1380_in[2] = op_hcompute_conv_stencil_13_port_controller_d[2];
assign arr__U1380_in[1] = op_hcompute_conv_stencil_13_port_controller_d[1];
assign arr__U1380_in[0] = op_hcompute_conv_stencil_13_port_controller_d[0];
array_delay_U1381 arr__U1380 (
    .clk(arr__U1380_clk),
    .in(arr__U1380_in),
    .out(arr__U1380_out)
);
assign arr__U1387_clk = clk;
assign arr__U1387_in[4] = arr__U1380_out[4];
assign arr__U1387_in[3] = arr__U1380_out[3];
assign arr__U1387_in[2] = arr__U1380_out[2];
assign arr__U1387_in[1] = arr__U1380_out[1];
assign arr__U1387_in[0] = arr__U1380_out[0];
array_delay_U1388 arr__U1387 (
    .clk(arr__U1387_clk),
    .in(arr__U1387_in),
    .out(arr__U1387_out)
);
assign arr__U1413_clk = clk;
assign arr__U1413_in[4] = op_hcompute_conv_stencil_13_port_controller_d[4];
assign arr__U1413_in[3] = op_hcompute_conv_stencil_13_port_controller_d[3];
assign arr__U1413_in[2] = op_hcompute_conv_stencil_13_port_controller_d[2];
assign arr__U1413_in[1] = op_hcompute_conv_stencil_13_port_controller_d[1];
assign arr__U1413_in[0] = op_hcompute_conv_stencil_13_port_controller_d[0];
array_delay_U1414 arr__U1413 (
    .clk(arr__U1413_clk),
    .in(arr__U1413_in),
    .out(arr__U1413_out)
);
assign arr__U1420_clk = clk;
assign arr__U1420_in[4] = arr__U1413_out[4];
assign arr__U1420_in[3] = arr__U1413_out[3];
assign arr__U1420_in[2] = arr__U1413_out[2];
assign arr__U1420_in[1] = arr__U1413_out[1];
assign arr__U1420_in[0] = arr__U1413_out[0];
array_delay_U1421 arr__U1420 (
    .clk(arr__U1420_clk),
    .in(arr__U1420_in),
    .out(arr__U1420_out)
);
assign arr__U1427_clk = clk;
assign arr__U1427_in[4] = arr__U1420_out[4];
assign arr__U1427_in[3] = arr__U1420_out[3];
assign arr__U1427_in[2] = arr__U1420_out[2];
assign arr__U1427_in[1] = arr__U1420_out[1];
assign arr__U1427_in[0] = arr__U1420_out[0];
array_delay_U1428 arr__U1427 (
    .clk(arr__U1427_clk),
    .in(arr__U1427_in),
    .out(arr__U1427_out)
);
assign arr__U1434_clk = clk;
assign arr__U1434_in[4] = arr__U1427_out[4];
assign arr__U1434_in[3] = arr__U1427_out[3];
assign arr__U1434_in[2] = arr__U1427_out[2];
assign arr__U1434_in[1] = arr__U1427_out[1];
assign arr__U1434_in[0] = arr__U1427_out[0];
array_delay_U1435 arr__U1434 (
    .clk(arr__U1434_clk),
    .in(arr__U1434_in),
    .out(arr__U1434_out)
);
assign arr__U1441_clk = clk;
assign arr__U1441_in[4] = arr__U1434_out[4];
assign arr__U1441_in[3] = arr__U1434_out[3];
assign arr__U1441_in[2] = arr__U1434_out[2];
assign arr__U1441_in[1] = arr__U1434_out[1];
assign arr__U1441_in[0] = arr__U1434_out[0];
array_delay_U1442 arr__U1441 (
    .clk(arr__U1441_clk),
    .in(arr__U1441_in),
    .out(arr__U1441_out)
);
assign arr__U1448_clk = clk;
assign arr__U1448_in[4] = arr__U1441_out[4];
assign arr__U1448_in[3] = arr__U1441_out[3];
assign arr__U1448_in[2] = arr__U1441_out[2];
assign arr__U1448_in[1] = arr__U1441_out[1];
assign arr__U1448_in[0] = arr__U1441_out[0];
array_delay_U1449 arr__U1448 (
    .clk(arr__U1448_clk),
    .in(arr__U1448_in),
    .out(arr__U1448_out)
);
assign arr__U1455_clk = clk;
assign arr__U1455_in[4] = arr__U1448_out[4];
assign arr__U1455_in[3] = arr__U1448_out[3];
assign arr__U1455_in[2] = arr__U1448_out[2];
assign arr__U1455_in[1] = arr__U1448_out[1];
assign arr__U1455_in[0] = arr__U1448_out[0];
array_delay_U1456 arr__U1455 (
    .clk(arr__U1455_clk),
    .in(arr__U1455_in),
    .out(arr__U1455_out)
);
assign arr__U1462_clk = clk;
assign arr__U1462_in[4] = arr__U1455_out[4];
assign arr__U1462_in[3] = arr__U1455_out[3];
assign arr__U1462_in[2] = arr__U1455_out[2];
assign arr__U1462_in[1] = arr__U1455_out[1];
assign arr__U1462_in[0] = arr__U1455_out[0];
array_delay_U1463 arr__U1462 (
    .clk(arr__U1462_clk),
    .in(arr__U1462_in),
    .out(arr__U1462_out)
);
assign arr__U1469_clk = clk;
assign arr__U1469_in[4] = arr__U1462_out[4];
assign arr__U1469_in[3] = arr__U1462_out[3];
assign arr__U1469_in[2] = arr__U1462_out[2];
assign arr__U1469_in[1] = arr__U1462_out[1];
assign arr__U1469_in[0] = arr__U1462_out[0];
array_delay_U1470 arr__U1469 (
    .clk(arr__U1469_clk),
    .in(arr__U1469_in),
    .out(arr__U1469_out)
);
assign arr__U1476_clk = clk;
assign arr__U1476_in[4] = arr__U1469_out[4];
assign arr__U1476_in[3] = arr__U1469_out[3];
assign arr__U1476_in[2] = arr__U1469_out[2];
assign arr__U1476_in[1] = arr__U1469_out[1];
assign arr__U1476_in[0] = arr__U1469_out[0];
array_delay_U1477 arr__U1476 (
    .clk(arr__U1476_clk),
    .in(arr__U1476_in),
    .out(arr__U1476_out)
);
assign arr__U1483_clk = clk;
assign arr__U1483_in[4] = arr__U1476_out[4];
assign arr__U1483_in[3] = arr__U1476_out[3];
assign arr__U1483_in[2] = arr__U1476_out[2];
assign arr__U1483_in[1] = arr__U1476_out[1];
assign arr__U1483_in[0] = arr__U1476_out[0];
array_delay_U1484 arr__U1483 (
    .clk(arr__U1483_clk),
    .in(arr__U1483_in),
    .out(arr__U1483_out)
);
assign arr__U1490_clk = clk;
assign arr__U1490_in[4] = arr__U1483_out[4];
assign arr__U1490_in[3] = arr__U1483_out[3];
assign arr__U1490_in[2] = arr__U1483_out[2];
assign arr__U1490_in[1] = arr__U1483_out[1];
assign arr__U1490_in[0] = arr__U1483_out[0];
array_delay_U1491 arr__U1490 (
    .clk(arr__U1490_clk),
    .in(arr__U1490_in),
    .out(arr__U1490_out)
);
assign arr__U1497_clk = clk;
assign arr__U1497_in[4] = arr__U1490_out[4];
assign arr__U1497_in[3] = arr__U1490_out[3];
assign arr__U1497_in[2] = arr__U1490_out[2];
assign arr__U1497_in[1] = arr__U1490_out[1];
assign arr__U1497_in[0] = arr__U1490_out[0];
array_delay_U1498 arr__U1497 (
    .clk(arr__U1497_clk),
    .in(arr__U1497_in),
    .out(arr__U1497_out)
);
assign arr__U1504_clk = clk;
assign arr__U1504_in[4] = arr__U1497_out[4];
assign arr__U1504_in[3] = arr__U1497_out[3];
assign arr__U1504_in[2] = arr__U1497_out[2];
assign arr__U1504_in[1] = arr__U1497_out[1];
assign arr__U1504_in[0] = arr__U1497_out[0];
array_delay_U1505 arr__U1504 (
    .clk(arr__U1504_clk),
    .in(arr__U1504_in),
    .out(arr__U1504_out)
);
assign arr__U1511_clk = clk;
assign arr__U1511_in[4] = arr__U1504_out[4];
assign arr__U1511_in[3] = arr__U1504_out[3];
assign arr__U1511_in[2] = arr__U1504_out[2];
assign arr__U1511_in[1] = arr__U1504_out[1];
assign arr__U1511_in[0] = arr__U1504_out[0];
array_delay_U1512 arr__U1511 (
    .clk(arr__U1511_clk),
    .in(arr__U1511_in),
    .out(arr__U1511_out)
);
assign arr__U1518_clk = clk;
assign arr__U1518_in[4] = arr__U1511_out[4];
assign arr__U1518_in[3] = arr__U1511_out[3];
assign arr__U1518_in[2] = arr__U1511_out[2];
assign arr__U1518_in[1] = arr__U1511_out[1];
assign arr__U1518_in[0] = arr__U1511_out[0];
array_delay_U1519 arr__U1518 (
    .clk(arr__U1518_clk),
    .in(arr__U1518_in),
    .out(arr__U1518_out)
);
assign arr__U1525_clk = clk;
assign arr__U1525_in[4] = arr__U1518_out[4];
assign arr__U1525_in[3] = arr__U1518_out[3];
assign arr__U1525_in[2] = arr__U1518_out[2];
assign arr__U1525_in[1] = arr__U1518_out[1];
assign arr__U1525_in[0] = arr__U1518_out[0];
array_delay_U1526 arr__U1525 (
    .clk(arr__U1525_clk),
    .in(arr__U1525_in),
    .out(arr__U1525_out)
);
assign arr__U1568_clk = clk;
assign arr__U1568_in[4] = op_hcompute_conv_stencil_14_port_controller_d[4];
assign arr__U1568_in[3] = op_hcompute_conv_stencil_14_port_controller_d[3];
assign arr__U1568_in[2] = op_hcompute_conv_stencil_14_port_controller_d[2];
assign arr__U1568_in[1] = op_hcompute_conv_stencil_14_port_controller_d[1];
assign arr__U1568_in[0] = op_hcompute_conv_stencil_14_port_controller_d[0];
array_delay_U1569 arr__U1568 (
    .clk(arr__U1568_clk),
    .in(arr__U1568_in),
    .out(arr__U1568_out)
);
assign arr__U1575_clk = clk;
assign arr__U1575_in[4] = arr__U1568_out[4];
assign arr__U1575_in[3] = arr__U1568_out[3];
assign arr__U1575_in[2] = arr__U1568_out[2];
assign arr__U1575_in[1] = arr__U1568_out[1];
assign arr__U1575_in[0] = arr__U1568_out[0];
array_delay_U1576 arr__U1575 (
    .clk(arr__U1575_clk),
    .in(arr__U1575_in),
    .out(arr__U1575_out)
);
assign arr__U1601_clk = clk;
assign arr__U1601_in[4] = op_hcompute_conv_stencil_14_port_controller_d[4];
assign arr__U1601_in[3] = op_hcompute_conv_stencil_14_port_controller_d[3];
assign arr__U1601_in[2] = op_hcompute_conv_stencil_14_port_controller_d[2];
assign arr__U1601_in[1] = op_hcompute_conv_stencil_14_port_controller_d[1];
assign arr__U1601_in[0] = op_hcompute_conv_stencil_14_port_controller_d[0];
array_delay_U1602 arr__U1601 (
    .clk(arr__U1601_clk),
    .in(arr__U1601_in),
    .out(arr__U1601_out)
);
assign arr__U1608_clk = clk;
assign arr__U1608_in[4] = arr__U1601_out[4];
assign arr__U1608_in[3] = arr__U1601_out[3];
assign arr__U1608_in[2] = arr__U1601_out[2];
assign arr__U1608_in[1] = arr__U1601_out[1];
assign arr__U1608_in[0] = arr__U1601_out[0];
array_delay_U1609 arr__U1608 (
    .clk(arr__U1608_clk),
    .in(arr__U1608_in),
    .out(arr__U1608_out)
);
assign arr__U1615_clk = clk;
assign arr__U1615_in[4] = arr__U1608_out[4];
assign arr__U1615_in[3] = arr__U1608_out[3];
assign arr__U1615_in[2] = arr__U1608_out[2];
assign arr__U1615_in[1] = arr__U1608_out[1];
assign arr__U1615_in[0] = arr__U1608_out[0];
array_delay_U1616 arr__U1615 (
    .clk(arr__U1615_clk),
    .in(arr__U1615_in),
    .out(arr__U1615_out)
);
assign arr__U1622_clk = clk;
assign arr__U1622_in[4] = arr__U1615_out[4];
assign arr__U1622_in[3] = arr__U1615_out[3];
assign arr__U1622_in[2] = arr__U1615_out[2];
assign arr__U1622_in[1] = arr__U1615_out[1];
assign arr__U1622_in[0] = arr__U1615_out[0];
array_delay_U1623 arr__U1622 (
    .clk(arr__U1622_clk),
    .in(arr__U1622_in),
    .out(arr__U1622_out)
);
assign arr__U1629_clk = clk;
assign arr__U1629_in[4] = arr__U1622_out[4];
assign arr__U1629_in[3] = arr__U1622_out[3];
assign arr__U1629_in[2] = arr__U1622_out[2];
assign arr__U1629_in[1] = arr__U1622_out[1];
assign arr__U1629_in[0] = arr__U1622_out[0];
array_delay_U1630 arr__U1629 (
    .clk(arr__U1629_clk),
    .in(arr__U1629_in),
    .out(arr__U1629_out)
);
assign arr__U1636_clk = clk;
assign arr__U1636_in[4] = arr__U1629_out[4];
assign arr__U1636_in[3] = arr__U1629_out[3];
assign arr__U1636_in[2] = arr__U1629_out[2];
assign arr__U1636_in[1] = arr__U1629_out[1];
assign arr__U1636_in[0] = arr__U1629_out[0];
array_delay_U1637 arr__U1636 (
    .clk(arr__U1636_clk),
    .in(arr__U1636_in),
    .out(arr__U1636_out)
);
assign arr__U1643_clk = clk;
assign arr__U1643_in[4] = arr__U1636_out[4];
assign arr__U1643_in[3] = arr__U1636_out[3];
assign arr__U1643_in[2] = arr__U1636_out[2];
assign arr__U1643_in[1] = arr__U1636_out[1];
assign arr__U1643_in[0] = arr__U1636_out[0];
array_delay_U1644 arr__U1643 (
    .clk(arr__U1643_clk),
    .in(arr__U1643_in),
    .out(arr__U1643_out)
);
assign arr__U1650_clk = clk;
assign arr__U1650_in[4] = arr__U1643_out[4];
assign arr__U1650_in[3] = arr__U1643_out[3];
assign arr__U1650_in[2] = arr__U1643_out[2];
assign arr__U1650_in[1] = arr__U1643_out[1];
assign arr__U1650_in[0] = arr__U1643_out[0];
array_delay_U1651 arr__U1650 (
    .clk(arr__U1650_clk),
    .in(arr__U1650_in),
    .out(arr__U1650_out)
);
assign arr__U1657_clk = clk;
assign arr__U1657_in[4] = arr__U1650_out[4];
assign arr__U1657_in[3] = arr__U1650_out[3];
assign arr__U1657_in[2] = arr__U1650_out[2];
assign arr__U1657_in[1] = arr__U1650_out[1];
assign arr__U1657_in[0] = arr__U1650_out[0];
array_delay_U1658 arr__U1657 (
    .clk(arr__U1657_clk),
    .in(arr__U1657_in),
    .out(arr__U1657_out)
);
assign arr__U1664_clk = clk;
assign arr__U1664_in[4] = arr__U1657_out[4];
assign arr__U1664_in[3] = arr__U1657_out[3];
assign arr__U1664_in[2] = arr__U1657_out[2];
assign arr__U1664_in[1] = arr__U1657_out[1];
assign arr__U1664_in[0] = arr__U1657_out[0];
array_delay_U1665 arr__U1664 (
    .clk(arr__U1664_clk),
    .in(arr__U1664_in),
    .out(arr__U1664_out)
);
assign arr__U1671_clk = clk;
assign arr__U1671_in[4] = arr__U1664_out[4];
assign arr__U1671_in[3] = arr__U1664_out[3];
assign arr__U1671_in[2] = arr__U1664_out[2];
assign arr__U1671_in[1] = arr__U1664_out[1];
assign arr__U1671_in[0] = arr__U1664_out[0];
array_delay_U1672 arr__U1671 (
    .clk(arr__U1671_clk),
    .in(arr__U1671_in),
    .out(arr__U1671_out)
);
assign arr__U1678_clk = clk;
assign arr__U1678_in[4] = arr__U1671_out[4];
assign arr__U1678_in[3] = arr__U1671_out[3];
assign arr__U1678_in[2] = arr__U1671_out[2];
assign arr__U1678_in[1] = arr__U1671_out[1];
assign arr__U1678_in[0] = arr__U1671_out[0];
array_delay_U1679 arr__U1678 (
    .clk(arr__U1678_clk),
    .in(arr__U1678_in),
    .out(arr__U1678_out)
);
assign arr__U1685_clk = clk;
assign arr__U1685_in[4] = arr__U1678_out[4];
assign arr__U1685_in[3] = arr__U1678_out[3];
assign arr__U1685_in[2] = arr__U1678_out[2];
assign arr__U1685_in[1] = arr__U1678_out[1];
assign arr__U1685_in[0] = arr__U1678_out[0];
array_delay_U1686 arr__U1685 (
    .clk(arr__U1685_clk),
    .in(arr__U1685_in),
    .out(arr__U1685_out)
);
assign arr__U1692_clk = clk;
assign arr__U1692_in[4] = arr__U1685_out[4];
assign arr__U1692_in[3] = arr__U1685_out[3];
assign arr__U1692_in[2] = arr__U1685_out[2];
assign arr__U1692_in[1] = arr__U1685_out[1];
assign arr__U1692_in[0] = arr__U1685_out[0];
array_delay_U1693 arr__U1692 (
    .clk(arr__U1692_clk),
    .in(arr__U1692_in),
    .out(arr__U1692_out)
);
assign arr__U1699_clk = clk;
assign arr__U1699_in[4] = arr__U1692_out[4];
assign arr__U1699_in[3] = arr__U1692_out[3];
assign arr__U1699_in[2] = arr__U1692_out[2];
assign arr__U1699_in[1] = arr__U1692_out[1];
assign arr__U1699_in[0] = arr__U1692_out[0];
array_delay_U1700 arr__U1699 (
    .clk(arr__U1699_clk),
    .in(arr__U1699_in),
    .out(arr__U1699_out)
);
assign arr__U1706_clk = clk;
assign arr__U1706_in[4] = arr__U1699_out[4];
assign arr__U1706_in[3] = arr__U1699_out[3];
assign arr__U1706_in[2] = arr__U1699_out[2];
assign arr__U1706_in[1] = arr__U1699_out[1];
assign arr__U1706_in[0] = arr__U1699_out[0];
array_delay_U1707 arr__U1706 (
    .clk(arr__U1706_clk),
    .in(arr__U1706_in),
    .out(arr__U1706_out)
);
assign arr__U1713_clk = clk;
assign arr__U1713_in[4] = arr__U1706_out[4];
assign arr__U1713_in[3] = arr__U1706_out[3];
assign arr__U1713_in[2] = arr__U1706_out[2];
assign arr__U1713_in[1] = arr__U1706_out[1];
assign arr__U1713_in[0] = arr__U1706_out[0];
array_delay_U1714 arr__U1713 (
    .clk(arr__U1713_clk),
    .in(arr__U1713_in),
    .out(arr__U1713_out)
);
assign arr__U1756_clk = clk;
assign arr__U1756_in[4] = op_hcompute_conv_stencil_15_port_controller_d[4];
assign arr__U1756_in[3] = op_hcompute_conv_stencil_15_port_controller_d[3];
assign arr__U1756_in[2] = op_hcompute_conv_stencil_15_port_controller_d[2];
assign arr__U1756_in[1] = op_hcompute_conv_stencil_15_port_controller_d[1];
assign arr__U1756_in[0] = op_hcompute_conv_stencil_15_port_controller_d[0];
array_delay_U1757 arr__U1756 (
    .clk(arr__U1756_clk),
    .in(arr__U1756_in),
    .out(arr__U1756_out)
);
assign arr__U1763_clk = clk;
assign arr__U1763_in[4] = arr__U1756_out[4];
assign arr__U1763_in[3] = arr__U1756_out[3];
assign arr__U1763_in[2] = arr__U1756_out[2];
assign arr__U1763_in[1] = arr__U1756_out[1];
assign arr__U1763_in[0] = arr__U1756_out[0];
array_delay_U1764 arr__U1763 (
    .clk(arr__U1763_clk),
    .in(arr__U1763_in),
    .out(arr__U1763_out)
);
assign arr__U1789_clk = clk;
assign arr__U1789_in[4] = op_hcompute_conv_stencil_15_port_controller_d[4];
assign arr__U1789_in[3] = op_hcompute_conv_stencil_15_port_controller_d[3];
assign arr__U1789_in[2] = op_hcompute_conv_stencil_15_port_controller_d[2];
assign arr__U1789_in[1] = op_hcompute_conv_stencil_15_port_controller_d[1];
assign arr__U1789_in[0] = op_hcompute_conv_stencil_15_port_controller_d[0];
array_delay_U1790 arr__U1789 (
    .clk(arr__U1789_clk),
    .in(arr__U1789_in),
    .out(arr__U1789_out)
);
assign arr__U1796_clk = clk;
assign arr__U1796_in[4] = arr__U1789_out[4];
assign arr__U1796_in[3] = arr__U1789_out[3];
assign arr__U1796_in[2] = arr__U1789_out[2];
assign arr__U1796_in[1] = arr__U1789_out[1];
assign arr__U1796_in[0] = arr__U1789_out[0];
array_delay_U1797 arr__U1796 (
    .clk(arr__U1796_clk),
    .in(arr__U1796_in),
    .out(arr__U1796_out)
);
assign arr__U1803_clk = clk;
assign arr__U1803_in[4] = arr__U1796_out[4];
assign arr__U1803_in[3] = arr__U1796_out[3];
assign arr__U1803_in[2] = arr__U1796_out[2];
assign arr__U1803_in[1] = arr__U1796_out[1];
assign arr__U1803_in[0] = arr__U1796_out[0];
array_delay_U1804 arr__U1803 (
    .clk(arr__U1803_clk),
    .in(arr__U1803_in),
    .out(arr__U1803_out)
);
assign arr__U1810_clk = clk;
assign arr__U1810_in[4] = arr__U1803_out[4];
assign arr__U1810_in[3] = arr__U1803_out[3];
assign arr__U1810_in[2] = arr__U1803_out[2];
assign arr__U1810_in[1] = arr__U1803_out[1];
assign arr__U1810_in[0] = arr__U1803_out[0];
array_delay_U1811 arr__U1810 (
    .clk(arr__U1810_clk),
    .in(arr__U1810_in),
    .out(arr__U1810_out)
);
assign arr__U1817_clk = clk;
assign arr__U1817_in[4] = arr__U1810_out[4];
assign arr__U1817_in[3] = arr__U1810_out[3];
assign arr__U1817_in[2] = arr__U1810_out[2];
assign arr__U1817_in[1] = arr__U1810_out[1];
assign arr__U1817_in[0] = arr__U1810_out[0];
array_delay_U1818 arr__U1817 (
    .clk(arr__U1817_clk),
    .in(arr__U1817_in),
    .out(arr__U1817_out)
);
assign arr__U1824_clk = clk;
assign arr__U1824_in[4] = arr__U1817_out[4];
assign arr__U1824_in[3] = arr__U1817_out[3];
assign arr__U1824_in[2] = arr__U1817_out[2];
assign arr__U1824_in[1] = arr__U1817_out[1];
assign arr__U1824_in[0] = arr__U1817_out[0];
array_delay_U1825 arr__U1824 (
    .clk(arr__U1824_clk),
    .in(arr__U1824_in),
    .out(arr__U1824_out)
);
assign arr__U1831_clk = clk;
assign arr__U1831_in[4] = arr__U1824_out[4];
assign arr__U1831_in[3] = arr__U1824_out[3];
assign arr__U1831_in[2] = arr__U1824_out[2];
assign arr__U1831_in[1] = arr__U1824_out[1];
assign arr__U1831_in[0] = arr__U1824_out[0];
array_delay_U1832 arr__U1831 (
    .clk(arr__U1831_clk),
    .in(arr__U1831_in),
    .out(arr__U1831_out)
);
assign arr__U1838_clk = clk;
assign arr__U1838_in[4] = arr__U1831_out[4];
assign arr__U1838_in[3] = arr__U1831_out[3];
assign arr__U1838_in[2] = arr__U1831_out[2];
assign arr__U1838_in[1] = arr__U1831_out[1];
assign arr__U1838_in[0] = arr__U1831_out[0];
array_delay_U1839 arr__U1838 (
    .clk(arr__U1838_clk),
    .in(arr__U1838_in),
    .out(arr__U1838_out)
);
assign arr__U1845_clk = clk;
assign arr__U1845_in[4] = arr__U1838_out[4];
assign arr__U1845_in[3] = arr__U1838_out[3];
assign arr__U1845_in[2] = arr__U1838_out[2];
assign arr__U1845_in[1] = arr__U1838_out[1];
assign arr__U1845_in[0] = arr__U1838_out[0];
array_delay_U1846 arr__U1845 (
    .clk(arr__U1845_clk),
    .in(arr__U1845_in),
    .out(arr__U1845_out)
);
assign arr__U1852_clk = clk;
assign arr__U1852_in[4] = arr__U1845_out[4];
assign arr__U1852_in[3] = arr__U1845_out[3];
assign arr__U1852_in[2] = arr__U1845_out[2];
assign arr__U1852_in[1] = arr__U1845_out[1];
assign arr__U1852_in[0] = arr__U1845_out[0];
array_delay_U1853 arr__U1852 (
    .clk(arr__U1852_clk),
    .in(arr__U1852_in),
    .out(arr__U1852_out)
);
assign arr__U1859_clk = clk;
assign arr__U1859_in[4] = arr__U1852_out[4];
assign arr__U1859_in[3] = arr__U1852_out[3];
assign arr__U1859_in[2] = arr__U1852_out[2];
assign arr__U1859_in[1] = arr__U1852_out[1];
assign arr__U1859_in[0] = arr__U1852_out[0];
array_delay_U1860 arr__U1859 (
    .clk(arr__U1859_clk),
    .in(arr__U1859_in),
    .out(arr__U1859_out)
);
assign arr__U1866_clk = clk;
assign arr__U1866_in[4] = arr__U1859_out[4];
assign arr__U1866_in[3] = arr__U1859_out[3];
assign arr__U1866_in[2] = arr__U1859_out[2];
assign arr__U1866_in[1] = arr__U1859_out[1];
assign arr__U1866_in[0] = arr__U1859_out[0];
array_delay_U1867 arr__U1866 (
    .clk(arr__U1866_clk),
    .in(arr__U1866_in),
    .out(arr__U1866_out)
);
assign arr__U1873_clk = clk;
assign arr__U1873_in[4] = arr__U1866_out[4];
assign arr__U1873_in[3] = arr__U1866_out[3];
assign arr__U1873_in[2] = arr__U1866_out[2];
assign arr__U1873_in[1] = arr__U1866_out[1];
assign arr__U1873_in[0] = arr__U1866_out[0];
array_delay_U1874 arr__U1873 (
    .clk(arr__U1873_clk),
    .in(arr__U1873_in),
    .out(arr__U1873_out)
);
assign arr__U1880_clk = clk;
assign arr__U1880_in[4] = arr__U1873_out[4];
assign arr__U1880_in[3] = arr__U1873_out[3];
assign arr__U1880_in[2] = arr__U1873_out[2];
assign arr__U1880_in[1] = arr__U1873_out[1];
assign arr__U1880_in[0] = arr__U1873_out[0];
array_delay_U1881 arr__U1880 (
    .clk(arr__U1880_clk),
    .in(arr__U1880_in),
    .out(arr__U1880_out)
);
assign arr__U1887_clk = clk;
assign arr__U1887_in[4] = arr__U1880_out[4];
assign arr__U1887_in[3] = arr__U1880_out[3];
assign arr__U1887_in[2] = arr__U1880_out[2];
assign arr__U1887_in[1] = arr__U1880_out[1];
assign arr__U1887_in[0] = arr__U1880_out[0];
array_delay_U1888 arr__U1887 (
    .clk(arr__U1887_clk),
    .in(arr__U1887_in),
    .out(arr__U1887_out)
);
assign arr__U1894_clk = clk;
assign arr__U1894_in[4] = arr__U1887_out[4];
assign arr__U1894_in[3] = arr__U1887_out[3];
assign arr__U1894_in[2] = arr__U1887_out[2];
assign arr__U1894_in[1] = arr__U1887_out[1];
assign arr__U1894_in[0] = arr__U1887_out[0];
array_delay_U1895 arr__U1894 (
    .clk(arr__U1894_clk),
    .in(arr__U1894_in),
    .out(arr__U1894_out)
);
assign arr__U1901_clk = clk;
assign arr__U1901_in[4] = arr__U1894_out[4];
assign arr__U1901_in[3] = arr__U1894_out[3];
assign arr__U1901_in[2] = arr__U1894_out[2];
assign arr__U1901_in[1] = arr__U1894_out[1];
assign arr__U1901_in[0] = arr__U1894_out[0];
array_delay_U1902 arr__U1901 (
    .clk(arr__U1901_clk),
    .in(arr__U1901_in),
    .out(arr__U1901_out)
);
assign arr__U1931_clk = clk;
assign arr__U1931_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U1931_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U1931_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U1932 arr__U1931 (
    .clk(arr__U1931_clk),
    .in(arr__U1931_in),
    .out(arr__U1931_out)
);
assign arr__U1936_clk = clk;
assign arr__U1936_in[2] = arr__U1931_out[2];
assign arr__U1936_in[1] = arr__U1931_out[1];
assign arr__U1936_in[0] = arr__U1931_out[0];
array_delay_U1937 arr__U1936 (
    .clk(arr__U1936_clk),
    .in(arr__U1936_in),
    .out(arr__U1936_out)
);
assign arr__U1945_clk = clk;
assign arr__U1945_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U1945_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U1945_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U1946 arr__U1945 (
    .clk(arr__U1945_clk),
    .in(arr__U1945_in),
    .out(arr__U1945_out)
);
assign arr__U1950_clk = clk;
assign arr__U1950_in[2] = arr__U1945_out[2];
assign arr__U1950_in[1] = arr__U1945_out[1];
assign arr__U1950_in[0] = arr__U1945_out[0];
array_delay_U1951 arr__U1950 (
    .clk(arr__U1950_clk),
    .in(arr__U1950_in),
    .out(arr__U1950_out)
);
assign arr__U1978_clk = clk;
assign arr__U1978_in[2] = op_hcompute_hw_output_stencil_1_port_controller_d[2];
assign arr__U1978_in[1] = op_hcompute_hw_output_stencil_1_port_controller_d[1];
assign arr__U1978_in[0] = op_hcompute_hw_output_stencil_1_port_controller_d[0];
array_delay_U1979 arr__U1978 (
    .clk(arr__U1978_clk),
    .in(arr__U1978_in),
    .out(arr__U1978_out)
);
assign arr__U1983_clk = clk;
assign arr__U1983_in[2] = arr__U1978_out[2];
assign arr__U1983_in[1] = arr__U1978_out[1];
assign arr__U1983_in[0] = arr__U1978_out[0];
array_delay_U1984 arr__U1983 (
    .clk(arr__U1983_clk),
    .in(arr__U1983_in),
    .out(arr__U1983_out)
);
assign arr__U1992_clk = clk;
assign arr__U1992_in[2] = op_hcompute_hw_output_stencil_1_port_controller_d[2];
assign arr__U1992_in[1] = op_hcompute_hw_output_stencil_1_port_controller_d[1];
assign arr__U1992_in[0] = op_hcompute_hw_output_stencil_1_port_controller_d[0];
array_delay_U1993 arr__U1992 (
    .clk(arr__U1992_clk),
    .in(arr__U1992_in),
    .out(arr__U1992_out)
);
assign arr__U1997_clk = clk;
assign arr__U1997_in[2] = arr__U1992_out[2];
assign arr__U1997_in[1] = arr__U1992_out[1];
assign arr__U1997_in[0] = arr__U1992_out[0];
array_delay_U1998 arr__U1997 (
    .clk(arr__U1997_clk),
    .in(arr__U1997_in),
    .out(arr__U1997_out)
);
assign arr__U2025_clk = clk;
assign arr__U2025_in[2] = op_hcompute_hw_output_stencil_2_port_controller_d[2];
assign arr__U2025_in[1] = op_hcompute_hw_output_stencil_2_port_controller_d[1];
assign arr__U2025_in[0] = op_hcompute_hw_output_stencil_2_port_controller_d[0];
array_delay_U2026 arr__U2025 (
    .clk(arr__U2025_clk),
    .in(arr__U2025_in),
    .out(arr__U2025_out)
);
assign arr__U2030_clk = clk;
assign arr__U2030_in[2] = arr__U2025_out[2];
assign arr__U2030_in[1] = arr__U2025_out[1];
assign arr__U2030_in[0] = arr__U2025_out[0];
array_delay_U2031 arr__U2030 (
    .clk(arr__U2030_clk),
    .in(arr__U2030_in),
    .out(arr__U2030_out)
);
assign arr__U2039_clk = clk;
assign arr__U2039_in[2] = op_hcompute_hw_output_stencil_2_port_controller_d[2];
assign arr__U2039_in[1] = op_hcompute_hw_output_stencil_2_port_controller_d[1];
assign arr__U2039_in[0] = op_hcompute_hw_output_stencil_2_port_controller_d[0];
array_delay_U2040 arr__U2039 (
    .clk(arr__U2039_clk),
    .in(arr__U2039_in),
    .out(arr__U2039_out)
);
assign arr__U2044_clk = clk;
assign arr__U2044_in[2] = arr__U2039_out[2];
assign arr__U2044_in[1] = arr__U2039_out[1];
assign arr__U2044_in[0] = arr__U2039_out[0];
array_delay_U2045 arr__U2044 (
    .clk(arr__U2044_clk),
    .in(arr__U2044_in),
    .out(arr__U2044_out)
);
assign arr__U2072_clk = clk;
assign arr__U2072_in[2] = op_hcompute_hw_output_stencil_3_port_controller_d[2];
assign arr__U2072_in[1] = op_hcompute_hw_output_stencil_3_port_controller_d[1];
assign arr__U2072_in[0] = op_hcompute_hw_output_stencil_3_port_controller_d[0];
array_delay_U2073 arr__U2072 (
    .clk(arr__U2072_clk),
    .in(arr__U2072_in),
    .out(arr__U2072_out)
);
assign arr__U2077_clk = clk;
assign arr__U2077_in[2] = arr__U2072_out[2];
assign arr__U2077_in[1] = arr__U2072_out[1];
assign arr__U2077_in[0] = arr__U2072_out[0];
array_delay_U2078 arr__U2077 (
    .clk(arr__U2077_clk),
    .in(arr__U2077_in),
    .out(arr__U2077_out)
);
assign arr__U2086_clk = clk;
assign arr__U2086_in[2] = op_hcompute_hw_output_stencil_3_port_controller_d[2];
assign arr__U2086_in[1] = op_hcompute_hw_output_stencil_3_port_controller_d[1];
assign arr__U2086_in[0] = op_hcompute_hw_output_stencil_3_port_controller_d[0];
array_delay_U2087 arr__U2086 (
    .clk(arr__U2086_clk),
    .in(arr__U2086_in),
    .out(arr__U2086_out)
);
assign arr__U2091_clk = clk;
assign arr__U2091_in[2] = arr__U2086_out[2];
assign arr__U2091_in[1] = arr__U2086_out[1];
assign arr__U2091_in[0] = arr__U2086_out[0];
array_delay_U2092 arr__U2091 (
    .clk(arr__U2091_clk),
    .in(arr__U2091_in),
    .out(arr__U2091_out)
);
assign arr__U2119_clk = clk;
assign arr__U2119_in[2] = op_hcompute_hw_output_stencil_4_port_controller_d[2];
assign arr__U2119_in[1] = op_hcompute_hw_output_stencil_4_port_controller_d[1];
assign arr__U2119_in[0] = op_hcompute_hw_output_stencil_4_port_controller_d[0];
array_delay_U2120 arr__U2119 (
    .clk(arr__U2119_clk),
    .in(arr__U2119_in),
    .out(arr__U2119_out)
);
assign arr__U2124_clk = clk;
assign arr__U2124_in[2] = arr__U2119_out[2];
assign arr__U2124_in[1] = arr__U2119_out[1];
assign arr__U2124_in[0] = arr__U2119_out[0];
array_delay_U2125 arr__U2124 (
    .clk(arr__U2124_clk),
    .in(arr__U2124_in),
    .out(arr__U2124_out)
);
assign arr__U2133_clk = clk;
assign arr__U2133_in[2] = op_hcompute_hw_output_stencil_4_port_controller_d[2];
assign arr__U2133_in[1] = op_hcompute_hw_output_stencil_4_port_controller_d[1];
assign arr__U2133_in[0] = op_hcompute_hw_output_stencil_4_port_controller_d[0];
array_delay_U2134 arr__U2133 (
    .clk(arr__U2133_clk),
    .in(arr__U2133_in),
    .out(arr__U2133_out)
);
assign arr__U2138_clk = clk;
assign arr__U2138_in[2] = arr__U2133_out[2];
assign arr__U2138_in[1] = arr__U2133_out[1];
assign arr__U2138_in[0] = arr__U2133_out[0];
array_delay_U2139 arr__U2138 (
    .clk(arr__U2138_clk),
    .in(arr__U2138_in),
    .out(arr__U2138_out)
);
assign arr__U2166_clk = clk;
assign arr__U2166_in[2] = op_hcompute_hw_output_stencil_5_port_controller_d[2];
assign arr__U2166_in[1] = op_hcompute_hw_output_stencil_5_port_controller_d[1];
assign arr__U2166_in[0] = op_hcompute_hw_output_stencil_5_port_controller_d[0];
array_delay_U2167 arr__U2166 (
    .clk(arr__U2166_clk),
    .in(arr__U2166_in),
    .out(arr__U2166_out)
);
assign arr__U2171_clk = clk;
assign arr__U2171_in[2] = arr__U2166_out[2];
assign arr__U2171_in[1] = arr__U2166_out[1];
assign arr__U2171_in[0] = arr__U2166_out[0];
array_delay_U2172 arr__U2171 (
    .clk(arr__U2171_clk),
    .in(arr__U2171_in),
    .out(arr__U2171_out)
);
assign arr__U2180_clk = clk;
assign arr__U2180_in[2] = op_hcompute_hw_output_stencil_5_port_controller_d[2];
assign arr__U2180_in[1] = op_hcompute_hw_output_stencil_5_port_controller_d[1];
assign arr__U2180_in[0] = op_hcompute_hw_output_stencil_5_port_controller_d[0];
array_delay_U2181 arr__U2180 (
    .clk(arr__U2180_clk),
    .in(arr__U2180_in),
    .out(arr__U2180_out)
);
assign arr__U2185_clk = clk;
assign arr__U2185_in[2] = arr__U2180_out[2];
assign arr__U2185_in[1] = arr__U2180_out[1];
assign arr__U2185_in[0] = arr__U2180_out[0];
array_delay_U2186 arr__U2185 (
    .clk(arr__U2185_clk),
    .in(arr__U2185_in),
    .out(arr__U2185_out)
);
assign arr__U2213_clk = clk;
assign arr__U2213_in[2] = op_hcompute_hw_output_stencil_6_port_controller_d[2];
assign arr__U2213_in[1] = op_hcompute_hw_output_stencil_6_port_controller_d[1];
assign arr__U2213_in[0] = op_hcompute_hw_output_stencil_6_port_controller_d[0];
array_delay_U2214 arr__U2213 (
    .clk(arr__U2213_clk),
    .in(arr__U2213_in),
    .out(arr__U2213_out)
);
assign arr__U2218_clk = clk;
assign arr__U2218_in[2] = arr__U2213_out[2];
assign arr__U2218_in[1] = arr__U2213_out[1];
assign arr__U2218_in[0] = arr__U2213_out[0];
array_delay_U2219 arr__U2218 (
    .clk(arr__U2218_clk),
    .in(arr__U2218_in),
    .out(arr__U2218_out)
);
assign arr__U2227_clk = clk;
assign arr__U2227_in[2] = op_hcompute_hw_output_stencil_6_port_controller_d[2];
assign arr__U2227_in[1] = op_hcompute_hw_output_stencil_6_port_controller_d[1];
assign arr__U2227_in[0] = op_hcompute_hw_output_stencil_6_port_controller_d[0];
array_delay_U2228 arr__U2227 (
    .clk(arr__U2227_clk),
    .in(arr__U2227_in),
    .out(arr__U2227_out)
);
assign arr__U2232_clk = clk;
assign arr__U2232_in[2] = arr__U2227_out[2];
assign arr__U2232_in[1] = arr__U2227_out[1];
assign arr__U2232_in[0] = arr__U2227_out[0];
array_delay_U2233 arr__U2232 (
    .clk(arr__U2232_clk),
    .in(arr__U2232_in),
    .out(arr__U2232_out)
);
assign arr__U2260_clk = clk;
assign arr__U2260_in[2] = op_hcompute_hw_output_stencil_7_port_controller_d[2];
assign arr__U2260_in[1] = op_hcompute_hw_output_stencil_7_port_controller_d[1];
assign arr__U2260_in[0] = op_hcompute_hw_output_stencil_7_port_controller_d[0];
array_delay_U2261 arr__U2260 (
    .clk(arr__U2260_clk),
    .in(arr__U2260_in),
    .out(arr__U2260_out)
);
assign arr__U2265_clk = clk;
assign arr__U2265_in[2] = arr__U2260_out[2];
assign arr__U2265_in[1] = arr__U2260_out[1];
assign arr__U2265_in[0] = arr__U2260_out[0];
array_delay_U2266 arr__U2265 (
    .clk(arr__U2265_clk),
    .in(arr__U2265_in),
    .out(arr__U2265_out)
);
assign arr__U2274_clk = clk;
assign arr__U2274_in[2] = op_hcompute_hw_output_stencil_7_port_controller_d[2];
assign arr__U2274_in[1] = op_hcompute_hw_output_stencil_7_port_controller_d[1];
assign arr__U2274_in[0] = op_hcompute_hw_output_stencil_7_port_controller_d[0];
array_delay_U2275 arr__U2274 (
    .clk(arr__U2274_clk),
    .in(arr__U2274_in),
    .out(arr__U2274_out)
);
assign arr__U2279_clk = clk;
assign arr__U2279_in[2] = arr__U2274_out[2];
assign arr__U2279_in[1] = arr__U2274_out[1];
assign arr__U2279_in[0] = arr__U2274_out[0];
array_delay_U2280 arr__U2279 (
    .clk(arr__U2279_clk),
    .in(arr__U2279_in),
    .out(arr__U2279_out)
);
assign arr__U440_clk = clk;
assign arr__U440_in[4] = op_hcompute_conv_stencil_8_port_controller_d[4];
assign arr__U440_in[3] = op_hcompute_conv_stencil_8_port_controller_d[3];
assign arr__U440_in[2] = op_hcompute_conv_stencil_8_port_controller_d[2];
assign arr__U440_in[1] = op_hcompute_conv_stencil_8_port_controller_d[1];
assign arr__U440_in[0] = op_hcompute_conv_stencil_8_port_controller_d[0];
array_delay_U441 arr__U440 (
    .clk(arr__U440_clk),
    .in(arr__U440_in),
    .out(arr__U440_out)
);
assign arr__U447_clk = clk;
assign arr__U447_in[4] = arr__U440_out[4];
assign arr__U447_in[3] = arr__U440_out[3];
assign arr__U447_in[2] = arr__U440_out[2];
assign arr__U447_in[1] = arr__U440_out[1];
assign arr__U447_in[0] = arr__U440_out[0];
array_delay_U448 arr__U447 (
    .clk(arr__U447_clk),
    .in(arr__U447_in),
    .out(arr__U447_out)
);
assign arr__U473_clk = clk;
assign arr__U473_in[4] = op_hcompute_conv_stencil_8_port_controller_d[4];
assign arr__U473_in[3] = op_hcompute_conv_stencil_8_port_controller_d[3];
assign arr__U473_in[2] = op_hcompute_conv_stencil_8_port_controller_d[2];
assign arr__U473_in[1] = op_hcompute_conv_stencil_8_port_controller_d[1];
assign arr__U473_in[0] = op_hcompute_conv_stencil_8_port_controller_d[0];
array_delay_U474 arr__U473 (
    .clk(arr__U473_clk),
    .in(arr__U473_in),
    .out(arr__U473_out)
);
assign arr__U480_clk = clk;
assign arr__U480_in[4] = arr__U473_out[4];
assign arr__U480_in[3] = arr__U473_out[3];
assign arr__U480_in[2] = arr__U473_out[2];
assign arr__U480_in[1] = arr__U473_out[1];
assign arr__U480_in[0] = arr__U473_out[0];
array_delay_U481 arr__U480 (
    .clk(arr__U480_clk),
    .in(arr__U480_in),
    .out(arr__U480_out)
);
assign arr__U487_clk = clk;
assign arr__U487_in[4] = arr__U480_out[4];
assign arr__U487_in[3] = arr__U480_out[3];
assign arr__U487_in[2] = arr__U480_out[2];
assign arr__U487_in[1] = arr__U480_out[1];
assign arr__U487_in[0] = arr__U480_out[0];
array_delay_U488 arr__U487 (
    .clk(arr__U487_clk),
    .in(arr__U487_in),
    .out(arr__U487_out)
);
assign arr__U494_clk = clk;
assign arr__U494_in[4] = arr__U487_out[4];
assign arr__U494_in[3] = arr__U487_out[3];
assign arr__U494_in[2] = arr__U487_out[2];
assign arr__U494_in[1] = arr__U487_out[1];
assign arr__U494_in[0] = arr__U487_out[0];
array_delay_U495 arr__U494 (
    .clk(arr__U494_clk),
    .in(arr__U494_in),
    .out(arr__U494_out)
);
assign arr__U501_clk = clk;
assign arr__U501_in[4] = arr__U494_out[4];
assign arr__U501_in[3] = arr__U494_out[3];
assign arr__U501_in[2] = arr__U494_out[2];
assign arr__U501_in[1] = arr__U494_out[1];
assign arr__U501_in[0] = arr__U494_out[0];
array_delay_U502 arr__U501 (
    .clk(arr__U501_clk),
    .in(arr__U501_in),
    .out(arr__U501_out)
);
assign arr__U508_clk = clk;
assign arr__U508_in[4] = arr__U501_out[4];
assign arr__U508_in[3] = arr__U501_out[3];
assign arr__U508_in[2] = arr__U501_out[2];
assign arr__U508_in[1] = arr__U501_out[1];
assign arr__U508_in[0] = arr__U501_out[0];
array_delay_U509 arr__U508 (
    .clk(arr__U508_clk),
    .in(arr__U508_in),
    .out(arr__U508_out)
);
assign arr__U515_clk = clk;
assign arr__U515_in[4] = arr__U508_out[4];
assign arr__U515_in[3] = arr__U508_out[3];
assign arr__U515_in[2] = arr__U508_out[2];
assign arr__U515_in[1] = arr__U508_out[1];
assign arr__U515_in[0] = arr__U508_out[0];
array_delay_U516 arr__U515 (
    .clk(arr__U515_clk),
    .in(arr__U515_in),
    .out(arr__U515_out)
);
assign arr__U522_clk = clk;
assign arr__U522_in[4] = arr__U515_out[4];
assign arr__U522_in[3] = arr__U515_out[3];
assign arr__U522_in[2] = arr__U515_out[2];
assign arr__U522_in[1] = arr__U515_out[1];
assign arr__U522_in[0] = arr__U515_out[0];
array_delay_U523 arr__U522 (
    .clk(arr__U522_clk),
    .in(arr__U522_in),
    .out(arr__U522_out)
);
assign arr__U529_clk = clk;
assign arr__U529_in[4] = arr__U522_out[4];
assign arr__U529_in[3] = arr__U522_out[3];
assign arr__U529_in[2] = arr__U522_out[2];
assign arr__U529_in[1] = arr__U522_out[1];
assign arr__U529_in[0] = arr__U522_out[0];
array_delay_U530 arr__U529 (
    .clk(arr__U529_clk),
    .in(arr__U529_in),
    .out(arr__U529_out)
);
assign arr__U536_clk = clk;
assign arr__U536_in[4] = arr__U529_out[4];
assign arr__U536_in[3] = arr__U529_out[3];
assign arr__U536_in[2] = arr__U529_out[2];
assign arr__U536_in[1] = arr__U529_out[1];
assign arr__U536_in[0] = arr__U529_out[0];
array_delay_U537 arr__U536 (
    .clk(arr__U536_clk),
    .in(arr__U536_in),
    .out(arr__U536_out)
);
assign arr__U543_clk = clk;
assign arr__U543_in[4] = arr__U536_out[4];
assign arr__U543_in[3] = arr__U536_out[3];
assign arr__U543_in[2] = arr__U536_out[2];
assign arr__U543_in[1] = arr__U536_out[1];
assign arr__U543_in[0] = arr__U536_out[0];
array_delay_U544 arr__U543 (
    .clk(arr__U543_clk),
    .in(arr__U543_in),
    .out(arr__U543_out)
);
assign arr__U550_clk = clk;
assign arr__U550_in[4] = arr__U543_out[4];
assign arr__U550_in[3] = arr__U543_out[3];
assign arr__U550_in[2] = arr__U543_out[2];
assign arr__U550_in[1] = arr__U543_out[1];
assign arr__U550_in[0] = arr__U543_out[0];
array_delay_U551 arr__U550 (
    .clk(arr__U550_clk),
    .in(arr__U550_in),
    .out(arr__U550_out)
);
assign arr__U557_clk = clk;
assign arr__U557_in[4] = arr__U550_out[4];
assign arr__U557_in[3] = arr__U550_out[3];
assign arr__U557_in[2] = arr__U550_out[2];
assign arr__U557_in[1] = arr__U550_out[1];
assign arr__U557_in[0] = arr__U550_out[0];
array_delay_U558 arr__U557 (
    .clk(arr__U557_clk),
    .in(arr__U557_in),
    .out(arr__U557_out)
);
assign arr__U564_clk = clk;
assign arr__U564_in[4] = arr__U557_out[4];
assign arr__U564_in[3] = arr__U557_out[3];
assign arr__U564_in[2] = arr__U557_out[2];
assign arr__U564_in[1] = arr__U557_out[1];
assign arr__U564_in[0] = arr__U557_out[0];
array_delay_U565 arr__U564 (
    .clk(arr__U564_clk),
    .in(arr__U564_in),
    .out(arr__U564_out)
);
assign arr__U571_clk = clk;
assign arr__U571_in[4] = arr__U564_out[4];
assign arr__U571_in[3] = arr__U564_out[3];
assign arr__U571_in[2] = arr__U564_out[2];
assign arr__U571_in[1] = arr__U564_out[1];
assign arr__U571_in[0] = arr__U564_out[0];
array_delay_U572 arr__U571 (
    .clk(arr__U571_clk),
    .in(arr__U571_in),
    .out(arr__U571_out)
);
assign arr__U578_clk = clk;
assign arr__U578_in[4] = arr__U571_out[4];
assign arr__U578_in[3] = arr__U571_out[3];
assign arr__U578_in[2] = arr__U571_out[2];
assign arr__U578_in[1] = arr__U571_out[1];
assign arr__U578_in[0] = arr__U571_out[0];
array_delay_U579 arr__U578 (
    .clk(arr__U578_clk),
    .in(arr__U578_in),
    .out(arr__U578_out)
);
assign arr__U585_clk = clk;
assign arr__U585_in[4] = arr__U578_out[4];
assign arr__U585_in[3] = arr__U578_out[3];
assign arr__U585_in[2] = arr__U578_out[2];
assign arr__U585_in[1] = arr__U578_out[1];
assign arr__U585_in[0] = arr__U578_out[0];
array_delay_U586 arr__U585 (
    .clk(arr__U585_clk),
    .in(arr__U585_in),
    .out(arr__U585_out)
);
assign arr__U628_clk = clk;
assign arr__U628_in[4] = op_hcompute_conv_stencil_9_port_controller_d[4];
assign arr__U628_in[3] = op_hcompute_conv_stencil_9_port_controller_d[3];
assign arr__U628_in[2] = op_hcompute_conv_stencil_9_port_controller_d[2];
assign arr__U628_in[1] = op_hcompute_conv_stencil_9_port_controller_d[1];
assign arr__U628_in[0] = op_hcompute_conv_stencil_9_port_controller_d[0];
array_delay_U629 arr__U628 (
    .clk(arr__U628_clk),
    .in(arr__U628_in),
    .out(arr__U628_out)
);
assign arr__U635_clk = clk;
assign arr__U635_in[4] = arr__U628_out[4];
assign arr__U635_in[3] = arr__U628_out[3];
assign arr__U635_in[2] = arr__U628_out[2];
assign arr__U635_in[1] = arr__U628_out[1];
assign arr__U635_in[0] = arr__U628_out[0];
array_delay_U636 arr__U635 (
    .clk(arr__U635_clk),
    .in(arr__U635_in),
    .out(arr__U635_out)
);
assign arr__U661_clk = clk;
assign arr__U661_in[4] = op_hcompute_conv_stencil_9_port_controller_d[4];
assign arr__U661_in[3] = op_hcompute_conv_stencil_9_port_controller_d[3];
assign arr__U661_in[2] = op_hcompute_conv_stencil_9_port_controller_d[2];
assign arr__U661_in[1] = op_hcompute_conv_stencil_9_port_controller_d[1];
assign arr__U661_in[0] = op_hcompute_conv_stencil_9_port_controller_d[0];
array_delay_U662 arr__U661 (
    .clk(arr__U661_clk),
    .in(arr__U661_in),
    .out(arr__U661_out)
);
assign arr__U668_clk = clk;
assign arr__U668_in[4] = arr__U661_out[4];
assign arr__U668_in[3] = arr__U661_out[3];
assign arr__U668_in[2] = arr__U661_out[2];
assign arr__U668_in[1] = arr__U661_out[1];
assign arr__U668_in[0] = arr__U661_out[0];
array_delay_U669 arr__U668 (
    .clk(arr__U668_clk),
    .in(arr__U668_in),
    .out(arr__U668_out)
);
assign arr__U675_clk = clk;
assign arr__U675_in[4] = arr__U668_out[4];
assign arr__U675_in[3] = arr__U668_out[3];
assign arr__U675_in[2] = arr__U668_out[2];
assign arr__U675_in[1] = arr__U668_out[1];
assign arr__U675_in[0] = arr__U668_out[0];
array_delay_U676 arr__U675 (
    .clk(arr__U675_clk),
    .in(arr__U675_in),
    .out(arr__U675_out)
);
assign arr__U682_clk = clk;
assign arr__U682_in[4] = arr__U675_out[4];
assign arr__U682_in[3] = arr__U675_out[3];
assign arr__U682_in[2] = arr__U675_out[2];
assign arr__U682_in[1] = arr__U675_out[1];
assign arr__U682_in[0] = arr__U675_out[0];
array_delay_U683 arr__U682 (
    .clk(arr__U682_clk),
    .in(arr__U682_in),
    .out(arr__U682_out)
);
assign arr__U689_clk = clk;
assign arr__U689_in[4] = arr__U682_out[4];
assign arr__U689_in[3] = arr__U682_out[3];
assign arr__U689_in[2] = arr__U682_out[2];
assign arr__U689_in[1] = arr__U682_out[1];
assign arr__U689_in[0] = arr__U682_out[0];
array_delay_U690 arr__U689 (
    .clk(arr__U689_clk),
    .in(arr__U689_in),
    .out(arr__U689_out)
);
assign arr__U696_clk = clk;
assign arr__U696_in[4] = arr__U689_out[4];
assign arr__U696_in[3] = arr__U689_out[3];
assign arr__U696_in[2] = arr__U689_out[2];
assign arr__U696_in[1] = arr__U689_out[1];
assign arr__U696_in[0] = arr__U689_out[0];
array_delay_U697 arr__U696 (
    .clk(arr__U696_clk),
    .in(arr__U696_in),
    .out(arr__U696_out)
);
assign arr__U703_clk = clk;
assign arr__U703_in[4] = arr__U696_out[4];
assign arr__U703_in[3] = arr__U696_out[3];
assign arr__U703_in[2] = arr__U696_out[2];
assign arr__U703_in[1] = arr__U696_out[1];
assign arr__U703_in[0] = arr__U696_out[0];
array_delay_U704 arr__U703 (
    .clk(arr__U703_clk),
    .in(arr__U703_in),
    .out(arr__U703_out)
);
assign arr__U710_clk = clk;
assign arr__U710_in[4] = arr__U703_out[4];
assign arr__U710_in[3] = arr__U703_out[3];
assign arr__U710_in[2] = arr__U703_out[2];
assign arr__U710_in[1] = arr__U703_out[1];
assign arr__U710_in[0] = arr__U703_out[0];
array_delay_U711 arr__U710 (
    .clk(arr__U710_clk),
    .in(arr__U710_in),
    .out(arr__U710_out)
);
assign arr__U717_clk = clk;
assign arr__U717_in[4] = arr__U710_out[4];
assign arr__U717_in[3] = arr__U710_out[3];
assign arr__U717_in[2] = arr__U710_out[2];
assign arr__U717_in[1] = arr__U710_out[1];
assign arr__U717_in[0] = arr__U710_out[0];
array_delay_U718 arr__U717 (
    .clk(arr__U717_clk),
    .in(arr__U717_in),
    .out(arr__U717_out)
);
assign arr__U724_clk = clk;
assign arr__U724_in[4] = arr__U717_out[4];
assign arr__U724_in[3] = arr__U717_out[3];
assign arr__U724_in[2] = arr__U717_out[2];
assign arr__U724_in[1] = arr__U717_out[1];
assign arr__U724_in[0] = arr__U717_out[0];
array_delay_U725 arr__U724 (
    .clk(arr__U724_clk),
    .in(arr__U724_in),
    .out(arr__U724_out)
);
assign arr__U731_clk = clk;
assign arr__U731_in[4] = arr__U724_out[4];
assign arr__U731_in[3] = arr__U724_out[3];
assign arr__U731_in[2] = arr__U724_out[2];
assign arr__U731_in[1] = arr__U724_out[1];
assign arr__U731_in[0] = arr__U724_out[0];
array_delay_U732 arr__U731 (
    .clk(arr__U731_clk),
    .in(arr__U731_in),
    .out(arr__U731_out)
);
assign arr__U738_clk = clk;
assign arr__U738_in[4] = arr__U731_out[4];
assign arr__U738_in[3] = arr__U731_out[3];
assign arr__U738_in[2] = arr__U731_out[2];
assign arr__U738_in[1] = arr__U731_out[1];
assign arr__U738_in[0] = arr__U731_out[0];
array_delay_U739 arr__U738 (
    .clk(arr__U738_clk),
    .in(arr__U738_in),
    .out(arr__U738_out)
);
assign arr__U745_clk = clk;
assign arr__U745_in[4] = arr__U738_out[4];
assign arr__U745_in[3] = arr__U738_out[3];
assign arr__U745_in[2] = arr__U738_out[2];
assign arr__U745_in[1] = arr__U738_out[1];
assign arr__U745_in[0] = arr__U738_out[0];
array_delay_U746 arr__U745 (
    .clk(arr__U745_clk),
    .in(arr__U745_in),
    .out(arr__U745_out)
);
assign arr__U752_clk = clk;
assign arr__U752_in[4] = arr__U745_out[4];
assign arr__U752_in[3] = arr__U745_out[3];
assign arr__U752_in[2] = arr__U745_out[2];
assign arr__U752_in[1] = arr__U745_out[1];
assign arr__U752_in[0] = arr__U745_out[0];
array_delay_U753 arr__U752 (
    .clk(arr__U752_clk),
    .in(arr__U752_in),
    .out(arr__U752_out)
);
assign arr__U759_clk = clk;
assign arr__U759_in[4] = arr__U752_out[4];
assign arr__U759_in[3] = arr__U752_out[3];
assign arr__U759_in[2] = arr__U752_out[2];
assign arr__U759_in[1] = arr__U752_out[1];
assign arr__U759_in[0] = arr__U752_out[0];
array_delay_U760 arr__U759 (
    .clk(arr__U759_clk),
    .in(arr__U759_in),
    .out(arr__U759_out)
);
assign arr__U766_clk = clk;
assign arr__U766_in[4] = arr__U759_out[4];
assign arr__U766_in[3] = arr__U759_out[3];
assign arr__U766_in[2] = arr__U759_out[2];
assign arr__U766_in[1] = arr__U759_out[1];
assign arr__U766_in[0] = arr__U759_out[0];
array_delay_U767 arr__U766 (
    .clk(arr__U766_clk),
    .in(arr__U766_in),
    .out(arr__U766_out)
);
assign arr__U773_clk = clk;
assign arr__U773_in[4] = arr__U766_out[4];
assign arr__U773_in[3] = arr__U766_out[3];
assign arr__U773_in[2] = arr__U766_out[2];
assign arr__U773_in[1] = arr__U766_out[1];
assign arr__U773_in[0] = arr__U766_out[0];
array_delay_U774 arr__U773 (
    .clk(arr__U773_clk),
    .in(arr__U773_in),
    .out(arr__U773_out)
);
assign arr__U816_clk = clk;
assign arr__U816_in[4] = op_hcompute_conv_stencil_10_port_controller_d[4];
assign arr__U816_in[3] = op_hcompute_conv_stencil_10_port_controller_d[3];
assign arr__U816_in[2] = op_hcompute_conv_stencil_10_port_controller_d[2];
assign arr__U816_in[1] = op_hcompute_conv_stencil_10_port_controller_d[1];
assign arr__U816_in[0] = op_hcompute_conv_stencil_10_port_controller_d[0];
array_delay_U817 arr__U816 (
    .clk(arr__U816_clk),
    .in(arr__U816_in),
    .out(arr__U816_out)
);
assign arr__U823_clk = clk;
assign arr__U823_in[4] = arr__U816_out[4];
assign arr__U823_in[3] = arr__U816_out[3];
assign arr__U823_in[2] = arr__U816_out[2];
assign arr__U823_in[1] = arr__U816_out[1];
assign arr__U823_in[0] = arr__U816_out[0];
array_delay_U824 arr__U823 (
    .clk(arr__U823_clk),
    .in(arr__U823_in),
    .out(arr__U823_out)
);
assign arr__U849_clk = clk;
assign arr__U849_in[4] = op_hcompute_conv_stencil_10_port_controller_d[4];
assign arr__U849_in[3] = op_hcompute_conv_stencil_10_port_controller_d[3];
assign arr__U849_in[2] = op_hcompute_conv_stencil_10_port_controller_d[2];
assign arr__U849_in[1] = op_hcompute_conv_stencil_10_port_controller_d[1];
assign arr__U849_in[0] = op_hcompute_conv_stencil_10_port_controller_d[0];
array_delay_U850 arr__U849 (
    .clk(arr__U849_clk),
    .in(arr__U849_in),
    .out(arr__U849_out)
);
assign arr__U856_clk = clk;
assign arr__U856_in[4] = arr__U849_out[4];
assign arr__U856_in[3] = arr__U849_out[3];
assign arr__U856_in[2] = arr__U849_out[2];
assign arr__U856_in[1] = arr__U849_out[1];
assign arr__U856_in[0] = arr__U849_out[0];
array_delay_U857 arr__U856 (
    .clk(arr__U856_clk),
    .in(arr__U856_in),
    .out(arr__U856_out)
);
assign arr__U863_clk = clk;
assign arr__U863_in[4] = arr__U856_out[4];
assign arr__U863_in[3] = arr__U856_out[3];
assign arr__U863_in[2] = arr__U856_out[2];
assign arr__U863_in[1] = arr__U856_out[1];
assign arr__U863_in[0] = arr__U856_out[0];
array_delay_U864 arr__U863 (
    .clk(arr__U863_clk),
    .in(arr__U863_in),
    .out(arr__U863_out)
);
assign arr__U870_clk = clk;
assign arr__U870_in[4] = arr__U863_out[4];
assign arr__U870_in[3] = arr__U863_out[3];
assign arr__U870_in[2] = arr__U863_out[2];
assign arr__U870_in[1] = arr__U863_out[1];
assign arr__U870_in[0] = arr__U863_out[0];
array_delay_U871 arr__U870 (
    .clk(arr__U870_clk),
    .in(arr__U870_in),
    .out(arr__U870_out)
);
assign arr__U877_clk = clk;
assign arr__U877_in[4] = arr__U870_out[4];
assign arr__U877_in[3] = arr__U870_out[3];
assign arr__U877_in[2] = arr__U870_out[2];
assign arr__U877_in[1] = arr__U870_out[1];
assign arr__U877_in[0] = arr__U870_out[0];
array_delay_U878 arr__U877 (
    .clk(arr__U877_clk),
    .in(arr__U877_in),
    .out(arr__U877_out)
);
assign arr__U884_clk = clk;
assign arr__U884_in[4] = arr__U877_out[4];
assign arr__U884_in[3] = arr__U877_out[3];
assign arr__U884_in[2] = arr__U877_out[2];
assign arr__U884_in[1] = arr__U877_out[1];
assign arr__U884_in[0] = arr__U877_out[0];
array_delay_U885 arr__U884 (
    .clk(arr__U884_clk),
    .in(arr__U884_in),
    .out(arr__U884_out)
);
assign arr__U891_clk = clk;
assign arr__U891_in[4] = arr__U884_out[4];
assign arr__U891_in[3] = arr__U884_out[3];
assign arr__U891_in[2] = arr__U884_out[2];
assign arr__U891_in[1] = arr__U884_out[1];
assign arr__U891_in[0] = arr__U884_out[0];
array_delay_U892 arr__U891 (
    .clk(arr__U891_clk),
    .in(arr__U891_in),
    .out(arr__U891_out)
);
assign arr__U898_clk = clk;
assign arr__U898_in[4] = arr__U891_out[4];
assign arr__U898_in[3] = arr__U891_out[3];
assign arr__U898_in[2] = arr__U891_out[2];
assign arr__U898_in[1] = arr__U891_out[1];
assign arr__U898_in[0] = arr__U891_out[0];
array_delay_U899 arr__U898 (
    .clk(arr__U898_clk),
    .in(arr__U898_in),
    .out(arr__U898_out)
);
assign arr__U905_clk = clk;
assign arr__U905_in[4] = arr__U898_out[4];
assign arr__U905_in[3] = arr__U898_out[3];
assign arr__U905_in[2] = arr__U898_out[2];
assign arr__U905_in[1] = arr__U898_out[1];
assign arr__U905_in[0] = arr__U898_out[0];
array_delay_U906 arr__U905 (
    .clk(arr__U905_clk),
    .in(arr__U905_in),
    .out(arr__U905_out)
);
assign arr__U912_clk = clk;
assign arr__U912_in[4] = arr__U905_out[4];
assign arr__U912_in[3] = arr__U905_out[3];
assign arr__U912_in[2] = arr__U905_out[2];
assign arr__U912_in[1] = arr__U905_out[1];
assign arr__U912_in[0] = arr__U905_out[0];
array_delay_U913 arr__U912 (
    .clk(arr__U912_clk),
    .in(arr__U912_in),
    .out(arr__U912_out)
);
assign arr__U919_clk = clk;
assign arr__U919_in[4] = arr__U912_out[4];
assign arr__U919_in[3] = arr__U912_out[3];
assign arr__U919_in[2] = arr__U912_out[2];
assign arr__U919_in[1] = arr__U912_out[1];
assign arr__U919_in[0] = arr__U912_out[0];
array_delay_U920 arr__U919 (
    .clk(arr__U919_clk),
    .in(arr__U919_in),
    .out(arr__U919_out)
);
assign arr__U926_clk = clk;
assign arr__U926_in[4] = arr__U919_out[4];
assign arr__U926_in[3] = arr__U919_out[3];
assign arr__U926_in[2] = arr__U919_out[2];
assign arr__U926_in[1] = arr__U919_out[1];
assign arr__U926_in[0] = arr__U919_out[0];
array_delay_U927 arr__U926 (
    .clk(arr__U926_clk),
    .in(arr__U926_in),
    .out(arr__U926_out)
);
assign arr__U933_clk = clk;
assign arr__U933_in[4] = arr__U926_out[4];
assign arr__U933_in[3] = arr__U926_out[3];
assign arr__U933_in[2] = arr__U926_out[2];
assign arr__U933_in[1] = arr__U926_out[1];
assign arr__U933_in[0] = arr__U926_out[0];
array_delay_U934 arr__U933 (
    .clk(arr__U933_clk),
    .in(arr__U933_in),
    .out(arr__U933_out)
);
assign arr__U940_clk = clk;
assign arr__U940_in[4] = arr__U933_out[4];
assign arr__U940_in[3] = arr__U933_out[3];
assign arr__U940_in[2] = arr__U933_out[2];
assign arr__U940_in[1] = arr__U933_out[1];
assign arr__U940_in[0] = arr__U933_out[0];
array_delay_U941 arr__U940 (
    .clk(arr__U940_clk),
    .in(arr__U940_in),
    .out(arr__U940_out)
);
assign arr__U947_clk = clk;
assign arr__U947_in[4] = arr__U940_out[4];
assign arr__U947_in[3] = arr__U940_out[3];
assign arr__U947_in[2] = arr__U940_out[2];
assign arr__U947_in[1] = arr__U940_out[1];
assign arr__U947_in[0] = arr__U940_out[0];
array_delay_U948 arr__U947 (
    .clk(arr__U947_clk),
    .in(arr__U947_in),
    .out(arr__U947_out)
);
assign arr__U954_clk = clk;
assign arr__U954_in[4] = arr__U947_out[4];
assign arr__U954_in[3] = arr__U947_out[3];
assign arr__U954_in[2] = arr__U947_out[2];
assign arr__U954_in[1] = arr__U947_out[1];
assign arr__U954_in[0] = arr__U947_out[0];
array_delay_U955 arr__U954 (
    .clk(arr__U954_clk),
    .in(arr__U954_in),
    .out(arr__U954_out)
);
assign arr__U961_clk = clk;
assign arr__U961_in[4] = arr__U954_out[4];
assign arr__U961_in[3] = arr__U954_out[3];
assign arr__U961_in[2] = arr__U954_out[2];
assign arr__U961_in[1] = arr__U954_out[1];
assign arr__U961_in[0] = arr__U954_out[0];
array_delay_U962 arr__U961 (
    .clk(arr__U961_clk),
    .in(arr__U961_in),
    .out(arr__U961_out)
);
assign conv_stencil_clk = clk;
assign conv_stencil_flush = flush;
assign conv_stencil_rst_n = rst_n;
assign conv_stencil_op_hcompute_conv_stencil_10_read_ren = op_hcompute_conv_stencil_10_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[4] = op_hcompute_conv_stencil_10_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[3] = op_hcompute_conv_stencil_10_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[2] = op_hcompute_conv_stencil_10_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[1] = op_hcompute_conv_stencil_10_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[0] = op_hcompute_conv_stencil_10_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_10_write_wen = op_hcompute_conv_stencil_10_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_10_write_ctrl_vars[4] = op_hcompute_conv_stencil_10_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_10_write_ctrl_vars[3] = op_hcompute_conv_stencil_10_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_10_write_ctrl_vars[2] = op_hcompute_conv_stencil_10_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_10_write_ctrl_vars[1] = op_hcompute_conv_stencil_10_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_10_write_ctrl_vars[0] = op_hcompute_conv_stencil_10_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_10_write[0] = op_hcompute_conv_stencil_10_conv_stencil_op_hcompute_conv_stencil_10_write[0];
assign conv_stencil_op_hcompute_conv_stencil_11_read_ren = op_hcompute_conv_stencil_11_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[4] = op_hcompute_conv_stencil_11_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[3] = op_hcompute_conv_stencil_11_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[2] = op_hcompute_conv_stencil_11_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[1] = op_hcompute_conv_stencil_11_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[0] = op_hcompute_conv_stencil_11_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_11_write_wen = op_hcompute_conv_stencil_11_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_11_write_ctrl_vars[4] = op_hcompute_conv_stencil_11_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_11_write_ctrl_vars[3] = op_hcompute_conv_stencil_11_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_11_write_ctrl_vars[2] = op_hcompute_conv_stencil_11_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_11_write_ctrl_vars[1] = op_hcompute_conv_stencil_11_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_11_write_ctrl_vars[0] = op_hcompute_conv_stencil_11_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_11_write[0] = op_hcompute_conv_stencil_11_conv_stencil_op_hcompute_conv_stencil_11_write[0];
assign conv_stencil_op_hcompute_conv_stencil_12_read_ren = op_hcompute_conv_stencil_12_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[4] = op_hcompute_conv_stencil_12_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[3] = op_hcompute_conv_stencil_12_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[2] = op_hcompute_conv_stencil_12_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[1] = op_hcompute_conv_stencil_12_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[0] = op_hcompute_conv_stencil_12_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_12_write_wen = op_hcompute_conv_stencil_12_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_12_write_ctrl_vars[4] = op_hcompute_conv_stencil_12_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_12_write_ctrl_vars[3] = op_hcompute_conv_stencil_12_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_12_write_ctrl_vars[2] = op_hcompute_conv_stencil_12_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_12_write_ctrl_vars[1] = op_hcompute_conv_stencil_12_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_12_write_ctrl_vars[0] = op_hcompute_conv_stencil_12_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_12_write[0] = op_hcompute_conv_stencil_12_conv_stencil_op_hcompute_conv_stencil_12_write[0];
assign conv_stencil_op_hcompute_conv_stencil_13_read_ren = op_hcompute_conv_stencil_13_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[4] = op_hcompute_conv_stencil_13_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[3] = op_hcompute_conv_stencil_13_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[2] = op_hcompute_conv_stencil_13_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[1] = op_hcompute_conv_stencil_13_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[0] = op_hcompute_conv_stencil_13_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_13_write_wen = op_hcompute_conv_stencil_13_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_13_write_ctrl_vars[4] = op_hcompute_conv_stencil_13_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_13_write_ctrl_vars[3] = op_hcompute_conv_stencil_13_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_13_write_ctrl_vars[2] = op_hcompute_conv_stencil_13_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_13_write_ctrl_vars[1] = op_hcompute_conv_stencil_13_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_13_write_ctrl_vars[0] = op_hcompute_conv_stencil_13_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_13_write[0] = op_hcompute_conv_stencil_13_conv_stencil_op_hcompute_conv_stencil_13_write[0];
assign conv_stencil_op_hcompute_conv_stencil_14_read_ren = op_hcompute_conv_stencil_14_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[4] = op_hcompute_conv_stencil_14_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[3] = op_hcompute_conv_stencil_14_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[2] = op_hcompute_conv_stencil_14_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[1] = op_hcompute_conv_stencil_14_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[0] = op_hcompute_conv_stencil_14_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_14_write_wen = op_hcompute_conv_stencil_14_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_14_write_ctrl_vars[4] = op_hcompute_conv_stencil_14_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_14_write_ctrl_vars[3] = op_hcompute_conv_stencil_14_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_14_write_ctrl_vars[2] = op_hcompute_conv_stencil_14_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_14_write_ctrl_vars[1] = op_hcompute_conv_stencil_14_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_14_write_ctrl_vars[0] = op_hcompute_conv_stencil_14_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_14_write[0] = op_hcompute_conv_stencil_14_conv_stencil_op_hcompute_conv_stencil_14_write[0];
assign conv_stencil_op_hcompute_conv_stencil_15_read_ren = op_hcompute_conv_stencil_15_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[4] = op_hcompute_conv_stencil_15_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[3] = op_hcompute_conv_stencil_15_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[2] = op_hcompute_conv_stencil_15_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[1] = op_hcompute_conv_stencil_15_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[0] = op_hcompute_conv_stencil_15_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_15_write_wen = op_hcompute_conv_stencil_15_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_15_write_ctrl_vars[4] = op_hcompute_conv_stencil_15_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_15_write_ctrl_vars[3] = op_hcompute_conv_stencil_15_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_15_write_ctrl_vars[2] = op_hcompute_conv_stencil_15_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_15_write_ctrl_vars[1] = op_hcompute_conv_stencil_15_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_15_write_ctrl_vars[0] = op_hcompute_conv_stencil_15_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_15_write[0] = op_hcompute_conv_stencil_15_conv_stencil_op_hcompute_conv_stencil_15_write[0];
assign conv_stencil_op_hcompute_conv_stencil_1_write_wen = op_hcompute_conv_stencil_1_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[2] = op_hcompute_conv_stencil_1_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[1] = op_hcompute_conv_stencil_1_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[0] = op_hcompute_conv_stencil_1_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write[0];
assign conv_stencil_op_hcompute_conv_stencil_2_write_wen = op_hcompute_conv_stencil_2_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[2] = op_hcompute_conv_stencil_2_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[1] = op_hcompute_conv_stencil_2_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[0] = op_hcompute_conv_stencil_2_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write[0];
assign conv_stencil_op_hcompute_conv_stencil_3_write_wen = op_hcompute_conv_stencil_3_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[2] = op_hcompute_conv_stencil_3_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[1] = op_hcompute_conv_stencil_3_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[0] = op_hcompute_conv_stencil_3_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write[0];
assign conv_stencil_op_hcompute_conv_stencil_4_write_wen = op_hcompute_conv_stencil_4_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[2] = op_hcompute_conv_stencil_4_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[1] = op_hcompute_conv_stencil_4_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[0] = op_hcompute_conv_stencil_4_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write[0];
assign conv_stencil_op_hcompute_conv_stencil_5_write_wen = op_hcompute_conv_stencil_5_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[2] = op_hcompute_conv_stencil_5_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[1] = op_hcompute_conv_stencil_5_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[0] = op_hcompute_conv_stencil_5_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write[0];
assign conv_stencil_op_hcompute_conv_stencil_6_write_wen = op_hcompute_conv_stencil_6_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_6_write_ctrl_vars[2] = op_hcompute_conv_stencil_6_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_6_write_ctrl_vars[1] = op_hcompute_conv_stencil_6_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_6_write_ctrl_vars[0] = op_hcompute_conv_stencil_6_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_6_write[0] = op_hcompute_conv_stencil_6_conv_stencil_op_hcompute_conv_stencil_6_write[0];
assign conv_stencil_op_hcompute_conv_stencil_7_write_wen = op_hcompute_conv_stencil_7_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_7_write_ctrl_vars[2] = op_hcompute_conv_stencil_7_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_7_write_ctrl_vars[1] = op_hcompute_conv_stencil_7_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_7_write_ctrl_vars[0] = op_hcompute_conv_stencil_7_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_7_write[0] = op_hcompute_conv_stencil_7_conv_stencil_op_hcompute_conv_stencil_7_write[0];
assign conv_stencil_op_hcompute_conv_stencil_8_read_ren = op_hcompute_conv_stencil_8_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[4] = op_hcompute_conv_stencil_8_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[3] = op_hcompute_conv_stencil_8_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[2] = op_hcompute_conv_stencil_8_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[1] = op_hcompute_conv_stencil_8_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[0] = op_hcompute_conv_stencil_8_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_8_write_wen = op_hcompute_conv_stencil_8_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_8_write_ctrl_vars[4] = op_hcompute_conv_stencil_8_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_8_write_ctrl_vars[3] = op_hcompute_conv_stencil_8_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_8_write_ctrl_vars[2] = op_hcompute_conv_stencil_8_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_8_write_ctrl_vars[1] = op_hcompute_conv_stencil_8_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_8_write_ctrl_vars[0] = op_hcompute_conv_stencil_8_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_8_write[0] = op_hcompute_conv_stencil_8_conv_stencil_op_hcompute_conv_stencil_8_write[0];
assign conv_stencil_op_hcompute_conv_stencil_9_read_ren = op_hcompute_conv_stencil_9_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[4] = op_hcompute_conv_stencil_9_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[3] = op_hcompute_conv_stencil_9_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[2] = op_hcompute_conv_stencil_9_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[1] = op_hcompute_conv_stencil_9_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[0] = op_hcompute_conv_stencil_9_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_9_write_wen = op_hcompute_conv_stencil_9_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_9_write_ctrl_vars[4] = op_hcompute_conv_stencil_9_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_9_write_ctrl_vars[3] = op_hcompute_conv_stencil_9_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_9_write_ctrl_vars[2] = op_hcompute_conv_stencil_9_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_9_write_ctrl_vars[1] = op_hcompute_conv_stencil_9_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_9_write_ctrl_vars[0] = op_hcompute_conv_stencil_9_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_9_write[0] = op_hcompute_conv_stencil_9_conv_stencil_op_hcompute_conv_stencil_9_write[0];
assign conv_stencil_op_hcompute_conv_stencil_write_wen = op_hcompute_conv_stencil_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[2] = op_hcompute_conv_stencil_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[1] = op_hcompute_conv_stencil_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[0] = op_hcompute_conv_stencil_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_write[0] = op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write[0];
assign conv_stencil_op_hcompute_hw_output_stencil_1_read_ren = op_hcompute_hw_output_stencil_1_read_start_out;
assign conv_stencil_op_hcompute_hw_output_stencil_1_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_1_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_1_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_1_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_1_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_1_port_controller_d[0];
assign conv_stencil_op_hcompute_hw_output_stencil_2_read_ren = op_hcompute_hw_output_stencil_2_read_start_out;
assign conv_stencil_op_hcompute_hw_output_stencil_2_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_2_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_2_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_2_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_2_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_2_port_controller_d[0];
assign conv_stencil_op_hcompute_hw_output_stencil_3_read_ren = op_hcompute_hw_output_stencil_3_read_start_out;
assign conv_stencil_op_hcompute_hw_output_stencil_3_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_3_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_3_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_3_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_3_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_3_port_controller_d[0];
assign conv_stencil_op_hcompute_hw_output_stencil_4_read_ren = op_hcompute_hw_output_stencil_4_read_start_out;
assign conv_stencil_op_hcompute_hw_output_stencil_4_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_4_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_4_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_4_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_4_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_4_port_controller_d[0];
assign conv_stencil_op_hcompute_hw_output_stencil_5_read_ren = op_hcompute_hw_output_stencil_5_read_start_out;
assign conv_stencil_op_hcompute_hw_output_stencil_5_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_5_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_5_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_5_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_5_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_5_port_controller_d[0];
assign conv_stencil_op_hcompute_hw_output_stencil_6_read_ren = op_hcompute_hw_output_stencil_6_read_start_out;
assign conv_stencil_op_hcompute_hw_output_stencil_6_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_6_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_6_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_6_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_6_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_6_port_controller_d[0];
assign conv_stencil_op_hcompute_hw_output_stencil_7_read_ren = op_hcompute_hw_output_stencil_7_read_start_out;
assign conv_stencil_op_hcompute_hw_output_stencil_7_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_7_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_7_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_7_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_7_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_7_port_controller_d[0];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ren = op_hcompute_hw_output_stencil_read_start_out;
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
conv_stencil_ub conv_stencil (
    .clk(conv_stencil_clk),
    .flush(conv_stencil_flush),
    .rst_n(conv_stencil_rst_n),
    .op_hcompute_conv_stencil_10_read_ren(conv_stencil_op_hcompute_conv_stencil_10_read_ren),
    .op_hcompute_conv_stencil_10_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars),
    .op_hcompute_conv_stencil_10_read(conv_stencil_op_hcompute_conv_stencil_10_read),
    .op_hcompute_conv_stencil_10_write_wen(conv_stencil_op_hcompute_conv_stencil_10_write_wen),
    .op_hcompute_conv_stencil_10_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_10_write_ctrl_vars),
    .op_hcompute_conv_stencil_10_write(conv_stencil_op_hcompute_conv_stencil_10_write),
    .op_hcompute_conv_stencil_11_read_ren(conv_stencil_op_hcompute_conv_stencil_11_read_ren),
    .op_hcompute_conv_stencil_11_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars),
    .op_hcompute_conv_stencil_11_read(conv_stencil_op_hcompute_conv_stencil_11_read),
    .op_hcompute_conv_stencil_11_write_wen(conv_stencil_op_hcompute_conv_stencil_11_write_wen),
    .op_hcompute_conv_stencil_11_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_11_write_ctrl_vars),
    .op_hcompute_conv_stencil_11_write(conv_stencil_op_hcompute_conv_stencil_11_write),
    .op_hcompute_conv_stencil_12_read_ren(conv_stencil_op_hcompute_conv_stencil_12_read_ren),
    .op_hcompute_conv_stencil_12_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars),
    .op_hcompute_conv_stencil_12_read(conv_stencil_op_hcompute_conv_stencil_12_read),
    .op_hcompute_conv_stencil_12_write_wen(conv_stencil_op_hcompute_conv_stencil_12_write_wen),
    .op_hcompute_conv_stencil_12_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_12_write_ctrl_vars),
    .op_hcompute_conv_stencil_12_write(conv_stencil_op_hcompute_conv_stencil_12_write),
    .op_hcompute_conv_stencil_13_read_ren(conv_stencil_op_hcompute_conv_stencil_13_read_ren),
    .op_hcompute_conv_stencil_13_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars),
    .op_hcompute_conv_stencil_13_read(conv_stencil_op_hcompute_conv_stencil_13_read),
    .op_hcompute_conv_stencil_13_write_wen(conv_stencil_op_hcompute_conv_stencil_13_write_wen),
    .op_hcompute_conv_stencil_13_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_13_write_ctrl_vars),
    .op_hcompute_conv_stencil_13_write(conv_stencil_op_hcompute_conv_stencil_13_write),
    .op_hcompute_conv_stencil_14_read_ren(conv_stencil_op_hcompute_conv_stencil_14_read_ren),
    .op_hcompute_conv_stencil_14_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars),
    .op_hcompute_conv_stencil_14_read(conv_stencil_op_hcompute_conv_stencil_14_read),
    .op_hcompute_conv_stencil_14_write_wen(conv_stencil_op_hcompute_conv_stencil_14_write_wen),
    .op_hcompute_conv_stencil_14_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_14_write_ctrl_vars),
    .op_hcompute_conv_stencil_14_write(conv_stencil_op_hcompute_conv_stencil_14_write),
    .op_hcompute_conv_stencil_15_read_ren(conv_stencil_op_hcompute_conv_stencil_15_read_ren),
    .op_hcompute_conv_stencil_15_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars),
    .op_hcompute_conv_stencil_15_read(conv_stencil_op_hcompute_conv_stencil_15_read),
    .op_hcompute_conv_stencil_15_write_wen(conv_stencil_op_hcompute_conv_stencil_15_write_wen),
    .op_hcompute_conv_stencil_15_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_15_write_ctrl_vars),
    .op_hcompute_conv_stencil_15_write(conv_stencil_op_hcompute_conv_stencil_15_write),
    .op_hcompute_conv_stencil_1_write_wen(conv_stencil_op_hcompute_conv_stencil_1_write_wen),
    .op_hcompute_conv_stencil_1_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars),
    .op_hcompute_conv_stencil_1_write(conv_stencil_op_hcompute_conv_stencil_1_write),
    .op_hcompute_conv_stencil_2_write_wen(conv_stencil_op_hcompute_conv_stencil_2_write_wen),
    .op_hcompute_conv_stencil_2_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars),
    .op_hcompute_conv_stencil_2_write(conv_stencil_op_hcompute_conv_stencil_2_write),
    .op_hcompute_conv_stencil_3_write_wen(conv_stencil_op_hcompute_conv_stencil_3_write_wen),
    .op_hcompute_conv_stencil_3_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars),
    .op_hcompute_conv_stencil_3_write(conv_stencil_op_hcompute_conv_stencil_3_write),
    .op_hcompute_conv_stencil_4_write_wen(conv_stencil_op_hcompute_conv_stencil_4_write_wen),
    .op_hcompute_conv_stencil_4_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars),
    .op_hcompute_conv_stencil_4_write(conv_stencil_op_hcompute_conv_stencil_4_write),
    .op_hcompute_conv_stencil_5_write_wen(conv_stencil_op_hcompute_conv_stencil_5_write_wen),
    .op_hcompute_conv_stencil_5_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars),
    .op_hcompute_conv_stencil_5_write(conv_stencil_op_hcompute_conv_stencil_5_write),
    .op_hcompute_conv_stencil_6_write_wen(conv_stencil_op_hcompute_conv_stencil_6_write_wen),
    .op_hcompute_conv_stencil_6_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_6_write_ctrl_vars),
    .op_hcompute_conv_stencil_6_write(conv_stencil_op_hcompute_conv_stencil_6_write),
    .op_hcompute_conv_stencil_7_write_wen(conv_stencil_op_hcompute_conv_stencil_7_write_wen),
    .op_hcompute_conv_stencil_7_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_7_write_ctrl_vars),
    .op_hcompute_conv_stencil_7_write(conv_stencil_op_hcompute_conv_stencil_7_write),
    .op_hcompute_conv_stencil_8_read_ren(conv_stencil_op_hcompute_conv_stencil_8_read_ren),
    .op_hcompute_conv_stencil_8_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars),
    .op_hcompute_conv_stencil_8_read(conv_stencil_op_hcompute_conv_stencil_8_read),
    .op_hcompute_conv_stencil_8_write_wen(conv_stencil_op_hcompute_conv_stencil_8_write_wen),
    .op_hcompute_conv_stencil_8_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_8_write_ctrl_vars),
    .op_hcompute_conv_stencil_8_write(conv_stencil_op_hcompute_conv_stencil_8_write),
    .op_hcompute_conv_stencil_9_read_ren(conv_stencil_op_hcompute_conv_stencil_9_read_ren),
    .op_hcompute_conv_stencil_9_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars),
    .op_hcompute_conv_stencil_9_read(conv_stencil_op_hcompute_conv_stencil_9_read),
    .op_hcompute_conv_stencil_9_write_wen(conv_stencil_op_hcompute_conv_stencil_9_write_wen),
    .op_hcompute_conv_stencil_9_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_9_write_ctrl_vars),
    .op_hcompute_conv_stencil_9_write(conv_stencil_op_hcompute_conv_stencil_9_write),
    .op_hcompute_conv_stencil_write_wen(conv_stencil_op_hcompute_conv_stencil_write_wen),
    .op_hcompute_conv_stencil_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars),
    .op_hcompute_conv_stencil_write(conv_stencil_op_hcompute_conv_stencil_write),
    .op_hcompute_hw_output_stencil_1_read_ren(conv_stencil_op_hcompute_hw_output_stencil_1_read_ren),
    .op_hcompute_hw_output_stencil_1_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_1_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_1_read(conv_stencil_op_hcompute_hw_output_stencil_1_read),
    .op_hcompute_hw_output_stencil_2_read_ren(conv_stencil_op_hcompute_hw_output_stencil_2_read_ren),
    .op_hcompute_hw_output_stencil_2_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_2_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_2_read(conv_stencil_op_hcompute_hw_output_stencil_2_read),
    .op_hcompute_hw_output_stencil_3_read_ren(conv_stencil_op_hcompute_hw_output_stencil_3_read_ren),
    .op_hcompute_hw_output_stencil_3_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_3_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_3_read(conv_stencil_op_hcompute_hw_output_stencil_3_read),
    .op_hcompute_hw_output_stencil_4_read_ren(conv_stencil_op_hcompute_hw_output_stencil_4_read_ren),
    .op_hcompute_hw_output_stencil_4_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_4_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_4_read(conv_stencil_op_hcompute_hw_output_stencil_4_read),
    .op_hcompute_hw_output_stencil_5_read_ren(conv_stencil_op_hcompute_hw_output_stencil_5_read_ren),
    .op_hcompute_hw_output_stencil_5_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_5_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_5_read(conv_stencil_op_hcompute_hw_output_stencil_5_read),
    .op_hcompute_hw_output_stencil_6_read_ren(conv_stencil_op_hcompute_hw_output_stencil_6_read_ren),
    .op_hcompute_hw_output_stencil_6_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_6_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_6_read(conv_stencil_op_hcompute_hw_output_stencil_6_read),
    .op_hcompute_hw_output_stencil_7_read_ren(conv_stencil_op_hcompute_hw_output_stencil_7_read_ren),
    .op_hcompute_hw_output_stencil_7_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_7_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_7_read(conv_stencil_op_hcompute_hw_output_stencil_7_read),
    .op_hcompute_hw_output_stencil_read_ren(conv_stencil_op_hcompute_hw_output_stencil_read_ren),
    .op_hcompute_hw_output_stencil_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_read(conv_stencil_op_hcompute_hw_output_stencil_read)
);
assign delay_reg__U1001_clk = clk;
assign delay_reg__U1001_in = op_hcompute_conv_stencil_11_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1001 (
    .clk(delay_reg__U1001_clk),
    .in(delay_reg__U1001_in),
    .out(delay_reg__U1001_out)
);
assign delay_reg__U1002_clk = clk;
assign delay_reg__U1002_in = delay_reg__U1001_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1002 (
    .clk(delay_reg__U1002_clk),
    .in(delay_reg__U1002_in),
    .out(delay_reg__U1002_out)
);
assign delay_reg__U1019_clk = clk;
assign delay_reg__U1019_in = op_hcompute_conv_stencil_11_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1019 (
    .clk(delay_reg__U1019_clk),
    .in(delay_reg__U1019_in),
    .out(delay_reg__U1019_out)
);
assign delay_reg__U1020_clk = clk;
assign delay_reg__U1020_in = delay_reg__U1019_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1020 (
    .clk(delay_reg__U1020_clk),
    .in(delay_reg__U1020_in),
    .out(delay_reg__U1020_out)
);
assign delay_reg__U1021_clk = clk;
assign delay_reg__U1021_in = delay_reg__U1020_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1021 (
    .clk(delay_reg__U1021_clk),
    .in(delay_reg__U1021_in),
    .out(delay_reg__U1021_out)
);
assign delay_reg__U1022_clk = clk;
assign delay_reg__U1022_in = delay_reg__U1021_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1022 (
    .clk(delay_reg__U1022_clk),
    .in(delay_reg__U1022_in),
    .out(delay_reg__U1022_out)
);
assign delay_reg__U1023_clk = clk;
assign delay_reg__U1023_in = delay_reg__U1022_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1023 (
    .clk(delay_reg__U1023_clk),
    .in(delay_reg__U1023_in),
    .out(delay_reg__U1023_out)
);
assign delay_reg__U1024_clk = clk;
assign delay_reg__U1024_in = delay_reg__U1023_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1024 (
    .clk(delay_reg__U1024_clk),
    .in(delay_reg__U1024_in),
    .out(delay_reg__U1024_out)
);
assign delay_reg__U1025_clk = clk;
assign delay_reg__U1025_in = delay_reg__U1024_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1025 (
    .clk(delay_reg__U1025_clk),
    .in(delay_reg__U1025_in),
    .out(delay_reg__U1025_out)
);
assign delay_reg__U1026_clk = clk;
assign delay_reg__U1026_in = delay_reg__U1025_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1026 (
    .clk(delay_reg__U1026_clk),
    .in(delay_reg__U1026_in),
    .out(delay_reg__U1026_out)
);
assign delay_reg__U1027_clk = clk;
assign delay_reg__U1027_in = delay_reg__U1026_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1027 (
    .clk(delay_reg__U1027_clk),
    .in(delay_reg__U1027_in),
    .out(delay_reg__U1027_out)
);
assign delay_reg__U1028_clk = clk;
assign delay_reg__U1028_in = delay_reg__U1027_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1028 (
    .clk(delay_reg__U1028_clk),
    .in(delay_reg__U1028_in),
    .out(delay_reg__U1028_out)
);
assign delay_reg__U1029_clk = clk;
assign delay_reg__U1029_in = delay_reg__U1028_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1029 (
    .clk(delay_reg__U1029_clk),
    .in(delay_reg__U1029_in),
    .out(delay_reg__U1029_out)
);
assign delay_reg__U1030_clk = clk;
assign delay_reg__U1030_in = delay_reg__U1029_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1030 (
    .clk(delay_reg__U1030_clk),
    .in(delay_reg__U1030_in),
    .out(delay_reg__U1030_out)
);
assign delay_reg__U1031_clk = clk;
assign delay_reg__U1031_in = delay_reg__U1030_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1031 (
    .clk(delay_reg__U1031_clk),
    .in(delay_reg__U1031_in),
    .out(delay_reg__U1031_out)
);
assign delay_reg__U1032_clk = clk;
assign delay_reg__U1032_in = delay_reg__U1031_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1032 (
    .clk(delay_reg__U1032_clk),
    .in(delay_reg__U1032_in),
    .out(delay_reg__U1032_out)
);
assign delay_reg__U1033_clk = clk;
assign delay_reg__U1033_in = delay_reg__U1032_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1033 (
    .clk(delay_reg__U1033_clk),
    .in(delay_reg__U1033_in),
    .out(delay_reg__U1033_out)
);
assign delay_reg__U1034_clk = clk;
assign delay_reg__U1034_in = delay_reg__U1033_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1034 (
    .clk(delay_reg__U1034_clk),
    .in(delay_reg__U1034_in),
    .out(delay_reg__U1034_out)
);
assign delay_reg__U1035_clk = clk;
assign delay_reg__U1035_in = delay_reg__U1034_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1035 (
    .clk(delay_reg__U1035_clk),
    .in(delay_reg__U1035_in),
    .out(delay_reg__U1035_out)
);
assign delay_reg__U1189_clk = clk;
assign delay_reg__U1189_in = op_hcompute_conv_stencil_12_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1189 (
    .clk(delay_reg__U1189_clk),
    .in(delay_reg__U1189_in),
    .out(delay_reg__U1189_out)
);
assign delay_reg__U1190_clk = clk;
assign delay_reg__U1190_in = delay_reg__U1189_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1190 (
    .clk(delay_reg__U1190_clk),
    .in(delay_reg__U1190_in),
    .out(delay_reg__U1190_out)
);
assign delay_reg__U1207_clk = clk;
assign delay_reg__U1207_in = op_hcompute_conv_stencil_12_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1207 (
    .clk(delay_reg__U1207_clk),
    .in(delay_reg__U1207_in),
    .out(delay_reg__U1207_out)
);
assign delay_reg__U1208_clk = clk;
assign delay_reg__U1208_in = delay_reg__U1207_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1208 (
    .clk(delay_reg__U1208_clk),
    .in(delay_reg__U1208_in),
    .out(delay_reg__U1208_out)
);
assign delay_reg__U1209_clk = clk;
assign delay_reg__U1209_in = delay_reg__U1208_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1209 (
    .clk(delay_reg__U1209_clk),
    .in(delay_reg__U1209_in),
    .out(delay_reg__U1209_out)
);
assign delay_reg__U1210_clk = clk;
assign delay_reg__U1210_in = delay_reg__U1209_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1210 (
    .clk(delay_reg__U1210_clk),
    .in(delay_reg__U1210_in),
    .out(delay_reg__U1210_out)
);
assign delay_reg__U1211_clk = clk;
assign delay_reg__U1211_in = delay_reg__U1210_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1211 (
    .clk(delay_reg__U1211_clk),
    .in(delay_reg__U1211_in),
    .out(delay_reg__U1211_out)
);
assign delay_reg__U1212_clk = clk;
assign delay_reg__U1212_in = delay_reg__U1211_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1212 (
    .clk(delay_reg__U1212_clk),
    .in(delay_reg__U1212_in),
    .out(delay_reg__U1212_out)
);
assign delay_reg__U1213_clk = clk;
assign delay_reg__U1213_in = delay_reg__U1212_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1213 (
    .clk(delay_reg__U1213_clk),
    .in(delay_reg__U1213_in),
    .out(delay_reg__U1213_out)
);
assign delay_reg__U1214_clk = clk;
assign delay_reg__U1214_in = delay_reg__U1213_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1214 (
    .clk(delay_reg__U1214_clk),
    .in(delay_reg__U1214_in),
    .out(delay_reg__U1214_out)
);
assign delay_reg__U1215_clk = clk;
assign delay_reg__U1215_in = delay_reg__U1214_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1215 (
    .clk(delay_reg__U1215_clk),
    .in(delay_reg__U1215_in),
    .out(delay_reg__U1215_out)
);
assign delay_reg__U1216_clk = clk;
assign delay_reg__U1216_in = delay_reg__U1215_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1216 (
    .clk(delay_reg__U1216_clk),
    .in(delay_reg__U1216_in),
    .out(delay_reg__U1216_out)
);
assign delay_reg__U1217_clk = clk;
assign delay_reg__U1217_in = delay_reg__U1216_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1217 (
    .clk(delay_reg__U1217_clk),
    .in(delay_reg__U1217_in),
    .out(delay_reg__U1217_out)
);
assign delay_reg__U1218_clk = clk;
assign delay_reg__U1218_in = delay_reg__U1217_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1218 (
    .clk(delay_reg__U1218_clk),
    .in(delay_reg__U1218_in),
    .out(delay_reg__U1218_out)
);
assign delay_reg__U1219_clk = clk;
assign delay_reg__U1219_in = delay_reg__U1218_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1219 (
    .clk(delay_reg__U1219_clk),
    .in(delay_reg__U1219_in),
    .out(delay_reg__U1219_out)
);
assign delay_reg__U1220_clk = clk;
assign delay_reg__U1220_in = delay_reg__U1219_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1220 (
    .clk(delay_reg__U1220_clk),
    .in(delay_reg__U1220_in),
    .out(delay_reg__U1220_out)
);
assign delay_reg__U1221_clk = clk;
assign delay_reg__U1221_in = delay_reg__U1220_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1221 (
    .clk(delay_reg__U1221_clk),
    .in(delay_reg__U1221_in),
    .out(delay_reg__U1221_out)
);
assign delay_reg__U1222_clk = clk;
assign delay_reg__U1222_in = delay_reg__U1221_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1222 (
    .clk(delay_reg__U1222_clk),
    .in(delay_reg__U1222_in),
    .out(delay_reg__U1222_out)
);
assign delay_reg__U1223_clk = clk;
assign delay_reg__U1223_in = delay_reg__U1222_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1223 (
    .clk(delay_reg__U1223_clk),
    .in(delay_reg__U1223_in),
    .out(delay_reg__U1223_out)
);
assign delay_reg__U1377_clk = clk;
assign delay_reg__U1377_in = op_hcompute_conv_stencil_13_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1377 (
    .clk(delay_reg__U1377_clk),
    .in(delay_reg__U1377_in),
    .out(delay_reg__U1377_out)
);
assign delay_reg__U1378_clk = clk;
assign delay_reg__U1378_in = delay_reg__U1377_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1378 (
    .clk(delay_reg__U1378_clk),
    .in(delay_reg__U1378_in),
    .out(delay_reg__U1378_out)
);
assign delay_reg__U1395_clk = clk;
assign delay_reg__U1395_in = op_hcompute_conv_stencil_13_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1395 (
    .clk(delay_reg__U1395_clk),
    .in(delay_reg__U1395_in),
    .out(delay_reg__U1395_out)
);
assign delay_reg__U1396_clk = clk;
assign delay_reg__U1396_in = delay_reg__U1395_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1396 (
    .clk(delay_reg__U1396_clk),
    .in(delay_reg__U1396_in),
    .out(delay_reg__U1396_out)
);
assign delay_reg__U1397_clk = clk;
assign delay_reg__U1397_in = delay_reg__U1396_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1397 (
    .clk(delay_reg__U1397_clk),
    .in(delay_reg__U1397_in),
    .out(delay_reg__U1397_out)
);
assign delay_reg__U1398_clk = clk;
assign delay_reg__U1398_in = delay_reg__U1397_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1398 (
    .clk(delay_reg__U1398_clk),
    .in(delay_reg__U1398_in),
    .out(delay_reg__U1398_out)
);
assign delay_reg__U1399_clk = clk;
assign delay_reg__U1399_in = delay_reg__U1398_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1399 (
    .clk(delay_reg__U1399_clk),
    .in(delay_reg__U1399_in),
    .out(delay_reg__U1399_out)
);
assign delay_reg__U1400_clk = clk;
assign delay_reg__U1400_in = delay_reg__U1399_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1400 (
    .clk(delay_reg__U1400_clk),
    .in(delay_reg__U1400_in),
    .out(delay_reg__U1400_out)
);
assign delay_reg__U1401_clk = clk;
assign delay_reg__U1401_in = delay_reg__U1400_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1401 (
    .clk(delay_reg__U1401_clk),
    .in(delay_reg__U1401_in),
    .out(delay_reg__U1401_out)
);
assign delay_reg__U1402_clk = clk;
assign delay_reg__U1402_in = delay_reg__U1401_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1402 (
    .clk(delay_reg__U1402_clk),
    .in(delay_reg__U1402_in),
    .out(delay_reg__U1402_out)
);
assign delay_reg__U1403_clk = clk;
assign delay_reg__U1403_in = delay_reg__U1402_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1403 (
    .clk(delay_reg__U1403_clk),
    .in(delay_reg__U1403_in),
    .out(delay_reg__U1403_out)
);
assign delay_reg__U1404_clk = clk;
assign delay_reg__U1404_in = delay_reg__U1403_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1404 (
    .clk(delay_reg__U1404_clk),
    .in(delay_reg__U1404_in),
    .out(delay_reg__U1404_out)
);
assign delay_reg__U1405_clk = clk;
assign delay_reg__U1405_in = delay_reg__U1404_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1405 (
    .clk(delay_reg__U1405_clk),
    .in(delay_reg__U1405_in),
    .out(delay_reg__U1405_out)
);
assign delay_reg__U1406_clk = clk;
assign delay_reg__U1406_in = delay_reg__U1405_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1406 (
    .clk(delay_reg__U1406_clk),
    .in(delay_reg__U1406_in),
    .out(delay_reg__U1406_out)
);
assign delay_reg__U1407_clk = clk;
assign delay_reg__U1407_in = delay_reg__U1406_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1407 (
    .clk(delay_reg__U1407_clk),
    .in(delay_reg__U1407_in),
    .out(delay_reg__U1407_out)
);
assign delay_reg__U1408_clk = clk;
assign delay_reg__U1408_in = delay_reg__U1407_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1408 (
    .clk(delay_reg__U1408_clk),
    .in(delay_reg__U1408_in),
    .out(delay_reg__U1408_out)
);
assign delay_reg__U1409_clk = clk;
assign delay_reg__U1409_in = delay_reg__U1408_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1409 (
    .clk(delay_reg__U1409_clk),
    .in(delay_reg__U1409_in),
    .out(delay_reg__U1409_out)
);
assign delay_reg__U1410_clk = clk;
assign delay_reg__U1410_in = delay_reg__U1409_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1410 (
    .clk(delay_reg__U1410_clk),
    .in(delay_reg__U1410_in),
    .out(delay_reg__U1410_out)
);
assign delay_reg__U1411_clk = clk;
assign delay_reg__U1411_in = delay_reg__U1410_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1411 (
    .clk(delay_reg__U1411_clk),
    .in(delay_reg__U1411_in),
    .out(delay_reg__U1411_out)
);
assign delay_reg__U1565_clk = clk;
assign delay_reg__U1565_in = op_hcompute_conv_stencil_14_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1565 (
    .clk(delay_reg__U1565_clk),
    .in(delay_reg__U1565_in),
    .out(delay_reg__U1565_out)
);
assign delay_reg__U1566_clk = clk;
assign delay_reg__U1566_in = delay_reg__U1565_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1566 (
    .clk(delay_reg__U1566_clk),
    .in(delay_reg__U1566_in),
    .out(delay_reg__U1566_out)
);
assign delay_reg__U1583_clk = clk;
assign delay_reg__U1583_in = op_hcompute_conv_stencil_14_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1583 (
    .clk(delay_reg__U1583_clk),
    .in(delay_reg__U1583_in),
    .out(delay_reg__U1583_out)
);
assign delay_reg__U1584_clk = clk;
assign delay_reg__U1584_in = delay_reg__U1583_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1584 (
    .clk(delay_reg__U1584_clk),
    .in(delay_reg__U1584_in),
    .out(delay_reg__U1584_out)
);
assign delay_reg__U1585_clk = clk;
assign delay_reg__U1585_in = delay_reg__U1584_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1585 (
    .clk(delay_reg__U1585_clk),
    .in(delay_reg__U1585_in),
    .out(delay_reg__U1585_out)
);
assign delay_reg__U1586_clk = clk;
assign delay_reg__U1586_in = delay_reg__U1585_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1586 (
    .clk(delay_reg__U1586_clk),
    .in(delay_reg__U1586_in),
    .out(delay_reg__U1586_out)
);
assign delay_reg__U1587_clk = clk;
assign delay_reg__U1587_in = delay_reg__U1586_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1587 (
    .clk(delay_reg__U1587_clk),
    .in(delay_reg__U1587_in),
    .out(delay_reg__U1587_out)
);
assign delay_reg__U1588_clk = clk;
assign delay_reg__U1588_in = delay_reg__U1587_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1588 (
    .clk(delay_reg__U1588_clk),
    .in(delay_reg__U1588_in),
    .out(delay_reg__U1588_out)
);
assign delay_reg__U1589_clk = clk;
assign delay_reg__U1589_in = delay_reg__U1588_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1589 (
    .clk(delay_reg__U1589_clk),
    .in(delay_reg__U1589_in),
    .out(delay_reg__U1589_out)
);
assign delay_reg__U1590_clk = clk;
assign delay_reg__U1590_in = delay_reg__U1589_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1590 (
    .clk(delay_reg__U1590_clk),
    .in(delay_reg__U1590_in),
    .out(delay_reg__U1590_out)
);
assign delay_reg__U1591_clk = clk;
assign delay_reg__U1591_in = delay_reg__U1590_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1591 (
    .clk(delay_reg__U1591_clk),
    .in(delay_reg__U1591_in),
    .out(delay_reg__U1591_out)
);
assign delay_reg__U1592_clk = clk;
assign delay_reg__U1592_in = delay_reg__U1591_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1592 (
    .clk(delay_reg__U1592_clk),
    .in(delay_reg__U1592_in),
    .out(delay_reg__U1592_out)
);
assign delay_reg__U1593_clk = clk;
assign delay_reg__U1593_in = delay_reg__U1592_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1593 (
    .clk(delay_reg__U1593_clk),
    .in(delay_reg__U1593_in),
    .out(delay_reg__U1593_out)
);
assign delay_reg__U1594_clk = clk;
assign delay_reg__U1594_in = delay_reg__U1593_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1594 (
    .clk(delay_reg__U1594_clk),
    .in(delay_reg__U1594_in),
    .out(delay_reg__U1594_out)
);
assign delay_reg__U1595_clk = clk;
assign delay_reg__U1595_in = delay_reg__U1594_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1595 (
    .clk(delay_reg__U1595_clk),
    .in(delay_reg__U1595_in),
    .out(delay_reg__U1595_out)
);
assign delay_reg__U1596_clk = clk;
assign delay_reg__U1596_in = delay_reg__U1595_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1596 (
    .clk(delay_reg__U1596_clk),
    .in(delay_reg__U1596_in),
    .out(delay_reg__U1596_out)
);
assign delay_reg__U1597_clk = clk;
assign delay_reg__U1597_in = delay_reg__U1596_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1597 (
    .clk(delay_reg__U1597_clk),
    .in(delay_reg__U1597_in),
    .out(delay_reg__U1597_out)
);
assign delay_reg__U1598_clk = clk;
assign delay_reg__U1598_in = delay_reg__U1597_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1598 (
    .clk(delay_reg__U1598_clk),
    .in(delay_reg__U1598_in),
    .out(delay_reg__U1598_out)
);
assign delay_reg__U1599_clk = clk;
assign delay_reg__U1599_in = delay_reg__U1598_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1599 (
    .clk(delay_reg__U1599_clk),
    .in(delay_reg__U1599_in),
    .out(delay_reg__U1599_out)
);
assign delay_reg__U1753_clk = clk;
assign delay_reg__U1753_in = op_hcompute_conv_stencil_15_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1753 (
    .clk(delay_reg__U1753_clk),
    .in(delay_reg__U1753_in),
    .out(delay_reg__U1753_out)
);
assign delay_reg__U1754_clk = clk;
assign delay_reg__U1754_in = delay_reg__U1753_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1754 (
    .clk(delay_reg__U1754_clk),
    .in(delay_reg__U1754_in),
    .out(delay_reg__U1754_out)
);
assign delay_reg__U1771_clk = clk;
assign delay_reg__U1771_in = op_hcompute_conv_stencil_15_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1771 (
    .clk(delay_reg__U1771_clk),
    .in(delay_reg__U1771_in),
    .out(delay_reg__U1771_out)
);
assign delay_reg__U1772_clk = clk;
assign delay_reg__U1772_in = delay_reg__U1771_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1772 (
    .clk(delay_reg__U1772_clk),
    .in(delay_reg__U1772_in),
    .out(delay_reg__U1772_out)
);
assign delay_reg__U1773_clk = clk;
assign delay_reg__U1773_in = delay_reg__U1772_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1773 (
    .clk(delay_reg__U1773_clk),
    .in(delay_reg__U1773_in),
    .out(delay_reg__U1773_out)
);
assign delay_reg__U1774_clk = clk;
assign delay_reg__U1774_in = delay_reg__U1773_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1774 (
    .clk(delay_reg__U1774_clk),
    .in(delay_reg__U1774_in),
    .out(delay_reg__U1774_out)
);
assign delay_reg__U1775_clk = clk;
assign delay_reg__U1775_in = delay_reg__U1774_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1775 (
    .clk(delay_reg__U1775_clk),
    .in(delay_reg__U1775_in),
    .out(delay_reg__U1775_out)
);
assign delay_reg__U1776_clk = clk;
assign delay_reg__U1776_in = delay_reg__U1775_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1776 (
    .clk(delay_reg__U1776_clk),
    .in(delay_reg__U1776_in),
    .out(delay_reg__U1776_out)
);
assign delay_reg__U1777_clk = clk;
assign delay_reg__U1777_in = delay_reg__U1776_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1777 (
    .clk(delay_reg__U1777_clk),
    .in(delay_reg__U1777_in),
    .out(delay_reg__U1777_out)
);
assign delay_reg__U1778_clk = clk;
assign delay_reg__U1778_in = delay_reg__U1777_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1778 (
    .clk(delay_reg__U1778_clk),
    .in(delay_reg__U1778_in),
    .out(delay_reg__U1778_out)
);
assign delay_reg__U1779_clk = clk;
assign delay_reg__U1779_in = delay_reg__U1778_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1779 (
    .clk(delay_reg__U1779_clk),
    .in(delay_reg__U1779_in),
    .out(delay_reg__U1779_out)
);
assign delay_reg__U1780_clk = clk;
assign delay_reg__U1780_in = delay_reg__U1779_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1780 (
    .clk(delay_reg__U1780_clk),
    .in(delay_reg__U1780_in),
    .out(delay_reg__U1780_out)
);
assign delay_reg__U1781_clk = clk;
assign delay_reg__U1781_in = delay_reg__U1780_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1781 (
    .clk(delay_reg__U1781_clk),
    .in(delay_reg__U1781_in),
    .out(delay_reg__U1781_out)
);
assign delay_reg__U1782_clk = clk;
assign delay_reg__U1782_in = delay_reg__U1781_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1782 (
    .clk(delay_reg__U1782_clk),
    .in(delay_reg__U1782_in),
    .out(delay_reg__U1782_out)
);
assign delay_reg__U1783_clk = clk;
assign delay_reg__U1783_in = delay_reg__U1782_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1783 (
    .clk(delay_reg__U1783_clk),
    .in(delay_reg__U1783_in),
    .out(delay_reg__U1783_out)
);
assign delay_reg__U1784_clk = clk;
assign delay_reg__U1784_in = delay_reg__U1783_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1784 (
    .clk(delay_reg__U1784_clk),
    .in(delay_reg__U1784_in),
    .out(delay_reg__U1784_out)
);
assign delay_reg__U1785_clk = clk;
assign delay_reg__U1785_in = delay_reg__U1784_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1785 (
    .clk(delay_reg__U1785_clk),
    .in(delay_reg__U1785_in),
    .out(delay_reg__U1785_out)
);
assign delay_reg__U1786_clk = clk;
assign delay_reg__U1786_in = delay_reg__U1785_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1786 (
    .clk(delay_reg__U1786_clk),
    .in(delay_reg__U1786_in),
    .out(delay_reg__U1786_out)
);
assign delay_reg__U1787_clk = clk;
assign delay_reg__U1787_in = delay_reg__U1786_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1787 (
    .clk(delay_reg__U1787_clk),
    .in(delay_reg__U1787_in),
    .out(delay_reg__U1787_out)
);
assign delay_reg__U1928_clk = clk;
assign delay_reg__U1928_in = op_hcompute_hw_output_stencil_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1928 (
    .clk(delay_reg__U1928_clk),
    .in(delay_reg__U1928_in),
    .out(delay_reg__U1928_out)
);
assign delay_reg__U1929_clk = clk;
assign delay_reg__U1929_in = delay_reg__U1928_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1929 (
    .clk(delay_reg__U1929_clk),
    .in(delay_reg__U1929_in),
    .out(delay_reg__U1929_out)
);
assign delay_reg__U1942_clk = clk;
assign delay_reg__U1942_in = op_hcompute_hw_output_stencil_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1942 (
    .clk(delay_reg__U1942_clk),
    .in(delay_reg__U1942_in),
    .out(delay_reg__U1942_out)
);
assign delay_reg__U1943_clk = clk;
assign delay_reg__U1943_in = delay_reg__U1942_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1943 (
    .clk(delay_reg__U1943_clk),
    .in(delay_reg__U1943_in),
    .out(delay_reg__U1943_out)
);
assign delay_reg__U1975_clk = clk;
assign delay_reg__U1975_in = op_hcompute_hw_output_stencil_1_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1975 (
    .clk(delay_reg__U1975_clk),
    .in(delay_reg__U1975_in),
    .out(delay_reg__U1975_out)
);
assign delay_reg__U1976_clk = clk;
assign delay_reg__U1976_in = delay_reg__U1975_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1976 (
    .clk(delay_reg__U1976_clk),
    .in(delay_reg__U1976_in),
    .out(delay_reg__U1976_out)
);
assign delay_reg__U1989_clk = clk;
assign delay_reg__U1989_in = op_hcompute_hw_output_stencil_1_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1989 (
    .clk(delay_reg__U1989_clk),
    .in(delay_reg__U1989_in),
    .out(delay_reg__U1989_out)
);
assign delay_reg__U1990_clk = clk;
assign delay_reg__U1990_in = delay_reg__U1989_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U1990 (
    .clk(delay_reg__U1990_clk),
    .in(delay_reg__U1990_in),
    .out(delay_reg__U1990_out)
);
assign delay_reg__U2022_clk = clk;
assign delay_reg__U2022_in = op_hcompute_hw_output_stencil_2_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2022 (
    .clk(delay_reg__U2022_clk),
    .in(delay_reg__U2022_in),
    .out(delay_reg__U2022_out)
);
assign delay_reg__U2023_clk = clk;
assign delay_reg__U2023_in = delay_reg__U2022_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2023 (
    .clk(delay_reg__U2023_clk),
    .in(delay_reg__U2023_in),
    .out(delay_reg__U2023_out)
);
assign delay_reg__U2036_clk = clk;
assign delay_reg__U2036_in = op_hcompute_hw_output_stencil_2_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2036 (
    .clk(delay_reg__U2036_clk),
    .in(delay_reg__U2036_in),
    .out(delay_reg__U2036_out)
);
assign delay_reg__U2037_clk = clk;
assign delay_reg__U2037_in = delay_reg__U2036_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2037 (
    .clk(delay_reg__U2037_clk),
    .in(delay_reg__U2037_in),
    .out(delay_reg__U2037_out)
);
assign delay_reg__U2069_clk = clk;
assign delay_reg__U2069_in = op_hcompute_hw_output_stencil_3_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2069 (
    .clk(delay_reg__U2069_clk),
    .in(delay_reg__U2069_in),
    .out(delay_reg__U2069_out)
);
assign delay_reg__U2070_clk = clk;
assign delay_reg__U2070_in = delay_reg__U2069_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2070 (
    .clk(delay_reg__U2070_clk),
    .in(delay_reg__U2070_in),
    .out(delay_reg__U2070_out)
);
assign delay_reg__U2083_clk = clk;
assign delay_reg__U2083_in = op_hcompute_hw_output_stencil_3_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2083 (
    .clk(delay_reg__U2083_clk),
    .in(delay_reg__U2083_in),
    .out(delay_reg__U2083_out)
);
assign delay_reg__U2084_clk = clk;
assign delay_reg__U2084_in = delay_reg__U2083_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2084 (
    .clk(delay_reg__U2084_clk),
    .in(delay_reg__U2084_in),
    .out(delay_reg__U2084_out)
);
assign delay_reg__U2116_clk = clk;
assign delay_reg__U2116_in = op_hcompute_hw_output_stencil_4_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2116 (
    .clk(delay_reg__U2116_clk),
    .in(delay_reg__U2116_in),
    .out(delay_reg__U2116_out)
);
assign delay_reg__U2117_clk = clk;
assign delay_reg__U2117_in = delay_reg__U2116_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2117 (
    .clk(delay_reg__U2117_clk),
    .in(delay_reg__U2117_in),
    .out(delay_reg__U2117_out)
);
assign delay_reg__U2130_clk = clk;
assign delay_reg__U2130_in = op_hcompute_hw_output_stencil_4_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2130 (
    .clk(delay_reg__U2130_clk),
    .in(delay_reg__U2130_in),
    .out(delay_reg__U2130_out)
);
assign delay_reg__U2131_clk = clk;
assign delay_reg__U2131_in = delay_reg__U2130_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2131 (
    .clk(delay_reg__U2131_clk),
    .in(delay_reg__U2131_in),
    .out(delay_reg__U2131_out)
);
assign delay_reg__U2163_clk = clk;
assign delay_reg__U2163_in = op_hcompute_hw_output_stencil_5_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2163 (
    .clk(delay_reg__U2163_clk),
    .in(delay_reg__U2163_in),
    .out(delay_reg__U2163_out)
);
assign delay_reg__U2164_clk = clk;
assign delay_reg__U2164_in = delay_reg__U2163_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2164 (
    .clk(delay_reg__U2164_clk),
    .in(delay_reg__U2164_in),
    .out(delay_reg__U2164_out)
);
assign delay_reg__U2177_clk = clk;
assign delay_reg__U2177_in = op_hcompute_hw_output_stencil_5_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2177 (
    .clk(delay_reg__U2177_clk),
    .in(delay_reg__U2177_in),
    .out(delay_reg__U2177_out)
);
assign delay_reg__U2178_clk = clk;
assign delay_reg__U2178_in = delay_reg__U2177_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2178 (
    .clk(delay_reg__U2178_clk),
    .in(delay_reg__U2178_in),
    .out(delay_reg__U2178_out)
);
assign delay_reg__U2210_clk = clk;
assign delay_reg__U2210_in = op_hcompute_hw_output_stencil_6_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2210 (
    .clk(delay_reg__U2210_clk),
    .in(delay_reg__U2210_in),
    .out(delay_reg__U2210_out)
);
assign delay_reg__U2211_clk = clk;
assign delay_reg__U2211_in = delay_reg__U2210_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2211 (
    .clk(delay_reg__U2211_clk),
    .in(delay_reg__U2211_in),
    .out(delay_reg__U2211_out)
);
assign delay_reg__U2224_clk = clk;
assign delay_reg__U2224_in = op_hcompute_hw_output_stencil_6_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2224 (
    .clk(delay_reg__U2224_clk),
    .in(delay_reg__U2224_in),
    .out(delay_reg__U2224_out)
);
assign delay_reg__U2225_clk = clk;
assign delay_reg__U2225_in = delay_reg__U2224_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2225 (
    .clk(delay_reg__U2225_clk),
    .in(delay_reg__U2225_in),
    .out(delay_reg__U2225_out)
);
assign delay_reg__U2257_clk = clk;
assign delay_reg__U2257_in = op_hcompute_hw_output_stencil_7_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2257 (
    .clk(delay_reg__U2257_clk),
    .in(delay_reg__U2257_in),
    .out(delay_reg__U2257_out)
);
assign delay_reg__U2258_clk = clk;
assign delay_reg__U2258_in = delay_reg__U2257_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2258 (
    .clk(delay_reg__U2258_clk),
    .in(delay_reg__U2258_in),
    .out(delay_reg__U2258_out)
);
assign delay_reg__U2271_clk = clk;
assign delay_reg__U2271_in = op_hcompute_hw_output_stencil_7_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2271 (
    .clk(delay_reg__U2271_clk),
    .in(delay_reg__U2271_in),
    .out(delay_reg__U2271_out)
);
assign delay_reg__U2272_clk = clk;
assign delay_reg__U2272_in = delay_reg__U2271_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U2272 (
    .clk(delay_reg__U2272_clk),
    .in(delay_reg__U2272_in),
    .out(delay_reg__U2272_out)
);
assign delay_reg__U437_clk = clk;
assign delay_reg__U437_in = op_hcompute_conv_stencil_8_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U437 (
    .clk(delay_reg__U437_clk),
    .in(delay_reg__U437_in),
    .out(delay_reg__U437_out)
);
assign delay_reg__U438_clk = clk;
assign delay_reg__U438_in = delay_reg__U437_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U438 (
    .clk(delay_reg__U438_clk),
    .in(delay_reg__U438_in),
    .out(delay_reg__U438_out)
);
assign delay_reg__U455_clk = clk;
assign delay_reg__U455_in = op_hcompute_conv_stencil_8_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U455 (
    .clk(delay_reg__U455_clk),
    .in(delay_reg__U455_in),
    .out(delay_reg__U455_out)
);
assign delay_reg__U456_clk = clk;
assign delay_reg__U456_in = delay_reg__U455_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U456 (
    .clk(delay_reg__U456_clk),
    .in(delay_reg__U456_in),
    .out(delay_reg__U456_out)
);
assign delay_reg__U457_clk = clk;
assign delay_reg__U457_in = delay_reg__U456_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U457 (
    .clk(delay_reg__U457_clk),
    .in(delay_reg__U457_in),
    .out(delay_reg__U457_out)
);
assign delay_reg__U458_clk = clk;
assign delay_reg__U458_in = delay_reg__U457_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U458 (
    .clk(delay_reg__U458_clk),
    .in(delay_reg__U458_in),
    .out(delay_reg__U458_out)
);
assign delay_reg__U459_clk = clk;
assign delay_reg__U459_in = delay_reg__U458_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U459 (
    .clk(delay_reg__U459_clk),
    .in(delay_reg__U459_in),
    .out(delay_reg__U459_out)
);
assign delay_reg__U460_clk = clk;
assign delay_reg__U460_in = delay_reg__U459_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U460 (
    .clk(delay_reg__U460_clk),
    .in(delay_reg__U460_in),
    .out(delay_reg__U460_out)
);
assign delay_reg__U461_clk = clk;
assign delay_reg__U461_in = delay_reg__U460_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U461 (
    .clk(delay_reg__U461_clk),
    .in(delay_reg__U461_in),
    .out(delay_reg__U461_out)
);
assign delay_reg__U462_clk = clk;
assign delay_reg__U462_in = delay_reg__U461_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U462 (
    .clk(delay_reg__U462_clk),
    .in(delay_reg__U462_in),
    .out(delay_reg__U462_out)
);
assign delay_reg__U463_clk = clk;
assign delay_reg__U463_in = delay_reg__U462_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U463 (
    .clk(delay_reg__U463_clk),
    .in(delay_reg__U463_in),
    .out(delay_reg__U463_out)
);
assign delay_reg__U464_clk = clk;
assign delay_reg__U464_in = delay_reg__U463_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U464 (
    .clk(delay_reg__U464_clk),
    .in(delay_reg__U464_in),
    .out(delay_reg__U464_out)
);
assign delay_reg__U465_clk = clk;
assign delay_reg__U465_in = delay_reg__U464_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U465 (
    .clk(delay_reg__U465_clk),
    .in(delay_reg__U465_in),
    .out(delay_reg__U465_out)
);
assign delay_reg__U466_clk = clk;
assign delay_reg__U466_in = delay_reg__U465_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U466 (
    .clk(delay_reg__U466_clk),
    .in(delay_reg__U466_in),
    .out(delay_reg__U466_out)
);
assign delay_reg__U467_clk = clk;
assign delay_reg__U467_in = delay_reg__U466_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U467 (
    .clk(delay_reg__U467_clk),
    .in(delay_reg__U467_in),
    .out(delay_reg__U467_out)
);
assign delay_reg__U468_clk = clk;
assign delay_reg__U468_in = delay_reg__U467_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U468 (
    .clk(delay_reg__U468_clk),
    .in(delay_reg__U468_in),
    .out(delay_reg__U468_out)
);
assign delay_reg__U469_clk = clk;
assign delay_reg__U469_in = delay_reg__U468_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U469 (
    .clk(delay_reg__U469_clk),
    .in(delay_reg__U469_in),
    .out(delay_reg__U469_out)
);
assign delay_reg__U470_clk = clk;
assign delay_reg__U470_in = delay_reg__U469_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U470 (
    .clk(delay_reg__U470_clk),
    .in(delay_reg__U470_in),
    .out(delay_reg__U470_out)
);
assign delay_reg__U471_clk = clk;
assign delay_reg__U471_in = delay_reg__U470_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U471 (
    .clk(delay_reg__U471_clk),
    .in(delay_reg__U471_in),
    .out(delay_reg__U471_out)
);
assign delay_reg__U625_clk = clk;
assign delay_reg__U625_in = op_hcompute_conv_stencil_9_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U625 (
    .clk(delay_reg__U625_clk),
    .in(delay_reg__U625_in),
    .out(delay_reg__U625_out)
);
assign delay_reg__U626_clk = clk;
assign delay_reg__U626_in = delay_reg__U625_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U626 (
    .clk(delay_reg__U626_clk),
    .in(delay_reg__U626_in),
    .out(delay_reg__U626_out)
);
assign delay_reg__U643_clk = clk;
assign delay_reg__U643_in = op_hcompute_conv_stencil_9_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U643 (
    .clk(delay_reg__U643_clk),
    .in(delay_reg__U643_in),
    .out(delay_reg__U643_out)
);
assign delay_reg__U644_clk = clk;
assign delay_reg__U644_in = delay_reg__U643_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U644 (
    .clk(delay_reg__U644_clk),
    .in(delay_reg__U644_in),
    .out(delay_reg__U644_out)
);
assign delay_reg__U645_clk = clk;
assign delay_reg__U645_in = delay_reg__U644_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U645 (
    .clk(delay_reg__U645_clk),
    .in(delay_reg__U645_in),
    .out(delay_reg__U645_out)
);
assign delay_reg__U646_clk = clk;
assign delay_reg__U646_in = delay_reg__U645_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U646 (
    .clk(delay_reg__U646_clk),
    .in(delay_reg__U646_in),
    .out(delay_reg__U646_out)
);
assign delay_reg__U647_clk = clk;
assign delay_reg__U647_in = delay_reg__U646_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U647 (
    .clk(delay_reg__U647_clk),
    .in(delay_reg__U647_in),
    .out(delay_reg__U647_out)
);
assign delay_reg__U648_clk = clk;
assign delay_reg__U648_in = delay_reg__U647_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U648 (
    .clk(delay_reg__U648_clk),
    .in(delay_reg__U648_in),
    .out(delay_reg__U648_out)
);
assign delay_reg__U649_clk = clk;
assign delay_reg__U649_in = delay_reg__U648_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U649 (
    .clk(delay_reg__U649_clk),
    .in(delay_reg__U649_in),
    .out(delay_reg__U649_out)
);
assign delay_reg__U650_clk = clk;
assign delay_reg__U650_in = delay_reg__U649_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U650 (
    .clk(delay_reg__U650_clk),
    .in(delay_reg__U650_in),
    .out(delay_reg__U650_out)
);
assign delay_reg__U651_clk = clk;
assign delay_reg__U651_in = delay_reg__U650_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U651 (
    .clk(delay_reg__U651_clk),
    .in(delay_reg__U651_in),
    .out(delay_reg__U651_out)
);
assign delay_reg__U652_clk = clk;
assign delay_reg__U652_in = delay_reg__U651_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U652 (
    .clk(delay_reg__U652_clk),
    .in(delay_reg__U652_in),
    .out(delay_reg__U652_out)
);
assign delay_reg__U653_clk = clk;
assign delay_reg__U653_in = delay_reg__U652_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U653 (
    .clk(delay_reg__U653_clk),
    .in(delay_reg__U653_in),
    .out(delay_reg__U653_out)
);
assign delay_reg__U654_clk = clk;
assign delay_reg__U654_in = delay_reg__U653_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U654 (
    .clk(delay_reg__U654_clk),
    .in(delay_reg__U654_in),
    .out(delay_reg__U654_out)
);
assign delay_reg__U655_clk = clk;
assign delay_reg__U655_in = delay_reg__U654_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U655 (
    .clk(delay_reg__U655_clk),
    .in(delay_reg__U655_in),
    .out(delay_reg__U655_out)
);
assign delay_reg__U656_clk = clk;
assign delay_reg__U656_in = delay_reg__U655_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U656 (
    .clk(delay_reg__U656_clk),
    .in(delay_reg__U656_in),
    .out(delay_reg__U656_out)
);
assign delay_reg__U657_clk = clk;
assign delay_reg__U657_in = delay_reg__U656_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U657 (
    .clk(delay_reg__U657_clk),
    .in(delay_reg__U657_in),
    .out(delay_reg__U657_out)
);
assign delay_reg__U658_clk = clk;
assign delay_reg__U658_in = delay_reg__U657_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U658 (
    .clk(delay_reg__U658_clk),
    .in(delay_reg__U658_in),
    .out(delay_reg__U658_out)
);
assign delay_reg__U659_clk = clk;
assign delay_reg__U659_in = delay_reg__U658_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U659 (
    .clk(delay_reg__U659_clk),
    .in(delay_reg__U659_in),
    .out(delay_reg__U659_out)
);
assign delay_reg__U813_clk = clk;
assign delay_reg__U813_in = op_hcompute_conv_stencil_10_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U813 (
    .clk(delay_reg__U813_clk),
    .in(delay_reg__U813_in),
    .out(delay_reg__U813_out)
);
assign delay_reg__U814_clk = clk;
assign delay_reg__U814_in = delay_reg__U813_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U814 (
    .clk(delay_reg__U814_clk),
    .in(delay_reg__U814_in),
    .out(delay_reg__U814_out)
);
assign delay_reg__U831_clk = clk;
assign delay_reg__U831_in = op_hcompute_conv_stencil_10_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U831 (
    .clk(delay_reg__U831_clk),
    .in(delay_reg__U831_in),
    .out(delay_reg__U831_out)
);
assign delay_reg__U832_clk = clk;
assign delay_reg__U832_in = delay_reg__U831_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U832 (
    .clk(delay_reg__U832_clk),
    .in(delay_reg__U832_in),
    .out(delay_reg__U832_out)
);
assign delay_reg__U833_clk = clk;
assign delay_reg__U833_in = delay_reg__U832_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U833 (
    .clk(delay_reg__U833_clk),
    .in(delay_reg__U833_in),
    .out(delay_reg__U833_out)
);
assign delay_reg__U834_clk = clk;
assign delay_reg__U834_in = delay_reg__U833_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U834 (
    .clk(delay_reg__U834_clk),
    .in(delay_reg__U834_in),
    .out(delay_reg__U834_out)
);
assign delay_reg__U835_clk = clk;
assign delay_reg__U835_in = delay_reg__U834_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U835 (
    .clk(delay_reg__U835_clk),
    .in(delay_reg__U835_in),
    .out(delay_reg__U835_out)
);
assign delay_reg__U836_clk = clk;
assign delay_reg__U836_in = delay_reg__U835_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U836 (
    .clk(delay_reg__U836_clk),
    .in(delay_reg__U836_in),
    .out(delay_reg__U836_out)
);
assign delay_reg__U837_clk = clk;
assign delay_reg__U837_in = delay_reg__U836_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U837 (
    .clk(delay_reg__U837_clk),
    .in(delay_reg__U837_in),
    .out(delay_reg__U837_out)
);
assign delay_reg__U838_clk = clk;
assign delay_reg__U838_in = delay_reg__U837_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U838 (
    .clk(delay_reg__U838_clk),
    .in(delay_reg__U838_in),
    .out(delay_reg__U838_out)
);
assign delay_reg__U839_clk = clk;
assign delay_reg__U839_in = delay_reg__U838_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U839 (
    .clk(delay_reg__U839_clk),
    .in(delay_reg__U839_in),
    .out(delay_reg__U839_out)
);
assign delay_reg__U840_clk = clk;
assign delay_reg__U840_in = delay_reg__U839_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U840 (
    .clk(delay_reg__U840_clk),
    .in(delay_reg__U840_in),
    .out(delay_reg__U840_out)
);
assign delay_reg__U841_clk = clk;
assign delay_reg__U841_in = delay_reg__U840_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U841 (
    .clk(delay_reg__U841_clk),
    .in(delay_reg__U841_in),
    .out(delay_reg__U841_out)
);
assign delay_reg__U842_clk = clk;
assign delay_reg__U842_in = delay_reg__U841_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U842 (
    .clk(delay_reg__U842_clk),
    .in(delay_reg__U842_in),
    .out(delay_reg__U842_out)
);
assign delay_reg__U843_clk = clk;
assign delay_reg__U843_in = delay_reg__U842_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U843 (
    .clk(delay_reg__U843_clk),
    .in(delay_reg__U843_in),
    .out(delay_reg__U843_out)
);
assign delay_reg__U844_clk = clk;
assign delay_reg__U844_in = delay_reg__U843_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U844 (
    .clk(delay_reg__U844_clk),
    .in(delay_reg__U844_in),
    .out(delay_reg__U844_out)
);
assign delay_reg__U845_clk = clk;
assign delay_reg__U845_in = delay_reg__U844_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U845 (
    .clk(delay_reg__U845_clk),
    .in(delay_reg__U845_in),
    .out(delay_reg__U845_out)
);
assign delay_reg__U846_clk = clk;
assign delay_reg__U846_in = delay_reg__U845_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U846 (
    .clk(delay_reg__U846_clk),
    .in(delay_reg__U846_in),
    .out(delay_reg__U846_out)
);
assign delay_reg__U847_clk = clk;
assign delay_reg__U847_in = delay_reg__U846_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U847 (
    .clk(delay_reg__U847_clk),
    .in(delay_reg__U847_in),
    .out(delay_reg__U847_out)
);
assign hw_input_global_wrapper_stencil_clk = clk;
assign hw_input_global_wrapper_stencil_flush = flush;
assign hw_input_global_wrapper_stencil_rst_n = rst_n;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ren = op_hcompute_conv_stencil_10_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[4] = op_hcompute_conv_stencil_10_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[3] = op_hcompute_conv_stencil_10_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[2] = op_hcompute_conv_stencil_10_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[1] = op_hcompute_conv_stencil_10_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[0] = op_hcompute_conv_stencil_10_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ren = op_hcompute_conv_stencil_11_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[4] = op_hcompute_conv_stencil_11_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[3] = op_hcompute_conv_stencil_11_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[2] = op_hcompute_conv_stencil_11_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[1] = op_hcompute_conv_stencil_11_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[0] = op_hcompute_conv_stencil_11_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ren = op_hcompute_conv_stencil_12_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[4] = op_hcompute_conv_stencil_12_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[3] = op_hcompute_conv_stencil_12_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[2] = op_hcompute_conv_stencil_12_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[1] = op_hcompute_conv_stencil_12_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[0] = op_hcompute_conv_stencil_12_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ren = op_hcompute_conv_stencil_13_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[4] = op_hcompute_conv_stencil_13_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[3] = op_hcompute_conv_stencil_13_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[2] = op_hcompute_conv_stencil_13_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[1] = op_hcompute_conv_stencil_13_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[0] = op_hcompute_conv_stencil_13_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ren = op_hcompute_conv_stencil_14_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[4] = op_hcompute_conv_stencil_14_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[3] = op_hcompute_conv_stencil_14_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[2] = op_hcompute_conv_stencil_14_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[1] = op_hcompute_conv_stencil_14_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[0] = op_hcompute_conv_stencil_14_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ren = op_hcompute_conv_stencil_15_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[4] = op_hcompute_conv_stencil_15_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[3] = op_hcompute_conv_stencil_15_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[2] = op_hcompute_conv_stencil_15_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[1] = op_hcompute_conv_stencil_15_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[0] = op_hcompute_conv_stencil_15_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ren = op_hcompute_conv_stencil_8_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[4] = op_hcompute_conv_stencil_8_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[3] = op_hcompute_conv_stencil_8_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[2] = op_hcompute_conv_stencil_8_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[1] = op_hcompute_conv_stencil_8_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[0] = op_hcompute_conv_stencil_8_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ren = op_hcompute_conv_stencil_9_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[4] = op_hcompute_conv_stencil_9_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[3] = op_hcompute_conv_stencil_9_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[2] = op_hcompute_conv_stencil_9_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[1] = op_hcompute_conv_stencil_9_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[0] = op_hcompute_conv_stencil_9_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write_wen = op_hcompute_hw_input_global_wrapper_stencil_1_write_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_out[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write[0] = op_hcompute_hw_input_global_wrapper_stencil_1_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write_wen = op_hcompute_hw_input_global_wrapper_stencil_2_write_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_out[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write[0] = op_hcompute_hw_input_global_wrapper_stencil_2_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write_wen = op_hcompute_hw_input_global_wrapper_stencil_3_write_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_out[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write[0] = op_hcompute_hw_input_global_wrapper_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write_wen = op_hcompute_hw_input_global_wrapper_stencil_4_write_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_out[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write[0] = op_hcompute_hw_input_global_wrapper_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write_wen = op_hcompute_hw_input_global_wrapper_stencil_5_write_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_out[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write[0] = op_hcompute_hw_input_global_wrapper_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write_wen = op_hcompute_hw_input_global_wrapper_stencil_6_write_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_out[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write[0] = op_hcompute_hw_input_global_wrapper_stencil_6_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write_wen = op_hcompute_hw_input_global_wrapper_stencil_7_write_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_out[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write[0] = op_hcompute_hw_input_global_wrapper_stencil_7_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen = op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0];
hw_input_global_wrapper_stencil_ub hw_input_global_wrapper_stencil (
    .clk(hw_input_global_wrapper_stencil_clk),
    .flush(hw_input_global_wrapper_stencil_flush),
    .rst_n(hw_input_global_wrapper_stencil_rst_n),
    .op_hcompute_conv_stencil_10_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ren),
    .op_hcompute_conv_stencil_10_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars),
    .op_hcompute_conv_stencil_10_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read),
    .op_hcompute_conv_stencil_11_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ren),
    .op_hcompute_conv_stencil_11_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars),
    .op_hcompute_conv_stencil_11_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read),
    .op_hcompute_conv_stencil_12_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ren),
    .op_hcompute_conv_stencil_12_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars),
    .op_hcompute_conv_stencil_12_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read),
    .op_hcompute_conv_stencil_13_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ren),
    .op_hcompute_conv_stencil_13_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars),
    .op_hcompute_conv_stencil_13_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read),
    .op_hcompute_conv_stencil_14_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ren),
    .op_hcompute_conv_stencil_14_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars),
    .op_hcompute_conv_stencil_14_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read),
    .op_hcompute_conv_stencil_15_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ren),
    .op_hcompute_conv_stencil_15_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars),
    .op_hcompute_conv_stencil_15_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read),
    .op_hcompute_conv_stencil_8_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ren),
    .op_hcompute_conv_stencil_8_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars),
    .op_hcompute_conv_stencil_8_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read),
    .op_hcompute_conv_stencil_9_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ren),
    .op_hcompute_conv_stencil_9_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars),
    .op_hcompute_conv_stencil_9_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read),
    .op_hcompute_hw_input_global_wrapper_stencil_1_write_wen(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write_wen),
    .op_hcompute_hw_input_global_wrapper_stencil_1_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_1_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write),
    .op_hcompute_hw_input_global_wrapper_stencil_2_write_wen(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write_wen),
    .op_hcompute_hw_input_global_wrapper_stencil_2_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_2_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write),
    .op_hcompute_hw_input_global_wrapper_stencil_3_write_wen(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write_wen),
    .op_hcompute_hw_input_global_wrapper_stencil_3_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_3_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write),
    .op_hcompute_hw_input_global_wrapper_stencil_4_write_wen(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write_wen),
    .op_hcompute_hw_input_global_wrapper_stencil_4_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_4_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write),
    .op_hcompute_hw_input_global_wrapper_stencil_5_write_wen(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write_wen),
    .op_hcompute_hw_input_global_wrapper_stencil_5_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_5_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write),
    .op_hcompute_hw_input_global_wrapper_stencil_6_write_wen(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write_wen),
    .op_hcompute_hw_input_global_wrapper_stencil_6_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_6_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write),
    .op_hcompute_hw_input_global_wrapper_stencil_7_write_wen(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write_wen),
    .op_hcompute_hw_input_global_wrapper_stencil_7_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_7_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write),
    .op_hcompute_hw_input_global_wrapper_stencil_write_wen(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen),
    .op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
assign hw_kernel_global_wrapper_stencil_clk = clk;
assign hw_kernel_global_wrapper_stencil_flush = flush;
assign hw_kernel_global_wrapper_stencil_rst_n = rst_n;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ren = op_hcompute_conv_stencil_10_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[4] = op_hcompute_conv_stencil_10_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[3] = op_hcompute_conv_stencil_10_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[2] = op_hcompute_conv_stencil_10_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[1] = op_hcompute_conv_stencil_10_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars[0] = op_hcompute_conv_stencil_10_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ren = op_hcompute_conv_stencil_11_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[4] = op_hcompute_conv_stencil_11_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[3] = op_hcompute_conv_stencil_11_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[2] = op_hcompute_conv_stencil_11_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[1] = op_hcompute_conv_stencil_11_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars[0] = op_hcompute_conv_stencil_11_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ren = op_hcompute_conv_stencil_12_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[4] = op_hcompute_conv_stencil_12_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[3] = op_hcompute_conv_stencil_12_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[2] = op_hcompute_conv_stencil_12_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[1] = op_hcompute_conv_stencil_12_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars[0] = op_hcompute_conv_stencil_12_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ren = op_hcompute_conv_stencil_13_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[4] = op_hcompute_conv_stencil_13_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[3] = op_hcompute_conv_stencil_13_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[2] = op_hcompute_conv_stencil_13_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[1] = op_hcompute_conv_stencil_13_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars[0] = op_hcompute_conv_stencil_13_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ren = op_hcompute_conv_stencil_14_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[4] = op_hcompute_conv_stencil_14_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[3] = op_hcompute_conv_stencil_14_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[2] = op_hcompute_conv_stencil_14_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[1] = op_hcompute_conv_stencil_14_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars[0] = op_hcompute_conv_stencil_14_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ren = op_hcompute_conv_stencil_15_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[4] = op_hcompute_conv_stencil_15_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[3] = op_hcompute_conv_stencil_15_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[2] = op_hcompute_conv_stencil_15_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[1] = op_hcompute_conv_stencil_15_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars[0] = op_hcompute_conv_stencil_15_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ren = op_hcompute_conv_stencil_8_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[4] = op_hcompute_conv_stencil_8_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[3] = op_hcompute_conv_stencil_8_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[2] = op_hcompute_conv_stencil_8_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[1] = op_hcompute_conv_stencil_8_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars[0] = op_hcompute_conv_stencil_8_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ren = op_hcompute_conv_stencil_9_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[4] = op_hcompute_conv_stencil_9_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[3] = op_hcompute_conv_stencil_9_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[2] = op_hcompute_conv_stencil_9_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[1] = op_hcompute_conv_stencil_9_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars[0] = op_hcompute_conv_stencil_9_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[4] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0];
hw_kernel_global_wrapper_stencil_ub hw_kernel_global_wrapper_stencil (
    .clk(hw_kernel_global_wrapper_stencil_clk),
    .flush(hw_kernel_global_wrapper_stencil_flush),
    .rst_n(hw_kernel_global_wrapper_stencil_rst_n),
    .op_hcompute_conv_stencil_10_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ren),
    .op_hcompute_conv_stencil_10_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read_ctrl_vars),
    .op_hcompute_conv_stencil_10_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read),
    .op_hcompute_conv_stencil_11_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ren),
    .op_hcompute_conv_stencil_11_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read_ctrl_vars),
    .op_hcompute_conv_stencil_11_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read),
    .op_hcompute_conv_stencil_12_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ren),
    .op_hcompute_conv_stencil_12_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read_ctrl_vars),
    .op_hcompute_conv_stencil_12_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read),
    .op_hcompute_conv_stencil_13_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ren),
    .op_hcompute_conv_stencil_13_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read_ctrl_vars),
    .op_hcompute_conv_stencil_13_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read),
    .op_hcompute_conv_stencil_14_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ren),
    .op_hcompute_conv_stencil_14_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read_ctrl_vars),
    .op_hcompute_conv_stencil_14_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read),
    .op_hcompute_conv_stencil_15_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ren),
    .op_hcompute_conv_stencil_15_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read_ctrl_vars),
    .op_hcompute_conv_stencil_15_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read),
    .op_hcompute_conv_stencil_8_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ren),
    .op_hcompute_conv_stencil_8_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read_ctrl_vars),
    .op_hcompute_conv_stencil_8_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read),
    .op_hcompute_conv_stencil_9_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ren),
    .op_hcompute_conv_stencil_9_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read_ctrl_vars),
    .op_hcompute_conv_stencil_9_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_wen(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
assign op_hcompute_conv_stencil_clk = clk;
cu_op_hcompute_conv_stencil op_hcompute_conv_stencil (
    .clk(op_hcompute_conv_stencil_clk),
    .conv_stencil_op_hcompute_conv_stencil_write(op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write)
);
assign op_hcompute_conv_stencil_1_clk = clk;
cu_op_hcompute_conv_stencil_1 op_hcompute_conv_stencil_1 (
    .clk(op_hcompute_conv_stencil_1_clk),
    .conv_stencil_op_hcompute_conv_stencil_1_write(op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write)
);
assign op_hcompute_conv_stencil_10_clk = clk;
assign op_hcompute_conv_stencil_10_conv_stencil_op_hcompute_conv_stencil_10_read[0] = conv_stencil_op_hcompute_conv_stencil_10_read[0];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[7];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[6];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[5];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[4];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[3];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[2];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[1];
assign op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[0];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[7];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[6];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[5];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[4];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[3];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[2];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[1];
assign op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read[0];
cu_op_hcompute_conv_stencil_10 op_hcompute_conv_stencil_10 (
    .clk(op_hcompute_conv_stencil_10_clk),
    .conv_stencil_op_hcompute_conv_stencil_10_read(op_hcompute_conv_stencil_10_conv_stencil_op_hcompute_conv_stencil_10_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read(op_hcompute_conv_stencil_10_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_10_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read(op_hcompute_conv_stencil_10_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_10_read),
    .conv_stencil_op_hcompute_conv_stencil_10_write(op_hcompute_conv_stencil_10_conv_stencil_op_hcompute_conv_stencil_10_write)
);
assign op_hcompute_conv_stencil_10_exe_start_in = delay_reg__U814_out;
op_hcompute_conv_stencil_10_exe_start_pt__U812 op_hcompute_conv_stencil_10_exe_start (
    .in(op_hcompute_conv_stencil_10_exe_start_in),
    .out(op_hcompute_conv_stencil_10_exe_start_out)
);
assign op_hcompute_conv_stencil_10_exe_start_control_vars_in[4] = arr__U823_out[4];
assign op_hcompute_conv_stencil_10_exe_start_control_vars_in[3] = arr__U823_out[3];
assign op_hcompute_conv_stencil_10_exe_start_control_vars_in[2] = arr__U823_out[2];
assign op_hcompute_conv_stencil_10_exe_start_control_vars_in[1] = arr__U823_out[1];
assign op_hcompute_conv_stencil_10_exe_start_control_vars_in[0] = arr__U823_out[0];
op_hcompute_conv_stencil_10_exe_start_control_vars_pt__U815 op_hcompute_conv_stencil_10_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_10_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_10_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_10_port_controller_clk = clk;
affine_controller__U780 op_hcompute_conv_stencil_10_port_controller (
    .clk(op_hcompute_conv_stencil_10_port_controller_clk),
    .valid(op_hcompute_conv_stencil_10_port_controller_valid),
    .d(op_hcompute_conv_stencil_10_port_controller_d)
);
assign op_hcompute_conv_stencil_10_read_start_in = op_hcompute_conv_stencil_10_port_controller_valid;
op_hcompute_conv_stencil_10_read_start_pt__U810 op_hcompute_conv_stencil_10_read_start (
    .in(op_hcompute_conv_stencil_10_read_start_in),
    .out(op_hcompute_conv_stencil_10_read_start_out)
);
assign op_hcompute_conv_stencil_10_read_start_control_vars_in[4] = op_hcompute_conv_stencil_10_port_controller_d[4];
assign op_hcompute_conv_stencil_10_read_start_control_vars_in[3] = op_hcompute_conv_stencil_10_port_controller_d[3];
assign op_hcompute_conv_stencil_10_read_start_control_vars_in[2] = op_hcompute_conv_stencil_10_port_controller_d[2];
assign op_hcompute_conv_stencil_10_read_start_control_vars_in[1] = op_hcompute_conv_stencil_10_port_controller_d[1];
assign op_hcompute_conv_stencil_10_read_start_control_vars_in[0] = op_hcompute_conv_stencil_10_port_controller_d[0];
op_hcompute_conv_stencil_10_read_start_control_vars_pt__U811 op_hcompute_conv_stencil_10_read_start_control_vars (
    .in(op_hcompute_conv_stencil_10_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_10_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_10_write_start_in = delay_reg__U847_out;
op_hcompute_conv_stencil_10_write_start_pt__U830 op_hcompute_conv_stencil_10_write_start (
    .in(op_hcompute_conv_stencil_10_write_start_in),
    .out(op_hcompute_conv_stencil_10_write_start_out)
);
assign op_hcompute_conv_stencil_10_write_start_control_vars_in[4] = arr__U961_out[4];
assign op_hcompute_conv_stencil_10_write_start_control_vars_in[3] = arr__U961_out[3];
assign op_hcompute_conv_stencil_10_write_start_control_vars_in[2] = arr__U961_out[2];
assign op_hcompute_conv_stencil_10_write_start_control_vars_in[1] = arr__U961_out[1];
assign op_hcompute_conv_stencil_10_write_start_control_vars_in[0] = arr__U961_out[0];
op_hcompute_conv_stencil_10_write_start_control_vars_pt__U848 op_hcompute_conv_stencil_10_write_start_control_vars (
    .in(op_hcompute_conv_stencil_10_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_10_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_11_clk = clk;
assign op_hcompute_conv_stencil_11_conv_stencil_op_hcompute_conv_stencil_11_read[0] = conv_stencil_op_hcompute_conv_stencil_11_read[0];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[7];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[6];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[5];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[4];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[3];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[2];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[1];
assign op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[0];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[7];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[6];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[5];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[4];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[3];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[2];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[1];
assign op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read[0];
cu_op_hcompute_conv_stencil_11 op_hcompute_conv_stencil_11 (
    .clk(op_hcompute_conv_stencil_11_clk),
    .conv_stencil_op_hcompute_conv_stencil_11_read(op_hcompute_conv_stencil_11_conv_stencil_op_hcompute_conv_stencil_11_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read(op_hcompute_conv_stencil_11_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_11_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read(op_hcompute_conv_stencil_11_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_11_read),
    .conv_stencil_op_hcompute_conv_stencil_11_write(op_hcompute_conv_stencil_11_conv_stencil_op_hcompute_conv_stencil_11_write)
);
assign op_hcompute_conv_stencil_11_exe_start_in = delay_reg__U1002_out;
op_hcompute_conv_stencil_11_exe_start_pt__U1000 op_hcompute_conv_stencil_11_exe_start (
    .in(op_hcompute_conv_stencil_11_exe_start_in),
    .out(op_hcompute_conv_stencil_11_exe_start_out)
);
assign op_hcompute_conv_stencil_11_exe_start_control_vars_in[4] = arr__U1011_out[4];
assign op_hcompute_conv_stencil_11_exe_start_control_vars_in[3] = arr__U1011_out[3];
assign op_hcompute_conv_stencil_11_exe_start_control_vars_in[2] = arr__U1011_out[2];
assign op_hcompute_conv_stencil_11_exe_start_control_vars_in[1] = arr__U1011_out[1];
assign op_hcompute_conv_stencil_11_exe_start_control_vars_in[0] = arr__U1011_out[0];
op_hcompute_conv_stencil_11_exe_start_control_vars_pt__U1003 op_hcompute_conv_stencil_11_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_11_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_11_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_11_port_controller_clk = clk;
affine_controller__U968 op_hcompute_conv_stencil_11_port_controller (
    .clk(op_hcompute_conv_stencil_11_port_controller_clk),
    .valid(op_hcompute_conv_stencil_11_port_controller_valid),
    .d(op_hcompute_conv_stencil_11_port_controller_d)
);
assign op_hcompute_conv_stencil_11_read_start_in = op_hcompute_conv_stencil_11_port_controller_valid;
op_hcompute_conv_stencil_11_read_start_pt__U998 op_hcompute_conv_stencil_11_read_start (
    .in(op_hcompute_conv_stencil_11_read_start_in),
    .out(op_hcompute_conv_stencil_11_read_start_out)
);
assign op_hcompute_conv_stencil_11_read_start_control_vars_in[4] = op_hcompute_conv_stencil_11_port_controller_d[4];
assign op_hcompute_conv_stencil_11_read_start_control_vars_in[3] = op_hcompute_conv_stencil_11_port_controller_d[3];
assign op_hcompute_conv_stencil_11_read_start_control_vars_in[2] = op_hcompute_conv_stencil_11_port_controller_d[2];
assign op_hcompute_conv_stencil_11_read_start_control_vars_in[1] = op_hcompute_conv_stencil_11_port_controller_d[1];
assign op_hcompute_conv_stencil_11_read_start_control_vars_in[0] = op_hcompute_conv_stencil_11_port_controller_d[0];
op_hcompute_conv_stencil_11_read_start_control_vars_pt__U999 op_hcompute_conv_stencil_11_read_start_control_vars (
    .in(op_hcompute_conv_stencil_11_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_11_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_11_write_start_in = delay_reg__U1035_out;
op_hcompute_conv_stencil_11_write_start_pt__U1018 op_hcompute_conv_stencil_11_write_start (
    .in(op_hcompute_conv_stencil_11_write_start_in),
    .out(op_hcompute_conv_stencil_11_write_start_out)
);
assign op_hcompute_conv_stencil_11_write_start_control_vars_in[4] = arr__U1149_out[4];
assign op_hcompute_conv_stencil_11_write_start_control_vars_in[3] = arr__U1149_out[3];
assign op_hcompute_conv_stencil_11_write_start_control_vars_in[2] = arr__U1149_out[2];
assign op_hcompute_conv_stencil_11_write_start_control_vars_in[1] = arr__U1149_out[1];
assign op_hcompute_conv_stencil_11_write_start_control_vars_in[0] = arr__U1149_out[0];
op_hcompute_conv_stencil_11_write_start_control_vars_pt__U1036 op_hcompute_conv_stencil_11_write_start_control_vars (
    .in(op_hcompute_conv_stencil_11_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_11_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_12_clk = clk;
assign op_hcompute_conv_stencil_12_conv_stencil_op_hcompute_conv_stencil_12_read[0] = conv_stencil_op_hcompute_conv_stencil_12_read[0];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[7];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[6];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[5];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[4];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[3];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[2];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[1];
assign op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[0];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[7];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[6];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[5];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[4];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[3];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[2];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[1];
assign op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read[0];
cu_op_hcompute_conv_stencil_12 op_hcompute_conv_stencil_12 (
    .clk(op_hcompute_conv_stencil_12_clk),
    .conv_stencil_op_hcompute_conv_stencil_12_read(op_hcompute_conv_stencil_12_conv_stencil_op_hcompute_conv_stencil_12_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read(op_hcompute_conv_stencil_12_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_12_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read(op_hcompute_conv_stencil_12_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_12_read),
    .conv_stencil_op_hcompute_conv_stencil_12_write(op_hcompute_conv_stencil_12_conv_stencil_op_hcompute_conv_stencil_12_write)
);
assign op_hcompute_conv_stencil_12_exe_start_in = delay_reg__U1190_out;
op_hcompute_conv_stencil_12_exe_start_pt__U1188 op_hcompute_conv_stencil_12_exe_start (
    .in(op_hcompute_conv_stencil_12_exe_start_in),
    .out(op_hcompute_conv_stencil_12_exe_start_out)
);
assign op_hcompute_conv_stencil_12_exe_start_control_vars_in[4] = arr__U1199_out[4];
assign op_hcompute_conv_stencil_12_exe_start_control_vars_in[3] = arr__U1199_out[3];
assign op_hcompute_conv_stencil_12_exe_start_control_vars_in[2] = arr__U1199_out[2];
assign op_hcompute_conv_stencil_12_exe_start_control_vars_in[1] = arr__U1199_out[1];
assign op_hcompute_conv_stencil_12_exe_start_control_vars_in[0] = arr__U1199_out[0];
op_hcompute_conv_stencil_12_exe_start_control_vars_pt__U1191 op_hcompute_conv_stencil_12_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_12_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_12_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_12_port_controller_clk = clk;
affine_controller__U1156 op_hcompute_conv_stencil_12_port_controller (
    .clk(op_hcompute_conv_stencil_12_port_controller_clk),
    .valid(op_hcompute_conv_stencil_12_port_controller_valid),
    .d(op_hcompute_conv_stencil_12_port_controller_d)
);
assign op_hcompute_conv_stencil_12_read_start_in = op_hcompute_conv_stencil_12_port_controller_valid;
op_hcompute_conv_stencil_12_read_start_pt__U1186 op_hcompute_conv_stencil_12_read_start (
    .in(op_hcompute_conv_stencil_12_read_start_in),
    .out(op_hcompute_conv_stencil_12_read_start_out)
);
assign op_hcompute_conv_stencil_12_read_start_control_vars_in[4] = op_hcompute_conv_stencil_12_port_controller_d[4];
assign op_hcompute_conv_stencil_12_read_start_control_vars_in[3] = op_hcompute_conv_stencil_12_port_controller_d[3];
assign op_hcompute_conv_stencil_12_read_start_control_vars_in[2] = op_hcompute_conv_stencil_12_port_controller_d[2];
assign op_hcompute_conv_stencil_12_read_start_control_vars_in[1] = op_hcompute_conv_stencil_12_port_controller_d[1];
assign op_hcompute_conv_stencil_12_read_start_control_vars_in[0] = op_hcompute_conv_stencil_12_port_controller_d[0];
op_hcompute_conv_stencil_12_read_start_control_vars_pt__U1187 op_hcompute_conv_stencil_12_read_start_control_vars (
    .in(op_hcompute_conv_stencil_12_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_12_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_12_write_start_in = delay_reg__U1223_out;
op_hcompute_conv_stencil_12_write_start_pt__U1206 op_hcompute_conv_stencil_12_write_start (
    .in(op_hcompute_conv_stencil_12_write_start_in),
    .out(op_hcompute_conv_stencil_12_write_start_out)
);
assign op_hcompute_conv_stencil_12_write_start_control_vars_in[4] = arr__U1337_out[4];
assign op_hcompute_conv_stencil_12_write_start_control_vars_in[3] = arr__U1337_out[3];
assign op_hcompute_conv_stencil_12_write_start_control_vars_in[2] = arr__U1337_out[2];
assign op_hcompute_conv_stencil_12_write_start_control_vars_in[1] = arr__U1337_out[1];
assign op_hcompute_conv_stencil_12_write_start_control_vars_in[0] = arr__U1337_out[0];
op_hcompute_conv_stencil_12_write_start_control_vars_pt__U1224 op_hcompute_conv_stencil_12_write_start_control_vars (
    .in(op_hcompute_conv_stencil_12_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_12_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_13_clk = clk;
assign op_hcompute_conv_stencil_13_conv_stencil_op_hcompute_conv_stencil_13_read[0] = conv_stencil_op_hcompute_conv_stencil_13_read[0];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[7];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[6];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[5];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[4];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[3];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[2];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[1];
assign op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[0];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[7];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[6];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[5];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[4];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[3];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[2];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[1];
assign op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read[0];
cu_op_hcompute_conv_stencil_13 op_hcompute_conv_stencil_13 (
    .clk(op_hcompute_conv_stencil_13_clk),
    .conv_stencil_op_hcompute_conv_stencil_13_read(op_hcompute_conv_stencil_13_conv_stencil_op_hcompute_conv_stencil_13_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read(op_hcompute_conv_stencil_13_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_13_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read(op_hcompute_conv_stencil_13_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_13_read),
    .conv_stencil_op_hcompute_conv_stencil_13_write(op_hcompute_conv_stencil_13_conv_stencil_op_hcompute_conv_stencil_13_write)
);
assign op_hcompute_conv_stencil_13_exe_start_in = delay_reg__U1378_out;
op_hcompute_conv_stencil_13_exe_start_pt__U1376 op_hcompute_conv_stencil_13_exe_start (
    .in(op_hcompute_conv_stencil_13_exe_start_in),
    .out(op_hcompute_conv_stencil_13_exe_start_out)
);
assign op_hcompute_conv_stencil_13_exe_start_control_vars_in[4] = arr__U1387_out[4];
assign op_hcompute_conv_stencil_13_exe_start_control_vars_in[3] = arr__U1387_out[3];
assign op_hcompute_conv_stencil_13_exe_start_control_vars_in[2] = arr__U1387_out[2];
assign op_hcompute_conv_stencil_13_exe_start_control_vars_in[1] = arr__U1387_out[1];
assign op_hcompute_conv_stencil_13_exe_start_control_vars_in[0] = arr__U1387_out[0];
op_hcompute_conv_stencil_13_exe_start_control_vars_pt__U1379 op_hcompute_conv_stencil_13_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_13_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_13_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_13_port_controller_clk = clk;
affine_controller__U1344 op_hcompute_conv_stencil_13_port_controller (
    .clk(op_hcompute_conv_stencil_13_port_controller_clk),
    .valid(op_hcompute_conv_stencil_13_port_controller_valid),
    .d(op_hcompute_conv_stencil_13_port_controller_d)
);
assign op_hcompute_conv_stencil_13_read_start_in = op_hcompute_conv_stencil_13_port_controller_valid;
op_hcompute_conv_stencil_13_read_start_pt__U1374 op_hcompute_conv_stencil_13_read_start (
    .in(op_hcompute_conv_stencil_13_read_start_in),
    .out(op_hcompute_conv_stencil_13_read_start_out)
);
assign op_hcompute_conv_stencil_13_read_start_control_vars_in[4] = op_hcompute_conv_stencil_13_port_controller_d[4];
assign op_hcompute_conv_stencil_13_read_start_control_vars_in[3] = op_hcompute_conv_stencil_13_port_controller_d[3];
assign op_hcompute_conv_stencil_13_read_start_control_vars_in[2] = op_hcompute_conv_stencil_13_port_controller_d[2];
assign op_hcompute_conv_stencil_13_read_start_control_vars_in[1] = op_hcompute_conv_stencil_13_port_controller_d[1];
assign op_hcompute_conv_stencil_13_read_start_control_vars_in[0] = op_hcompute_conv_stencil_13_port_controller_d[0];
op_hcompute_conv_stencil_13_read_start_control_vars_pt__U1375 op_hcompute_conv_stencil_13_read_start_control_vars (
    .in(op_hcompute_conv_stencil_13_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_13_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_13_write_start_in = delay_reg__U1411_out;
op_hcompute_conv_stencil_13_write_start_pt__U1394 op_hcompute_conv_stencil_13_write_start (
    .in(op_hcompute_conv_stencil_13_write_start_in),
    .out(op_hcompute_conv_stencil_13_write_start_out)
);
assign op_hcompute_conv_stencil_13_write_start_control_vars_in[4] = arr__U1525_out[4];
assign op_hcompute_conv_stencil_13_write_start_control_vars_in[3] = arr__U1525_out[3];
assign op_hcompute_conv_stencil_13_write_start_control_vars_in[2] = arr__U1525_out[2];
assign op_hcompute_conv_stencil_13_write_start_control_vars_in[1] = arr__U1525_out[1];
assign op_hcompute_conv_stencil_13_write_start_control_vars_in[0] = arr__U1525_out[0];
op_hcompute_conv_stencil_13_write_start_control_vars_pt__U1412 op_hcompute_conv_stencil_13_write_start_control_vars (
    .in(op_hcompute_conv_stencil_13_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_13_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_14_clk = clk;
assign op_hcompute_conv_stencil_14_conv_stencil_op_hcompute_conv_stencil_14_read[0] = conv_stencil_op_hcompute_conv_stencil_14_read[0];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[7];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[6];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[5];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[4];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[3];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[2];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[1];
assign op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[0];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[7];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[6];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[5];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[4];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[3];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[2];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[1];
assign op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read[0];
cu_op_hcompute_conv_stencil_14 op_hcompute_conv_stencil_14 (
    .clk(op_hcompute_conv_stencil_14_clk),
    .conv_stencil_op_hcompute_conv_stencil_14_read(op_hcompute_conv_stencil_14_conv_stencil_op_hcompute_conv_stencil_14_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read(op_hcompute_conv_stencil_14_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_14_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read(op_hcompute_conv_stencil_14_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_14_read),
    .conv_stencil_op_hcompute_conv_stencil_14_write(op_hcompute_conv_stencil_14_conv_stencil_op_hcompute_conv_stencil_14_write)
);
assign op_hcompute_conv_stencil_14_exe_start_in = delay_reg__U1566_out;
op_hcompute_conv_stencil_14_exe_start_pt__U1564 op_hcompute_conv_stencil_14_exe_start (
    .in(op_hcompute_conv_stencil_14_exe_start_in),
    .out(op_hcompute_conv_stencil_14_exe_start_out)
);
assign op_hcompute_conv_stencil_14_exe_start_control_vars_in[4] = arr__U1575_out[4];
assign op_hcompute_conv_stencil_14_exe_start_control_vars_in[3] = arr__U1575_out[3];
assign op_hcompute_conv_stencil_14_exe_start_control_vars_in[2] = arr__U1575_out[2];
assign op_hcompute_conv_stencil_14_exe_start_control_vars_in[1] = arr__U1575_out[1];
assign op_hcompute_conv_stencil_14_exe_start_control_vars_in[0] = arr__U1575_out[0];
op_hcompute_conv_stencil_14_exe_start_control_vars_pt__U1567 op_hcompute_conv_stencil_14_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_14_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_14_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_14_port_controller_clk = clk;
affine_controller__U1532 op_hcompute_conv_stencil_14_port_controller (
    .clk(op_hcompute_conv_stencil_14_port_controller_clk),
    .valid(op_hcompute_conv_stencil_14_port_controller_valid),
    .d(op_hcompute_conv_stencil_14_port_controller_d)
);
assign op_hcompute_conv_stencil_14_read_start_in = op_hcompute_conv_stencil_14_port_controller_valid;
op_hcompute_conv_stencil_14_read_start_pt__U1562 op_hcompute_conv_stencil_14_read_start (
    .in(op_hcompute_conv_stencil_14_read_start_in),
    .out(op_hcompute_conv_stencil_14_read_start_out)
);
assign op_hcompute_conv_stencil_14_read_start_control_vars_in[4] = op_hcompute_conv_stencil_14_port_controller_d[4];
assign op_hcompute_conv_stencil_14_read_start_control_vars_in[3] = op_hcompute_conv_stencil_14_port_controller_d[3];
assign op_hcompute_conv_stencil_14_read_start_control_vars_in[2] = op_hcompute_conv_stencil_14_port_controller_d[2];
assign op_hcompute_conv_stencil_14_read_start_control_vars_in[1] = op_hcompute_conv_stencil_14_port_controller_d[1];
assign op_hcompute_conv_stencil_14_read_start_control_vars_in[0] = op_hcompute_conv_stencil_14_port_controller_d[0];
op_hcompute_conv_stencil_14_read_start_control_vars_pt__U1563 op_hcompute_conv_stencil_14_read_start_control_vars (
    .in(op_hcompute_conv_stencil_14_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_14_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_14_write_start_in = delay_reg__U1599_out;
op_hcompute_conv_stencil_14_write_start_pt__U1582 op_hcompute_conv_stencil_14_write_start (
    .in(op_hcompute_conv_stencil_14_write_start_in),
    .out(op_hcompute_conv_stencil_14_write_start_out)
);
assign op_hcompute_conv_stencil_14_write_start_control_vars_in[4] = arr__U1713_out[4];
assign op_hcompute_conv_stencil_14_write_start_control_vars_in[3] = arr__U1713_out[3];
assign op_hcompute_conv_stencil_14_write_start_control_vars_in[2] = arr__U1713_out[2];
assign op_hcompute_conv_stencil_14_write_start_control_vars_in[1] = arr__U1713_out[1];
assign op_hcompute_conv_stencil_14_write_start_control_vars_in[0] = arr__U1713_out[0];
op_hcompute_conv_stencil_14_write_start_control_vars_pt__U1600 op_hcompute_conv_stencil_14_write_start_control_vars (
    .in(op_hcompute_conv_stencil_14_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_14_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_15_clk = clk;
assign op_hcompute_conv_stencil_15_conv_stencil_op_hcompute_conv_stencil_15_read[0] = conv_stencil_op_hcompute_conv_stencil_15_read[0];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[7];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[6];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[5];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[4];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[3];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[2];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[1];
assign op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[0];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[7];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[6];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[5];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[4];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[3];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[2];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[1];
assign op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read[0];
cu_op_hcompute_conv_stencil_15 op_hcompute_conv_stencil_15 (
    .clk(op_hcompute_conv_stencil_15_clk),
    .conv_stencil_op_hcompute_conv_stencil_15_read(op_hcompute_conv_stencil_15_conv_stencil_op_hcompute_conv_stencil_15_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read(op_hcompute_conv_stencil_15_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_15_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read(op_hcompute_conv_stencil_15_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_15_read),
    .conv_stencil_op_hcompute_conv_stencil_15_write(op_hcompute_conv_stencil_15_conv_stencil_op_hcompute_conv_stencil_15_write)
);
assign op_hcompute_conv_stencil_15_exe_start_in = delay_reg__U1754_out;
op_hcompute_conv_stencil_15_exe_start_pt__U1752 op_hcompute_conv_stencil_15_exe_start (
    .in(op_hcompute_conv_stencil_15_exe_start_in),
    .out(op_hcompute_conv_stencil_15_exe_start_out)
);
assign op_hcompute_conv_stencil_15_exe_start_control_vars_in[4] = arr__U1763_out[4];
assign op_hcompute_conv_stencil_15_exe_start_control_vars_in[3] = arr__U1763_out[3];
assign op_hcompute_conv_stencil_15_exe_start_control_vars_in[2] = arr__U1763_out[2];
assign op_hcompute_conv_stencil_15_exe_start_control_vars_in[1] = arr__U1763_out[1];
assign op_hcompute_conv_stencil_15_exe_start_control_vars_in[0] = arr__U1763_out[0];
op_hcompute_conv_stencil_15_exe_start_control_vars_pt__U1755 op_hcompute_conv_stencil_15_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_15_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_15_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_15_port_controller_clk = clk;
affine_controller__U1720 op_hcompute_conv_stencil_15_port_controller (
    .clk(op_hcompute_conv_stencil_15_port_controller_clk),
    .valid(op_hcompute_conv_stencil_15_port_controller_valid),
    .d(op_hcompute_conv_stencil_15_port_controller_d)
);
assign op_hcompute_conv_stencil_15_read_start_in = op_hcompute_conv_stencil_15_port_controller_valid;
op_hcompute_conv_stencil_15_read_start_pt__U1750 op_hcompute_conv_stencil_15_read_start (
    .in(op_hcompute_conv_stencil_15_read_start_in),
    .out(op_hcompute_conv_stencil_15_read_start_out)
);
assign op_hcompute_conv_stencil_15_read_start_control_vars_in[4] = op_hcompute_conv_stencil_15_port_controller_d[4];
assign op_hcompute_conv_stencil_15_read_start_control_vars_in[3] = op_hcompute_conv_stencil_15_port_controller_d[3];
assign op_hcompute_conv_stencil_15_read_start_control_vars_in[2] = op_hcompute_conv_stencil_15_port_controller_d[2];
assign op_hcompute_conv_stencil_15_read_start_control_vars_in[1] = op_hcompute_conv_stencil_15_port_controller_d[1];
assign op_hcompute_conv_stencil_15_read_start_control_vars_in[0] = op_hcompute_conv_stencil_15_port_controller_d[0];
op_hcompute_conv_stencil_15_read_start_control_vars_pt__U1751 op_hcompute_conv_stencil_15_read_start_control_vars (
    .in(op_hcompute_conv_stencil_15_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_15_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_15_write_start_in = delay_reg__U1787_out;
op_hcompute_conv_stencil_15_write_start_pt__U1770 op_hcompute_conv_stencil_15_write_start (
    .in(op_hcompute_conv_stencil_15_write_start_in),
    .out(op_hcompute_conv_stencil_15_write_start_out)
);
assign op_hcompute_conv_stencil_15_write_start_control_vars_in[4] = arr__U1901_out[4];
assign op_hcompute_conv_stencil_15_write_start_control_vars_in[3] = arr__U1901_out[3];
assign op_hcompute_conv_stencil_15_write_start_control_vars_in[2] = arr__U1901_out[2];
assign op_hcompute_conv_stencil_15_write_start_control_vars_in[1] = arr__U1901_out[1];
assign op_hcompute_conv_stencil_15_write_start_control_vars_in[0] = arr__U1901_out[0];
op_hcompute_conv_stencil_15_write_start_control_vars_pt__U1788 op_hcompute_conv_stencil_15_write_start_control_vars (
    .in(op_hcompute_conv_stencil_15_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_15_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_exe_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_exe_start_pt__U262 op_hcompute_conv_stencil_1_exe_start (
    .in(op_hcompute_conv_stencil_1_exe_start_in),
    .out(op_hcompute_conv_stencil_1_exe_start_out)
);
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U263 op_hcompute_conv_stencil_1_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_1_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_port_controller_clk = clk;
affine_controller__U243 op_hcompute_conv_stencil_1_port_controller (
    .clk(op_hcompute_conv_stencil_1_port_controller_clk),
    .valid(op_hcompute_conv_stencil_1_port_controller_valid),
    .d(op_hcompute_conv_stencil_1_port_controller_d)
);
assign op_hcompute_conv_stencil_1_read_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_read_start_pt__U260 op_hcompute_conv_stencil_1_read_start (
    .in(op_hcompute_conv_stencil_1_read_start_in),
    .out(op_hcompute_conv_stencil_1_read_start_out)
);
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_read_start_control_vars_pt__U261 op_hcompute_conv_stencil_1_read_start_control_vars (
    .in(op_hcompute_conv_stencil_1_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_write_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_write_start_pt__U264 op_hcompute_conv_stencil_1_write_start (
    .in(op_hcompute_conv_stencil_1_write_start_in),
    .out(op_hcompute_conv_stencil_1_write_start_out)
);
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_write_start_control_vars_pt__U265 op_hcompute_conv_stencil_1_write_start_control_vars (
    .in(op_hcompute_conv_stencil_1_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_clk = clk;
cu_op_hcompute_conv_stencil_2 op_hcompute_conv_stencil_2 (
    .clk(op_hcompute_conv_stencil_2_clk),
    .conv_stencil_op_hcompute_conv_stencil_2_write(op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write)
);
assign op_hcompute_conv_stencil_2_exe_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_exe_start_pt__U285 op_hcompute_conv_stencil_2_exe_start (
    .in(op_hcompute_conv_stencil_2_exe_start_in),
    .out(op_hcompute_conv_stencil_2_exe_start_out)
);
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U286 op_hcompute_conv_stencil_2_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_2_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_port_controller_clk = clk;
affine_controller__U266 op_hcompute_conv_stencil_2_port_controller (
    .clk(op_hcompute_conv_stencil_2_port_controller_clk),
    .valid(op_hcompute_conv_stencil_2_port_controller_valid),
    .d(op_hcompute_conv_stencil_2_port_controller_d)
);
assign op_hcompute_conv_stencil_2_read_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_read_start_pt__U283 op_hcompute_conv_stencil_2_read_start (
    .in(op_hcompute_conv_stencil_2_read_start_in),
    .out(op_hcompute_conv_stencil_2_read_start_out)
);
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_read_start_control_vars_pt__U284 op_hcompute_conv_stencil_2_read_start_control_vars (
    .in(op_hcompute_conv_stencil_2_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_write_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_write_start_pt__U287 op_hcompute_conv_stencil_2_write_start (
    .in(op_hcompute_conv_stencil_2_write_start_in),
    .out(op_hcompute_conv_stencil_2_write_start_out)
);
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_write_start_control_vars_pt__U288 op_hcompute_conv_stencil_2_write_start_control_vars (
    .in(op_hcompute_conv_stencil_2_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_clk = clk;
cu_op_hcompute_conv_stencil_3 op_hcompute_conv_stencil_3 (
    .clk(op_hcompute_conv_stencil_3_clk),
    .conv_stencil_op_hcompute_conv_stencil_3_write(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write)
);
assign op_hcompute_conv_stencil_3_exe_start_in = op_hcompute_conv_stencil_3_port_controller_valid;
op_hcompute_conv_stencil_3_exe_start_pt__U308 op_hcompute_conv_stencil_3_exe_start (
    .in(op_hcompute_conv_stencil_3_exe_start_in),
    .out(op_hcompute_conv_stencil_3_exe_start_out)
);
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U309 op_hcompute_conv_stencil_3_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_3_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_port_controller_clk = clk;
affine_controller__U289 op_hcompute_conv_stencil_3_port_controller (
    .clk(op_hcompute_conv_stencil_3_port_controller_clk),
    .valid(op_hcompute_conv_stencil_3_port_controller_valid),
    .d(op_hcompute_conv_stencil_3_port_controller_d)
);
assign op_hcompute_conv_stencil_3_read_start_in = op_hcompute_conv_stencil_3_port_controller_valid;
op_hcompute_conv_stencil_3_read_start_pt__U306 op_hcompute_conv_stencil_3_read_start (
    .in(op_hcompute_conv_stencil_3_read_start_in),
    .out(op_hcompute_conv_stencil_3_read_start_out)
);
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
op_hcompute_conv_stencil_3_read_start_control_vars_pt__U307 op_hcompute_conv_stencil_3_read_start_control_vars (
    .in(op_hcompute_conv_stencil_3_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_write_start_in = op_hcompute_conv_stencil_3_port_controller_valid;
op_hcompute_conv_stencil_3_write_start_pt__U310 op_hcompute_conv_stencil_3_write_start (
    .in(op_hcompute_conv_stencil_3_write_start_in),
    .out(op_hcompute_conv_stencil_3_write_start_out)
);
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
op_hcompute_conv_stencil_3_write_start_control_vars_pt__U311 op_hcompute_conv_stencil_3_write_start_control_vars (
    .in(op_hcompute_conv_stencil_3_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_clk = clk;
cu_op_hcompute_conv_stencil_4 op_hcompute_conv_stencil_4 (
    .clk(op_hcompute_conv_stencil_4_clk),
    .conv_stencil_op_hcompute_conv_stencil_4_write(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write)
);
assign op_hcompute_conv_stencil_4_exe_start_in = op_hcompute_conv_stencil_4_port_controller_valid;
op_hcompute_conv_stencil_4_exe_start_pt__U331 op_hcompute_conv_stencil_4_exe_start (
    .in(op_hcompute_conv_stencil_4_exe_start_in),
    .out(op_hcompute_conv_stencil_4_exe_start_out)
);
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U332 op_hcompute_conv_stencil_4_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_4_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_port_controller_clk = clk;
affine_controller__U312 op_hcompute_conv_stencil_4_port_controller (
    .clk(op_hcompute_conv_stencil_4_port_controller_clk),
    .valid(op_hcompute_conv_stencil_4_port_controller_valid),
    .d(op_hcompute_conv_stencil_4_port_controller_d)
);
assign op_hcompute_conv_stencil_4_read_start_in = op_hcompute_conv_stencil_4_port_controller_valid;
op_hcompute_conv_stencil_4_read_start_pt__U329 op_hcompute_conv_stencil_4_read_start (
    .in(op_hcompute_conv_stencil_4_read_start_in),
    .out(op_hcompute_conv_stencil_4_read_start_out)
);
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
op_hcompute_conv_stencil_4_read_start_control_vars_pt__U330 op_hcompute_conv_stencil_4_read_start_control_vars (
    .in(op_hcompute_conv_stencil_4_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_write_start_in = op_hcompute_conv_stencil_4_port_controller_valid;
op_hcompute_conv_stencil_4_write_start_pt__U333 op_hcompute_conv_stencil_4_write_start (
    .in(op_hcompute_conv_stencil_4_write_start_in),
    .out(op_hcompute_conv_stencil_4_write_start_out)
);
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
op_hcompute_conv_stencil_4_write_start_control_vars_pt__U334 op_hcompute_conv_stencil_4_write_start_control_vars (
    .in(op_hcompute_conv_stencil_4_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_clk = clk;
cu_op_hcompute_conv_stencil_5 op_hcompute_conv_stencil_5 (
    .clk(op_hcompute_conv_stencil_5_clk),
    .conv_stencil_op_hcompute_conv_stencil_5_write(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write)
);
assign op_hcompute_conv_stencil_5_exe_start_in = op_hcompute_conv_stencil_5_port_controller_valid;
op_hcompute_conv_stencil_5_exe_start_pt__U354 op_hcompute_conv_stencil_5_exe_start (
    .in(op_hcompute_conv_stencil_5_exe_start_in),
    .out(op_hcompute_conv_stencil_5_exe_start_out)
);
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U355 op_hcompute_conv_stencil_5_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_5_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_port_controller_clk = clk;
affine_controller__U335 op_hcompute_conv_stencil_5_port_controller (
    .clk(op_hcompute_conv_stencil_5_port_controller_clk),
    .valid(op_hcompute_conv_stencil_5_port_controller_valid),
    .d(op_hcompute_conv_stencil_5_port_controller_d)
);
assign op_hcompute_conv_stencil_5_read_start_in = op_hcompute_conv_stencil_5_port_controller_valid;
op_hcompute_conv_stencil_5_read_start_pt__U352 op_hcompute_conv_stencil_5_read_start (
    .in(op_hcompute_conv_stencil_5_read_start_in),
    .out(op_hcompute_conv_stencil_5_read_start_out)
);
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
op_hcompute_conv_stencil_5_read_start_control_vars_pt__U353 op_hcompute_conv_stencil_5_read_start_control_vars (
    .in(op_hcompute_conv_stencil_5_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_write_start_in = op_hcompute_conv_stencil_5_port_controller_valid;
op_hcompute_conv_stencil_5_write_start_pt__U356 op_hcompute_conv_stencil_5_write_start (
    .in(op_hcompute_conv_stencil_5_write_start_in),
    .out(op_hcompute_conv_stencil_5_write_start_out)
);
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
op_hcompute_conv_stencil_5_write_start_control_vars_pt__U357 op_hcompute_conv_stencil_5_write_start_control_vars (
    .in(op_hcompute_conv_stencil_5_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_6_clk = clk;
cu_op_hcompute_conv_stencil_6 op_hcompute_conv_stencil_6 (
    .clk(op_hcompute_conv_stencil_6_clk),
    .conv_stencil_op_hcompute_conv_stencil_6_write(op_hcompute_conv_stencil_6_conv_stencil_op_hcompute_conv_stencil_6_write)
);
assign op_hcompute_conv_stencil_6_exe_start_in = op_hcompute_conv_stencil_6_port_controller_valid;
op_hcompute_conv_stencil_6_exe_start_pt__U377 op_hcompute_conv_stencil_6_exe_start (
    .in(op_hcompute_conv_stencil_6_exe_start_in),
    .out(op_hcompute_conv_stencil_6_exe_start_out)
);
assign op_hcompute_conv_stencil_6_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_6_port_controller_d[2];
assign op_hcompute_conv_stencil_6_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_6_port_controller_d[1];
assign op_hcompute_conv_stencil_6_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_6_port_controller_d[0];
op_hcompute_conv_stencil_6_exe_start_control_vars_pt__U378 op_hcompute_conv_stencil_6_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_6_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_6_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_6_port_controller_clk = clk;
affine_controller__U358 op_hcompute_conv_stencil_6_port_controller (
    .clk(op_hcompute_conv_stencil_6_port_controller_clk),
    .valid(op_hcompute_conv_stencil_6_port_controller_valid),
    .d(op_hcompute_conv_stencil_6_port_controller_d)
);
assign op_hcompute_conv_stencil_6_read_start_in = op_hcompute_conv_stencil_6_port_controller_valid;
op_hcompute_conv_stencil_6_read_start_pt__U375 op_hcompute_conv_stencil_6_read_start (
    .in(op_hcompute_conv_stencil_6_read_start_in),
    .out(op_hcompute_conv_stencil_6_read_start_out)
);
assign op_hcompute_conv_stencil_6_read_start_control_vars_in[2] = op_hcompute_conv_stencil_6_port_controller_d[2];
assign op_hcompute_conv_stencil_6_read_start_control_vars_in[1] = op_hcompute_conv_stencil_6_port_controller_d[1];
assign op_hcompute_conv_stencil_6_read_start_control_vars_in[0] = op_hcompute_conv_stencil_6_port_controller_d[0];
op_hcompute_conv_stencil_6_read_start_control_vars_pt__U376 op_hcompute_conv_stencil_6_read_start_control_vars (
    .in(op_hcompute_conv_stencil_6_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_6_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_6_write_start_in = op_hcompute_conv_stencil_6_port_controller_valid;
op_hcompute_conv_stencil_6_write_start_pt__U379 op_hcompute_conv_stencil_6_write_start (
    .in(op_hcompute_conv_stencil_6_write_start_in),
    .out(op_hcompute_conv_stencil_6_write_start_out)
);
assign op_hcompute_conv_stencil_6_write_start_control_vars_in[2] = op_hcompute_conv_stencil_6_port_controller_d[2];
assign op_hcompute_conv_stencil_6_write_start_control_vars_in[1] = op_hcompute_conv_stencil_6_port_controller_d[1];
assign op_hcompute_conv_stencil_6_write_start_control_vars_in[0] = op_hcompute_conv_stencil_6_port_controller_d[0];
op_hcompute_conv_stencil_6_write_start_control_vars_pt__U380 op_hcompute_conv_stencil_6_write_start_control_vars (
    .in(op_hcompute_conv_stencil_6_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_6_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_7_clk = clk;
cu_op_hcompute_conv_stencil_7 op_hcompute_conv_stencil_7 (
    .clk(op_hcompute_conv_stencil_7_clk),
    .conv_stencil_op_hcompute_conv_stencil_7_write(op_hcompute_conv_stencil_7_conv_stencil_op_hcompute_conv_stencil_7_write)
);
assign op_hcompute_conv_stencil_7_exe_start_in = op_hcompute_conv_stencil_7_port_controller_valid;
op_hcompute_conv_stencil_7_exe_start_pt__U400 op_hcompute_conv_stencil_7_exe_start (
    .in(op_hcompute_conv_stencil_7_exe_start_in),
    .out(op_hcompute_conv_stencil_7_exe_start_out)
);
assign op_hcompute_conv_stencil_7_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_7_port_controller_d[2];
assign op_hcompute_conv_stencil_7_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_7_port_controller_d[1];
assign op_hcompute_conv_stencil_7_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_7_port_controller_d[0];
op_hcompute_conv_stencil_7_exe_start_control_vars_pt__U401 op_hcompute_conv_stencil_7_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_7_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_7_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_7_port_controller_clk = clk;
affine_controller__U381 op_hcompute_conv_stencil_7_port_controller (
    .clk(op_hcompute_conv_stencil_7_port_controller_clk),
    .valid(op_hcompute_conv_stencil_7_port_controller_valid),
    .d(op_hcompute_conv_stencil_7_port_controller_d)
);
assign op_hcompute_conv_stencil_7_read_start_in = op_hcompute_conv_stencil_7_port_controller_valid;
op_hcompute_conv_stencil_7_read_start_pt__U398 op_hcompute_conv_stencil_7_read_start (
    .in(op_hcompute_conv_stencil_7_read_start_in),
    .out(op_hcompute_conv_stencil_7_read_start_out)
);
assign op_hcompute_conv_stencil_7_read_start_control_vars_in[2] = op_hcompute_conv_stencil_7_port_controller_d[2];
assign op_hcompute_conv_stencil_7_read_start_control_vars_in[1] = op_hcompute_conv_stencil_7_port_controller_d[1];
assign op_hcompute_conv_stencil_7_read_start_control_vars_in[0] = op_hcompute_conv_stencil_7_port_controller_d[0];
op_hcompute_conv_stencil_7_read_start_control_vars_pt__U399 op_hcompute_conv_stencil_7_read_start_control_vars (
    .in(op_hcompute_conv_stencil_7_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_7_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_7_write_start_in = op_hcompute_conv_stencil_7_port_controller_valid;
op_hcompute_conv_stencil_7_write_start_pt__U402 op_hcompute_conv_stencil_7_write_start (
    .in(op_hcompute_conv_stencil_7_write_start_in),
    .out(op_hcompute_conv_stencil_7_write_start_out)
);
assign op_hcompute_conv_stencil_7_write_start_control_vars_in[2] = op_hcompute_conv_stencil_7_port_controller_d[2];
assign op_hcompute_conv_stencil_7_write_start_control_vars_in[1] = op_hcompute_conv_stencil_7_port_controller_d[1];
assign op_hcompute_conv_stencil_7_write_start_control_vars_in[0] = op_hcompute_conv_stencil_7_port_controller_d[0];
op_hcompute_conv_stencil_7_write_start_control_vars_pt__U403 op_hcompute_conv_stencil_7_write_start_control_vars (
    .in(op_hcompute_conv_stencil_7_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_7_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_8_clk = clk;
assign op_hcompute_conv_stencil_8_conv_stencil_op_hcompute_conv_stencil_8_read[0] = conv_stencil_op_hcompute_conv_stencil_8_read[0];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[7];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[6];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[5];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[4];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[3];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[2];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[1];
assign op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[0];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[7];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[6];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[5];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[4];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[3];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[2];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[1];
assign op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read[0];
cu_op_hcompute_conv_stencil_8 op_hcompute_conv_stencil_8 (
    .clk(op_hcompute_conv_stencil_8_clk),
    .conv_stencil_op_hcompute_conv_stencil_8_read(op_hcompute_conv_stencil_8_conv_stencil_op_hcompute_conv_stencil_8_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read(op_hcompute_conv_stencil_8_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_8_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read(op_hcompute_conv_stencil_8_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_8_read),
    .conv_stencil_op_hcompute_conv_stencil_8_write(op_hcompute_conv_stencil_8_conv_stencil_op_hcompute_conv_stencil_8_write)
);
assign op_hcompute_conv_stencil_8_exe_start_in = delay_reg__U438_out;
op_hcompute_conv_stencil_8_exe_start_pt__U436 op_hcompute_conv_stencil_8_exe_start (
    .in(op_hcompute_conv_stencil_8_exe_start_in),
    .out(op_hcompute_conv_stencil_8_exe_start_out)
);
assign op_hcompute_conv_stencil_8_exe_start_control_vars_in[4] = arr__U447_out[4];
assign op_hcompute_conv_stencil_8_exe_start_control_vars_in[3] = arr__U447_out[3];
assign op_hcompute_conv_stencil_8_exe_start_control_vars_in[2] = arr__U447_out[2];
assign op_hcompute_conv_stencil_8_exe_start_control_vars_in[1] = arr__U447_out[1];
assign op_hcompute_conv_stencil_8_exe_start_control_vars_in[0] = arr__U447_out[0];
op_hcompute_conv_stencil_8_exe_start_control_vars_pt__U439 op_hcompute_conv_stencil_8_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_8_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_8_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_8_port_controller_clk = clk;
affine_controller__U404 op_hcompute_conv_stencil_8_port_controller (
    .clk(op_hcompute_conv_stencil_8_port_controller_clk),
    .valid(op_hcompute_conv_stencil_8_port_controller_valid),
    .d(op_hcompute_conv_stencil_8_port_controller_d)
);
assign op_hcompute_conv_stencil_8_read_start_in = op_hcompute_conv_stencil_8_port_controller_valid;
op_hcompute_conv_stencil_8_read_start_pt__U434 op_hcompute_conv_stencil_8_read_start (
    .in(op_hcompute_conv_stencil_8_read_start_in),
    .out(op_hcompute_conv_stencil_8_read_start_out)
);
assign op_hcompute_conv_stencil_8_read_start_control_vars_in[4] = op_hcompute_conv_stencil_8_port_controller_d[4];
assign op_hcompute_conv_stencil_8_read_start_control_vars_in[3] = op_hcompute_conv_stencil_8_port_controller_d[3];
assign op_hcompute_conv_stencil_8_read_start_control_vars_in[2] = op_hcompute_conv_stencil_8_port_controller_d[2];
assign op_hcompute_conv_stencil_8_read_start_control_vars_in[1] = op_hcompute_conv_stencil_8_port_controller_d[1];
assign op_hcompute_conv_stencil_8_read_start_control_vars_in[0] = op_hcompute_conv_stencil_8_port_controller_d[0];
op_hcompute_conv_stencil_8_read_start_control_vars_pt__U435 op_hcompute_conv_stencil_8_read_start_control_vars (
    .in(op_hcompute_conv_stencil_8_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_8_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_8_write_start_in = delay_reg__U471_out;
op_hcompute_conv_stencil_8_write_start_pt__U454 op_hcompute_conv_stencil_8_write_start (
    .in(op_hcompute_conv_stencil_8_write_start_in),
    .out(op_hcompute_conv_stencil_8_write_start_out)
);
assign op_hcompute_conv_stencil_8_write_start_control_vars_in[4] = arr__U585_out[4];
assign op_hcompute_conv_stencil_8_write_start_control_vars_in[3] = arr__U585_out[3];
assign op_hcompute_conv_stencil_8_write_start_control_vars_in[2] = arr__U585_out[2];
assign op_hcompute_conv_stencil_8_write_start_control_vars_in[1] = arr__U585_out[1];
assign op_hcompute_conv_stencil_8_write_start_control_vars_in[0] = arr__U585_out[0];
op_hcompute_conv_stencil_8_write_start_control_vars_pt__U472 op_hcompute_conv_stencil_8_write_start_control_vars (
    .in(op_hcompute_conv_stencil_8_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_8_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_9_clk = clk;
assign op_hcompute_conv_stencil_9_conv_stencil_op_hcompute_conv_stencil_9_read[0] = conv_stencil_op_hcompute_conv_stencil_9_read[0];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[7];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[6];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[5];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[4];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[3];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[2];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[1];
assign op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[0];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[7];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[6];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[5];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[4];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[3];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[2];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[1];
assign op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read[0];
cu_op_hcompute_conv_stencil_9 op_hcompute_conv_stencil_9 (
    .clk(op_hcompute_conv_stencil_9_clk),
    .conv_stencil_op_hcompute_conv_stencil_9_read(op_hcompute_conv_stencil_9_conv_stencil_op_hcompute_conv_stencil_9_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read(op_hcompute_conv_stencil_9_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_9_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read(op_hcompute_conv_stencil_9_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_9_read),
    .conv_stencil_op_hcompute_conv_stencil_9_write(op_hcompute_conv_stencil_9_conv_stencil_op_hcompute_conv_stencil_9_write)
);
assign op_hcompute_conv_stencil_9_exe_start_in = delay_reg__U626_out;
op_hcompute_conv_stencil_9_exe_start_pt__U624 op_hcompute_conv_stencil_9_exe_start (
    .in(op_hcompute_conv_stencil_9_exe_start_in),
    .out(op_hcompute_conv_stencil_9_exe_start_out)
);
assign op_hcompute_conv_stencil_9_exe_start_control_vars_in[4] = arr__U635_out[4];
assign op_hcompute_conv_stencil_9_exe_start_control_vars_in[3] = arr__U635_out[3];
assign op_hcompute_conv_stencil_9_exe_start_control_vars_in[2] = arr__U635_out[2];
assign op_hcompute_conv_stencil_9_exe_start_control_vars_in[1] = arr__U635_out[1];
assign op_hcompute_conv_stencil_9_exe_start_control_vars_in[0] = arr__U635_out[0];
op_hcompute_conv_stencil_9_exe_start_control_vars_pt__U627 op_hcompute_conv_stencil_9_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_9_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_9_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_9_port_controller_clk = clk;
affine_controller__U592 op_hcompute_conv_stencil_9_port_controller (
    .clk(op_hcompute_conv_stencil_9_port_controller_clk),
    .valid(op_hcompute_conv_stencil_9_port_controller_valid),
    .d(op_hcompute_conv_stencil_9_port_controller_d)
);
assign op_hcompute_conv_stencil_9_read_start_in = op_hcompute_conv_stencil_9_port_controller_valid;
op_hcompute_conv_stencil_9_read_start_pt__U622 op_hcompute_conv_stencil_9_read_start (
    .in(op_hcompute_conv_stencil_9_read_start_in),
    .out(op_hcompute_conv_stencil_9_read_start_out)
);
assign op_hcompute_conv_stencil_9_read_start_control_vars_in[4] = op_hcompute_conv_stencil_9_port_controller_d[4];
assign op_hcompute_conv_stencil_9_read_start_control_vars_in[3] = op_hcompute_conv_stencil_9_port_controller_d[3];
assign op_hcompute_conv_stencil_9_read_start_control_vars_in[2] = op_hcompute_conv_stencil_9_port_controller_d[2];
assign op_hcompute_conv_stencil_9_read_start_control_vars_in[1] = op_hcompute_conv_stencil_9_port_controller_d[1];
assign op_hcompute_conv_stencil_9_read_start_control_vars_in[0] = op_hcompute_conv_stencil_9_port_controller_d[0];
op_hcompute_conv_stencil_9_read_start_control_vars_pt__U623 op_hcompute_conv_stencil_9_read_start_control_vars (
    .in(op_hcompute_conv_stencil_9_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_9_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_9_write_start_in = delay_reg__U659_out;
op_hcompute_conv_stencil_9_write_start_pt__U642 op_hcompute_conv_stencil_9_write_start (
    .in(op_hcompute_conv_stencil_9_write_start_in),
    .out(op_hcompute_conv_stencil_9_write_start_out)
);
assign op_hcompute_conv_stencil_9_write_start_control_vars_in[4] = arr__U773_out[4];
assign op_hcompute_conv_stencil_9_write_start_control_vars_in[3] = arr__U773_out[3];
assign op_hcompute_conv_stencil_9_write_start_control_vars_in[2] = arr__U773_out[2];
assign op_hcompute_conv_stencil_9_write_start_control_vars_in[1] = arr__U773_out[1];
assign op_hcompute_conv_stencil_9_write_start_control_vars_in[0] = arr__U773_out[0];
op_hcompute_conv_stencil_9_write_start_control_vars_pt__U660 op_hcompute_conv_stencil_9_write_start_control_vars (
    .in(op_hcompute_conv_stencil_9_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_9_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_exe_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_exe_start_pt__U239 op_hcompute_conv_stencil_exe_start (
    .in(op_hcompute_conv_stencil_exe_start_in),
    .out(op_hcompute_conv_stencil_exe_start_out)
);
assign op_hcompute_conv_stencil_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_exe_start_control_vars_pt__U240 op_hcompute_conv_stencil_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_port_controller_clk = clk;
affine_controller__U220 op_hcompute_conv_stencil_port_controller (
    .clk(op_hcompute_conv_stencil_port_controller_clk),
    .valid(op_hcompute_conv_stencil_port_controller_valid),
    .d(op_hcompute_conv_stencil_port_controller_d)
);
assign op_hcompute_conv_stencil_read_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_read_start_pt__U237 op_hcompute_conv_stencil_read_start (
    .in(op_hcompute_conv_stencil_read_start_in),
    .out(op_hcompute_conv_stencil_read_start_out)
);
assign op_hcompute_conv_stencil_read_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_read_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_read_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_read_start_control_vars_pt__U238 op_hcompute_conv_stencil_read_start_control_vars (
    .in(op_hcompute_conv_stencil_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_write_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_write_start_pt__U241 op_hcompute_conv_stencil_write_start (
    .in(op_hcompute_conv_stencil_write_start_in),
    .out(op_hcompute_conv_stencil_write_start_out)
);
assign op_hcompute_conv_stencil_write_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_write_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_write_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_write_start_control_vars_pt__U242 op_hcompute_conv_stencil_write_start_control_vars (
    .in(op_hcompute_conv_stencil_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read[0] = hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil op_hcompute_hw_input_global_wrapper_stencil (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_clk),
    .hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read(op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write(op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
assign op_hcompute_hw_input_global_wrapper_stencil_1_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_1_hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read[0] = hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil_1 op_hcompute_hw_input_global_wrapper_stencil_1 (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_1_clk),
    .hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read(op_hcompute_hw_input_global_wrapper_stencil_1_hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write(op_hcompute_hw_input_global_wrapper_stencil_1_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_1_write)
);
assign op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_in = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_pt__U42 op_hcompute_hw_input_global_wrapper_stencil_1_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_pt__U43 op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_1_exe_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_clk = clk;
affine_controller__U23 op_hcompute_hw_input_global_wrapper_stencil_1_port_controller (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d)
);
assign op_hcompute_hw_input_global_wrapper_stencil_1_read_start_in = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_1_read_start_pt__U40 op_hcompute_hw_input_global_wrapper_stencil_1_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_1_read_start_in),
    .out(hw_input_stencil_clkwrk_1_op_hcompute_hw_input_global_wrapper_stencil_1_read_en)
);
assign op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_pt__U41 op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_1_read_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_1_write_start_in = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_1_write_start_pt__U44 op_hcompute_hw_input_global_wrapper_stencil_1_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_1_write_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_1_write_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_1_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_pt__U45 op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_1_write_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_2_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_2_hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read[0] = hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil_2 op_hcompute_hw_input_global_wrapper_stencil_2 (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_2_clk),
    .hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read(op_hcompute_hw_input_global_wrapper_stencil_2_hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write(op_hcompute_hw_input_global_wrapper_stencil_2_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_2_write)
);
assign op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_in = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_pt__U65 op_hcompute_hw_input_global_wrapper_stencil_2_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_pt__U66 op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_2_exe_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_clk = clk;
affine_controller__U46 op_hcompute_hw_input_global_wrapper_stencil_2_port_controller (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d)
);
assign op_hcompute_hw_input_global_wrapper_stencil_2_read_start_in = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_2_read_start_pt__U63 op_hcompute_hw_input_global_wrapper_stencil_2_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_2_read_start_in),
    .out(hw_input_stencil_clkwrk_2_op_hcompute_hw_input_global_wrapper_stencil_2_read_en)
);
assign op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_pt__U64 op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_2_read_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_2_write_start_in = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_2_write_start_pt__U67 op_hcompute_hw_input_global_wrapper_stencil_2_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_2_write_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_2_write_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_2_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_pt__U68 op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_2_write_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_3_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_3_hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read[0] = hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil_3 op_hcompute_hw_input_global_wrapper_stencil_3 (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_3_clk),
    .hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read(op_hcompute_hw_input_global_wrapper_stencil_3_hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write(op_hcompute_hw_input_global_wrapper_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_3_write)
);
assign op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_in = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_pt__U88 op_hcompute_hw_input_global_wrapper_stencil_3_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_pt__U89 op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_3_exe_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_clk = clk;
affine_controller__U69 op_hcompute_hw_input_global_wrapper_stencil_3_port_controller (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d)
);
assign op_hcompute_hw_input_global_wrapper_stencil_3_read_start_in = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_3_read_start_pt__U86 op_hcompute_hw_input_global_wrapper_stencil_3_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_3_read_start_in),
    .out(hw_input_stencil_clkwrk_3_op_hcompute_hw_input_global_wrapper_stencil_3_read_en)
);
assign op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_pt__U87 op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_3_read_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_3_write_start_in = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_3_write_start_pt__U90 op_hcompute_hw_input_global_wrapper_stencil_3_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_3_write_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_3_write_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_3_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_pt__U91 op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_3_write_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_4_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_4_hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read[0] = hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil_4 op_hcompute_hw_input_global_wrapper_stencil_4 (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_4_clk),
    .hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read(op_hcompute_hw_input_global_wrapper_stencil_4_hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write(op_hcompute_hw_input_global_wrapper_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_4_write)
);
assign op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_in = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_pt__U111 op_hcompute_hw_input_global_wrapper_stencil_4_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_pt__U112 op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_4_exe_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_clk = clk;
affine_controller__U92 op_hcompute_hw_input_global_wrapper_stencil_4_port_controller (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d)
);
assign op_hcompute_hw_input_global_wrapper_stencil_4_read_start_in = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_4_read_start_pt__U109 op_hcompute_hw_input_global_wrapper_stencil_4_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_4_read_start_in),
    .out(hw_input_stencil_clkwrk_4_op_hcompute_hw_input_global_wrapper_stencil_4_read_en)
);
assign op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_pt__U110 op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_4_read_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_4_write_start_in = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_4_write_start_pt__U113 op_hcompute_hw_input_global_wrapper_stencil_4_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_4_write_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_4_write_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_4_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_pt__U114 op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_4_write_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_5_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_5_hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read[0] = hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil_5 op_hcompute_hw_input_global_wrapper_stencil_5 (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_5_clk),
    .hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read(op_hcompute_hw_input_global_wrapper_stencil_5_hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write(op_hcompute_hw_input_global_wrapper_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_5_write)
);
assign op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_in = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_pt__U134 op_hcompute_hw_input_global_wrapper_stencil_5_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_pt__U135 op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_5_exe_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_clk = clk;
affine_controller__U115 op_hcompute_hw_input_global_wrapper_stencil_5_port_controller (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d)
);
assign op_hcompute_hw_input_global_wrapper_stencil_5_read_start_in = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_5_read_start_pt__U132 op_hcompute_hw_input_global_wrapper_stencil_5_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_5_read_start_in),
    .out(hw_input_stencil_clkwrk_5_op_hcompute_hw_input_global_wrapper_stencil_5_read_en)
);
assign op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_pt__U133 op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_5_read_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_5_write_start_in = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_5_write_start_pt__U136 op_hcompute_hw_input_global_wrapper_stencil_5_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_5_write_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_5_write_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_5_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_pt__U137 op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_5_write_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_6_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_6_hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read[0] = hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil_6 op_hcompute_hw_input_global_wrapper_stencil_6 (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_6_clk),
    .hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read(op_hcompute_hw_input_global_wrapper_stencil_6_hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write(op_hcompute_hw_input_global_wrapper_stencil_6_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_6_write)
);
assign op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_in = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_pt__U157 op_hcompute_hw_input_global_wrapper_stencil_6_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_pt__U158 op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_6_exe_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_clk = clk;
affine_controller__U138 op_hcompute_hw_input_global_wrapper_stencil_6_port_controller (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d)
);
assign op_hcompute_hw_input_global_wrapper_stencil_6_read_start_in = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_6_read_start_pt__U155 op_hcompute_hw_input_global_wrapper_stencil_6_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_6_read_start_in),
    .out(hw_input_stencil_clkwrk_6_op_hcompute_hw_input_global_wrapper_stencil_6_read_en)
);
assign op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_pt__U156 op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_6_read_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_6_write_start_in = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_6_write_start_pt__U159 op_hcompute_hw_input_global_wrapper_stencil_6_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_6_write_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_6_write_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_6_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_pt__U160 op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_6_write_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_7_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_7_hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read[0] = hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil_7 op_hcompute_hw_input_global_wrapper_stencil_7 (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_7_clk),
    .hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read(op_hcompute_hw_input_global_wrapper_stencil_7_hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write(op_hcompute_hw_input_global_wrapper_stencil_7_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_7_write)
);
assign op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_in = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_pt__U180 op_hcompute_hw_input_global_wrapper_stencil_7_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_pt__U181 op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_7_exe_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_clk = clk;
affine_controller__U161 op_hcompute_hw_input_global_wrapper_stencil_7_port_controller (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d)
);
assign op_hcompute_hw_input_global_wrapper_stencil_7_read_start_in = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_7_read_start_pt__U178 op_hcompute_hw_input_global_wrapper_stencil_7_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_7_read_start_in),
    .out(hw_input_stencil_clkwrk_7_op_hcompute_hw_input_global_wrapper_stencil_7_read_en)
);
assign op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_pt__U179 op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_7_read_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_7_write_start_in = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_7_write_start_pt__U182 op_hcompute_hw_input_global_wrapper_stencil_7_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_7_write_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_7_write_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_7_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_pt__U183 op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_7_write_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U19 op_hcompute_hw_input_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U20 op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk = clk;
affine_controller__U0 op_hcompute_hw_input_global_wrapper_stencil_port_controller (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_port_controller_d)
);
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U17 op_hcompute_hw_input_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_in),
    .out(hw_input_stencil_clkwrk_0_op_hcompute_hw_input_global_wrapper_stencil_read_en)
);
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U18 op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U21 op_hcompute_hw_input_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U22 op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_clk = clk;
assign op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_kernel_global_wrapper_stencil op_hcompute_hw_kernel_global_wrapper_stencil (
    .clk(op_hcompute_hw_kernel_global_wrapper_stencil_clk),
    .hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U216 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U217 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk = clk;
affine_controller__U184 op_hcompute_hw_kernel_global_wrapper_stencil_port_controller (
    .clk(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk),
    .valid(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U214 op_hcompute_hw_kernel_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in),
    .out(hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U215 op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U218 op_hcompute_hw_kernel_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U219 op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_clk = clk;
assign op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
cu_op_hcompute_hw_output_stencil op_hcompute_hw_output_stencil (
    .clk(op_hcompute_hw_output_stencil_clk),
    .conv_stencil_op_hcompute_hw_output_stencil_read(op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read),
    .hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write(op_hcompute_hw_output_stencil_hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write)
);
assign op_hcompute_hw_output_stencil_1_clk = clk;
assign op_hcompute_hw_output_stencil_1_conv_stencil_op_hcompute_hw_output_stencil_1_read[0] = conv_stencil_op_hcompute_hw_output_stencil_1_read[0];
cu_op_hcompute_hw_output_stencil_1 op_hcompute_hw_output_stencil_1 (
    .clk(op_hcompute_hw_output_stencil_1_clk),
    .conv_stencil_op_hcompute_hw_output_stencil_1_read(op_hcompute_hw_output_stencil_1_conv_stencil_op_hcompute_hw_output_stencil_1_read),
    .hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write(op_hcompute_hw_output_stencil_1_hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write)
);
assign op_hcompute_hw_output_stencil_1_exe_start_in = delay_reg__U1976_out;
op_hcompute_hw_output_stencil_1_exe_start_pt__U1974 op_hcompute_hw_output_stencil_1_exe_start (
    .in(op_hcompute_hw_output_stencil_1_exe_start_in),
    .out(op_hcompute_hw_output_stencil_1_exe_start_out)
);
assign op_hcompute_hw_output_stencil_1_exe_start_control_vars_in[2] = arr__U1983_out[2];
assign op_hcompute_hw_output_stencil_1_exe_start_control_vars_in[1] = arr__U1983_out[1];
assign op_hcompute_hw_output_stencil_1_exe_start_control_vars_in[0] = arr__U1983_out[0];
op_hcompute_hw_output_stencil_1_exe_start_control_vars_pt__U1977 op_hcompute_hw_output_stencil_1_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_1_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_1_exe_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_1_port_controller_clk = clk;
affine_controller__U1955 op_hcompute_hw_output_stencil_1_port_controller (
    .clk(op_hcompute_hw_output_stencil_1_port_controller_clk),
    .valid(op_hcompute_hw_output_stencil_1_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_1_port_controller_d)
);
assign op_hcompute_hw_output_stencil_1_read_start_in = op_hcompute_hw_output_stencil_1_port_controller_valid;
op_hcompute_hw_output_stencil_1_read_start_pt__U1972 op_hcompute_hw_output_stencil_1_read_start (
    .in(op_hcompute_hw_output_stencil_1_read_start_in),
    .out(op_hcompute_hw_output_stencil_1_read_start_out)
);
assign op_hcompute_hw_output_stencil_1_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_1_port_controller_d[2];
assign op_hcompute_hw_output_stencil_1_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_1_port_controller_d[1];
assign op_hcompute_hw_output_stencil_1_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_1_port_controller_d[0];
op_hcompute_hw_output_stencil_1_read_start_control_vars_pt__U1973 op_hcompute_hw_output_stencil_1_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_1_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_1_read_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_1_write_start_in = delay_reg__U1990_out;
op_hcompute_hw_output_stencil_1_write_start_pt__U1988 op_hcompute_hw_output_stencil_1_write_start (
    .in(op_hcompute_hw_output_stencil_1_write_start_in),
    .out(hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write_valid)
);
assign op_hcompute_hw_output_stencil_1_write_start_control_vars_in[2] = arr__U1997_out[2];
assign op_hcompute_hw_output_stencil_1_write_start_control_vars_in[1] = arr__U1997_out[1];
assign op_hcompute_hw_output_stencil_1_write_start_control_vars_in[0] = arr__U1997_out[0];
op_hcompute_hw_output_stencil_1_write_start_control_vars_pt__U1991 op_hcompute_hw_output_stencil_1_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_1_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_1_write_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_2_clk = clk;
assign op_hcompute_hw_output_stencil_2_conv_stencil_op_hcompute_hw_output_stencil_2_read[0] = conv_stencil_op_hcompute_hw_output_stencil_2_read[0];
cu_op_hcompute_hw_output_stencil_2 op_hcompute_hw_output_stencil_2 (
    .clk(op_hcompute_hw_output_stencil_2_clk),
    .conv_stencil_op_hcompute_hw_output_stencil_2_read(op_hcompute_hw_output_stencil_2_conv_stencil_op_hcompute_hw_output_stencil_2_read),
    .hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write(op_hcompute_hw_output_stencil_2_hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write)
);
assign op_hcompute_hw_output_stencil_2_exe_start_in = delay_reg__U2023_out;
op_hcompute_hw_output_stencil_2_exe_start_pt__U2021 op_hcompute_hw_output_stencil_2_exe_start (
    .in(op_hcompute_hw_output_stencil_2_exe_start_in),
    .out(op_hcompute_hw_output_stencil_2_exe_start_out)
);
assign op_hcompute_hw_output_stencil_2_exe_start_control_vars_in[2] = arr__U2030_out[2];
assign op_hcompute_hw_output_stencil_2_exe_start_control_vars_in[1] = arr__U2030_out[1];
assign op_hcompute_hw_output_stencil_2_exe_start_control_vars_in[0] = arr__U2030_out[0];
op_hcompute_hw_output_stencil_2_exe_start_control_vars_pt__U2024 op_hcompute_hw_output_stencil_2_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_2_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_2_exe_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_2_port_controller_clk = clk;
affine_controller__U2002 op_hcompute_hw_output_stencil_2_port_controller (
    .clk(op_hcompute_hw_output_stencil_2_port_controller_clk),
    .valid(op_hcompute_hw_output_stencil_2_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_2_port_controller_d)
);
assign op_hcompute_hw_output_stencil_2_read_start_in = op_hcompute_hw_output_stencil_2_port_controller_valid;
op_hcompute_hw_output_stencil_2_read_start_pt__U2019 op_hcompute_hw_output_stencil_2_read_start (
    .in(op_hcompute_hw_output_stencil_2_read_start_in),
    .out(op_hcompute_hw_output_stencil_2_read_start_out)
);
assign op_hcompute_hw_output_stencil_2_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_2_port_controller_d[2];
assign op_hcompute_hw_output_stencil_2_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_2_port_controller_d[1];
assign op_hcompute_hw_output_stencil_2_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_2_port_controller_d[0];
op_hcompute_hw_output_stencil_2_read_start_control_vars_pt__U2020 op_hcompute_hw_output_stencil_2_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_2_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_2_read_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_2_write_start_in = delay_reg__U2037_out;
op_hcompute_hw_output_stencil_2_write_start_pt__U2035 op_hcompute_hw_output_stencil_2_write_start (
    .in(op_hcompute_hw_output_stencil_2_write_start_in),
    .out(hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write_valid)
);
assign op_hcompute_hw_output_stencil_2_write_start_control_vars_in[2] = arr__U2044_out[2];
assign op_hcompute_hw_output_stencil_2_write_start_control_vars_in[1] = arr__U2044_out[1];
assign op_hcompute_hw_output_stencil_2_write_start_control_vars_in[0] = arr__U2044_out[0];
op_hcompute_hw_output_stencil_2_write_start_control_vars_pt__U2038 op_hcompute_hw_output_stencil_2_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_2_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_2_write_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_3_clk = clk;
assign op_hcompute_hw_output_stencil_3_conv_stencil_op_hcompute_hw_output_stencil_3_read[0] = conv_stencil_op_hcompute_hw_output_stencil_3_read[0];
cu_op_hcompute_hw_output_stencil_3 op_hcompute_hw_output_stencil_3 (
    .clk(op_hcompute_hw_output_stencil_3_clk),
    .conv_stencil_op_hcompute_hw_output_stencil_3_read(op_hcompute_hw_output_stencil_3_conv_stencil_op_hcompute_hw_output_stencil_3_read),
    .hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write(op_hcompute_hw_output_stencil_3_hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write)
);
assign op_hcompute_hw_output_stencil_3_exe_start_in = delay_reg__U2070_out;
op_hcompute_hw_output_stencil_3_exe_start_pt__U2068 op_hcompute_hw_output_stencil_3_exe_start (
    .in(op_hcompute_hw_output_stencil_3_exe_start_in),
    .out(op_hcompute_hw_output_stencil_3_exe_start_out)
);
assign op_hcompute_hw_output_stencil_3_exe_start_control_vars_in[2] = arr__U2077_out[2];
assign op_hcompute_hw_output_stencil_3_exe_start_control_vars_in[1] = arr__U2077_out[1];
assign op_hcompute_hw_output_stencil_3_exe_start_control_vars_in[0] = arr__U2077_out[0];
op_hcompute_hw_output_stencil_3_exe_start_control_vars_pt__U2071 op_hcompute_hw_output_stencil_3_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_3_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_3_exe_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_3_port_controller_clk = clk;
affine_controller__U2049 op_hcompute_hw_output_stencil_3_port_controller (
    .clk(op_hcompute_hw_output_stencil_3_port_controller_clk),
    .valid(op_hcompute_hw_output_stencil_3_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_3_port_controller_d)
);
assign op_hcompute_hw_output_stencil_3_read_start_in = op_hcompute_hw_output_stencil_3_port_controller_valid;
op_hcompute_hw_output_stencil_3_read_start_pt__U2066 op_hcompute_hw_output_stencil_3_read_start (
    .in(op_hcompute_hw_output_stencil_3_read_start_in),
    .out(op_hcompute_hw_output_stencil_3_read_start_out)
);
assign op_hcompute_hw_output_stencil_3_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_3_port_controller_d[2];
assign op_hcompute_hw_output_stencil_3_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_3_port_controller_d[1];
assign op_hcompute_hw_output_stencil_3_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_3_port_controller_d[0];
op_hcompute_hw_output_stencil_3_read_start_control_vars_pt__U2067 op_hcompute_hw_output_stencil_3_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_3_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_3_read_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_3_write_start_in = delay_reg__U2084_out;
op_hcompute_hw_output_stencil_3_write_start_pt__U2082 op_hcompute_hw_output_stencil_3_write_start (
    .in(op_hcompute_hw_output_stencil_3_write_start_in),
    .out(hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write_valid)
);
assign op_hcompute_hw_output_stencil_3_write_start_control_vars_in[2] = arr__U2091_out[2];
assign op_hcompute_hw_output_stencil_3_write_start_control_vars_in[1] = arr__U2091_out[1];
assign op_hcompute_hw_output_stencil_3_write_start_control_vars_in[0] = arr__U2091_out[0];
op_hcompute_hw_output_stencil_3_write_start_control_vars_pt__U2085 op_hcompute_hw_output_stencil_3_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_3_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_3_write_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_4_clk = clk;
assign op_hcompute_hw_output_stencil_4_conv_stencil_op_hcompute_hw_output_stencil_4_read[0] = conv_stencil_op_hcompute_hw_output_stencil_4_read[0];
cu_op_hcompute_hw_output_stencil_4 op_hcompute_hw_output_stencil_4 (
    .clk(op_hcompute_hw_output_stencil_4_clk),
    .conv_stencil_op_hcompute_hw_output_stencil_4_read(op_hcompute_hw_output_stencil_4_conv_stencil_op_hcompute_hw_output_stencil_4_read),
    .hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write(op_hcompute_hw_output_stencil_4_hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write)
);
assign op_hcompute_hw_output_stencil_4_exe_start_in = delay_reg__U2117_out;
op_hcompute_hw_output_stencil_4_exe_start_pt__U2115 op_hcompute_hw_output_stencil_4_exe_start (
    .in(op_hcompute_hw_output_stencil_4_exe_start_in),
    .out(op_hcompute_hw_output_stencil_4_exe_start_out)
);
assign op_hcompute_hw_output_stencil_4_exe_start_control_vars_in[2] = arr__U2124_out[2];
assign op_hcompute_hw_output_stencil_4_exe_start_control_vars_in[1] = arr__U2124_out[1];
assign op_hcompute_hw_output_stencil_4_exe_start_control_vars_in[0] = arr__U2124_out[0];
op_hcompute_hw_output_stencil_4_exe_start_control_vars_pt__U2118 op_hcompute_hw_output_stencil_4_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_4_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_4_exe_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_4_port_controller_clk = clk;
affine_controller__U2096 op_hcompute_hw_output_stencil_4_port_controller (
    .clk(op_hcompute_hw_output_stencil_4_port_controller_clk),
    .valid(op_hcompute_hw_output_stencil_4_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_4_port_controller_d)
);
assign op_hcompute_hw_output_stencil_4_read_start_in = op_hcompute_hw_output_stencil_4_port_controller_valid;
op_hcompute_hw_output_stencil_4_read_start_pt__U2113 op_hcompute_hw_output_stencil_4_read_start (
    .in(op_hcompute_hw_output_stencil_4_read_start_in),
    .out(op_hcompute_hw_output_stencil_4_read_start_out)
);
assign op_hcompute_hw_output_stencil_4_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_4_port_controller_d[2];
assign op_hcompute_hw_output_stencil_4_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_4_port_controller_d[1];
assign op_hcompute_hw_output_stencil_4_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_4_port_controller_d[0];
op_hcompute_hw_output_stencil_4_read_start_control_vars_pt__U2114 op_hcompute_hw_output_stencil_4_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_4_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_4_read_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_4_write_start_in = delay_reg__U2131_out;
op_hcompute_hw_output_stencil_4_write_start_pt__U2129 op_hcompute_hw_output_stencil_4_write_start (
    .in(op_hcompute_hw_output_stencil_4_write_start_in),
    .out(hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write_valid)
);
assign op_hcompute_hw_output_stencil_4_write_start_control_vars_in[2] = arr__U2138_out[2];
assign op_hcompute_hw_output_stencil_4_write_start_control_vars_in[1] = arr__U2138_out[1];
assign op_hcompute_hw_output_stencil_4_write_start_control_vars_in[0] = arr__U2138_out[0];
op_hcompute_hw_output_stencil_4_write_start_control_vars_pt__U2132 op_hcompute_hw_output_stencil_4_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_4_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_4_write_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_5_clk = clk;
assign op_hcompute_hw_output_stencil_5_conv_stencil_op_hcompute_hw_output_stencil_5_read[0] = conv_stencil_op_hcompute_hw_output_stencil_5_read[0];
cu_op_hcompute_hw_output_stencil_5 op_hcompute_hw_output_stencil_5 (
    .clk(op_hcompute_hw_output_stencil_5_clk),
    .conv_stencil_op_hcompute_hw_output_stencil_5_read(op_hcompute_hw_output_stencil_5_conv_stencil_op_hcompute_hw_output_stencil_5_read),
    .hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write(op_hcompute_hw_output_stencil_5_hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write)
);
assign op_hcompute_hw_output_stencil_5_exe_start_in = delay_reg__U2164_out;
op_hcompute_hw_output_stencil_5_exe_start_pt__U2162 op_hcompute_hw_output_stencil_5_exe_start (
    .in(op_hcompute_hw_output_stencil_5_exe_start_in),
    .out(op_hcompute_hw_output_stencil_5_exe_start_out)
);
assign op_hcompute_hw_output_stencil_5_exe_start_control_vars_in[2] = arr__U2171_out[2];
assign op_hcompute_hw_output_stencil_5_exe_start_control_vars_in[1] = arr__U2171_out[1];
assign op_hcompute_hw_output_stencil_5_exe_start_control_vars_in[0] = arr__U2171_out[0];
op_hcompute_hw_output_stencil_5_exe_start_control_vars_pt__U2165 op_hcompute_hw_output_stencil_5_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_5_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_5_exe_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_5_port_controller_clk = clk;
affine_controller__U2143 op_hcompute_hw_output_stencil_5_port_controller (
    .clk(op_hcompute_hw_output_stencil_5_port_controller_clk),
    .valid(op_hcompute_hw_output_stencil_5_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_5_port_controller_d)
);
assign op_hcompute_hw_output_stencil_5_read_start_in = op_hcompute_hw_output_stencil_5_port_controller_valid;
op_hcompute_hw_output_stencil_5_read_start_pt__U2160 op_hcompute_hw_output_stencil_5_read_start (
    .in(op_hcompute_hw_output_stencil_5_read_start_in),
    .out(op_hcompute_hw_output_stencil_5_read_start_out)
);
assign op_hcompute_hw_output_stencil_5_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_5_port_controller_d[2];
assign op_hcompute_hw_output_stencil_5_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_5_port_controller_d[1];
assign op_hcompute_hw_output_stencil_5_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_5_port_controller_d[0];
op_hcompute_hw_output_stencil_5_read_start_control_vars_pt__U2161 op_hcompute_hw_output_stencil_5_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_5_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_5_read_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_5_write_start_in = delay_reg__U2178_out;
op_hcompute_hw_output_stencil_5_write_start_pt__U2176 op_hcompute_hw_output_stencil_5_write_start (
    .in(op_hcompute_hw_output_stencil_5_write_start_in),
    .out(hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write_valid)
);
assign op_hcompute_hw_output_stencil_5_write_start_control_vars_in[2] = arr__U2185_out[2];
assign op_hcompute_hw_output_stencil_5_write_start_control_vars_in[1] = arr__U2185_out[1];
assign op_hcompute_hw_output_stencil_5_write_start_control_vars_in[0] = arr__U2185_out[0];
op_hcompute_hw_output_stencil_5_write_start_control_vars_pt__U2179 op_hcompute_hw_output_stencil_5_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_5_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_5_write_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_6_clk = clk;
assign op_hcompute_hw_output_stencil_6_conv_stencil_op_hcompute_hw_output_stencil_6_read[0] = conv_stencil_op_hcompute_hw_output_stencil_6_read[0];
cu_op_hcompute_hw_output_stencil_6 op_hcompute_hw_output_stencil_6 (
    .clk(op_hcompute_hw_output_stencil_6_clk),
    .conv_stencil_op_hcompute_hw_output_stencil_6_read(op_hcompute_hw_output_stencil_6_conv_stencil_op_hcompute_hw_output_stencil_6_read),
    .hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write(op_hcompute_hw_output_stencil_6_hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write)
);
assign op_hcompute_hw_output_stencil_6_exe_start_in = delay_reg__U2211_out;
op_hcompute_hw_output_stencil_6_exe_start_pt__U2209 op_hcompute_hw_output_stencil_6_exe_start (
    .in(op_hcompute_hw_output_stencil_6_exe_start_in),
    .out(op_hcompute_hw_output_stencil_6_exe_start_out)
);
assign op_hcompute_hw_output_stencil_6_exe_start_control_vars_in[2] = arr__U2218_out[2];
assign op_hcompute_hw_output_stencil_6_exe_start_control_vars_in[1] = arr__U2218_out[1];
assign op_hcompute_hw_output_stencil_6_exe_start_control_vars_in[0] = arr__U2218_out[0];
op_hcompute_hw_output_stencil_6_exe_start_control_vars_pt__U2212 op_hcompute_hw_output_stencil_6_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_6_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_6_exe_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_6_port_controller_clk = clk;
affine_controller__U2190 op_hcompute_hw_output_stencil_6_port_controller (
    .clk(op_hcompute_hw_output_stencil_6_port_controller_clk),
    .valid(op_hcompute_hw_output_stencil_6_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_6_port_controller_d)
);
assign op_hcompute_hw_output_stencil_6_read_start_in = op_hcompute_hw_output_stencil_6_port_controller_valid;
op_hcompute_hw_output_stencil_6_read_start_pt__U2207 op_hcompute_hw_output_stencil_6_read_start (
    .in(op_hcompute_hw_output_stencil_6_read_start_in),
    .out(op_hcompute_hw_output_stencil_6_read_start_out)
);
assign op_hcompute_hw_output_stencil_6_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_6_port_controller_d[2];
assign op_hcompute_hw_output_stencil_6_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_6_port_controller_d[1];
assign op_hcompute_hw_output_stencil_6_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_6_port_controller_d[0];
op_hcompute_hw_output_stencil_6_read_start_control_vars_pt__U2208 op_hcompute_hw_output_stencil_6_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_6_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_6_read_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_6_write_start_in = delay_reg__U2225_out;
op_hcompute_hw_output_stencil_6_write_start_pt__U2223 op_hcompute_hw_output_stencil_6_write_start (
    .in(op_hcompute_hw_output_stencil_6_write_start_in),
    .out(hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write_valid)
);
assign op_hcompute_hw_output_stencil_6_write_start_control_vars_in[2] = arr__U2232_out[2];
assign op_hcompute_hw_output_stencil_6_write_start_control_vars_in[1] = arr__U2232_out[1];
assign op_hcompute_hw_output_stencil_6_write_start_control_vars_in[0] = arr__U2232_out[0];
op_hcompute_hw_output_stencil_6_write_start_control_vars_pt__U2226 op_hcompute_hw_output_stencil_6_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_6_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_6_write_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_7_clk = clk;
assign op_hcompute_hw_output_stencil_7_conv_stencil_op_hcompute_hw_output_stencil_7_read[0] = conv_stencil_op_hcompute_hw_output_stencil_7_read[0];
cu_op_hcompute_hw_output_stencil_7 op_hcompute_hw_output_stencil_7 (
    .clk(op_hcompute_hw_output_stencil_7_clk),
    .conv_stencil_op_hcompute_hw_output_stencil_7_read(op_hcompute_hw_output_stencil_7_conv_stencil_op_hcompute_hw_output_stencil_7_read),
    .hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write(op_hcompute_hw_output_stencil_7_hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write)
);
assign op_hcompute_hw_output_stencil_7_exe_start_in = delay_reg__U2258_out;
op_hcompute_hw_output_stencil_7_exe_start_pt__U2256 op_hcompute_hw_output_stencil_7_exe_start (
    .in(op_hcompute_hw_output_stencil_7_exe_start_in),
    .out(op_hcompute_hw_output_stencil_7_exe_start_out)
);
assign op_hcompute_hw_output_stencil_7_exe_start_control_vars_in[2] = arr__U2265_out[2];
assign op_hcompute_hw_output_stencil_7_exe_start_control_vars_in[1] = arr__U2265_out[1];
assign op_hcompute_hw_output_stencil_7_exe_start_control_vars_in[0] = arr__U2265_out[0];
op_hcompute_hw_output_stencil_7_exe_start_control_vars_pt__U2259 op_hcompute_hw_output_stencil_7_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_7_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_7_exe_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_7_port_controller_clk = clk;
affine_controller__U2237 op_hcompute_hw_output_stencil_7_port_controller (
    .clk(op_hcompute_hw_output_stencil_7_port_controller_clk),
    .valid(op_hcompute_hw_output_stencil_7_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_7_port_controller_d)
);
assign op_hcompute_hw_output_stencil_7_read_start_in = op_hcompute_hw_output_stencil_7_port_controller_valid;
op_hcompute_hw_output_stencil_7_read_start_pt__U2254 op_hcompute_hw_output_stencil_7_read_start (
    .in(op_hcompute_hw_output_stencil_7_read_start_in),
    .out(op_hcompute_hw_output_stencil_7_read_start_out)
);
assign op_hcompute_hw_output_stencil_7_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_7_port_controller_d[2];
assign op_hcompute_hw_output_stencil_7_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_7_port_controller_d[1];
assign op_hcompute_hw_output_stencil_7_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_7_port_controller_d[0];
op_hcompute_hw_output_stencil_7_read_start_control_vars_pt__U2255 op_hcompute_hw_output_stencil_7_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_7_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_7_read_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_7_write_start_in = delay_reg__U2272_out;
op_hcompute_hw_output_stencil_7_write_start_pt__U2270 op_hcompute_hw_output_stencil_7_write_start (
    .in(op_hcompute_hw_output_stencil_7_write_start_in),
    .out(hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write_valid)
);
assign op_hcompute_hw_output_stencil_7_write_start_control_vars_in[2] = arr__U2279_out[2];
assign op_hcompute_hw_output_stencil_7_write_start_control_vars_in[1] = arr__U2279_out[1];
assign op_hcompute_hw_output_stencil_7_write_start_control_vars_in[0] = arr__U2279_out[0];
op_hcompute_hw_output_stencil_7_write_start_control_vars_pt__U2273 op_hcompute_hw_output_stencil_7_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_7_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_7_write_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_exe_start_in = delay_reg__U1929_out;
op_hcompute_hw_output_stencil_exe_start_pt__U1927 op_hcompute_hw_output_stencil_exe_start (
    .in(op_hcompute_hw_output_stencil_exe_start_in),
    .out(op_hcompute_hw_output_stencil_exe_start_out)
);
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[2] = arr__U1936_out[2];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[1] = arr__U1936_out[1];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[0] = arr__U1936_out[0];
op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U1930 op_hcompute_hw_output_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_port_controller_clk = clk;
affine_controller__U1908 op_hcompute_hw_output_stencil_port_controller (
    .clk(op_hcompute_hw_output_stencil_port_controller_clk),
    .valid(op_hcompute_hw_output_stencil_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_port_controller_d)
);
assign op_hcompute_hw_output_stencil_read_start_in = op_hcompute_hw_output_stencil_port_controller_valid;
op_hcompute_hw_output_stencil_read_start_pt__U1925 op_hcompute_hw_output_stencil_read_start (
    .in(op_hcompute_hw_output_stencil_read_start_in),
    .out(op_hcompute_hw_output_stencil_read_start_out)
);
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
op_hcompute_hw_output_stencil_read_start_control_vars_pt__U1926 op_hcompute_hw_output_stencil_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_write_start_in = delay_reg__U1943_out;
op_hcompute_hw_output_stencil_write_start_pt__U1941 op_hcompute_hw_output_stencil_write_start (
    .in(op_hcompute_hw_output_stencil_write_start_in),
    .out(hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write_valid)
);
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[2] = arr__U1950_out[2];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[1] = arr__U1950_out[1];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[0] = arr__U1950_out[0];
op_hcompute_hw_output_stencil_write_start_control_vars_pt__U1944 op_hcompute_hw_output_stencil_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_write_start_control_vars_out)
);
assign hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write[0] = op_hcompute_hw_output_stencil_2_hw_output_stencil_clkwrk_10_op_hcompute_hw_output_stencil_2_write[0];
assign hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write[0] = op_hcompute_hw_output_stencil_3_hw_output_stencil_clkwrk_11_op_hcompute_hw_output_stencil_3_write[0];
assign hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write[0] = op_hcompute_hw_output_stencil_4_hw_output_stencil_clkwrk_12_op_hcompute_hw_output_stencil_4_write[0];
assign hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write[0] = op_hcompute_hw_output_stencil_5_hw_output_stencil_clkwrk_13_op_hcompute_hw_output_stencil_5_write[0];
assign hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write[0] = op_hcompute_hw_output_stencil_6_hw_output_stencil_clkwrk_14_op_hcompute_hw_output_stencil_6_write[0];
assign hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write[0] = op_hcompute_hw_output_stencil_7_hw_output_stencil_clkwrk_15_op_hcompute_hw_output_stencil_7_write[0];
assign hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write[0] = op_hcompute_hw_output_stencil_hw_output_stencil_clkwrk_8_op_hcompute_hw_output_stencil_write[0];
assign hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write[0] = op_hcompute_hw_output_stencil_1_hw_output_stencil_clkwrk_9_op_hcompute_hw_output_stencil_1_write[0];
endmodule

