module bright_gauss_blur_1_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1265;
    end
  end

endmodule


module bright_gauss_blur_1_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (1259 - d0 >= 0) ? (1263) : (-1260 + d0 == 0) ? (1263) : 0;
    end
  end

endmodule


module bright_weights_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_update_0_write_wdata(output [31:0] bright_update_0_write_wdata);

endmodule


module bright(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] bright_update_0_write_wdata, input [31:0] bright_weights_update_0_read_dummy, input [287:0] bright_gauss_blur_1_update_0_read_dummy, input [0:0] bright_update_0_write_wen, output [287:0] bright_gauss_blur_1_update_0_read_rdata, input [31:0] bright_laplace_diff_0_update_0_read_dummy, output [31:0] bright_laplace_diff_0_update_0_read_rdata, output [31:0] bright_weights_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;
  logic [31:0] rd_6;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;
  reg [31:0] rd_6_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;
      rd_6_stage_1 <= rd_6;


    end

  end


  // Data processing units...
  // selector_bright_gauss_blur_1_rd1_select
  logic [0:0] selector_bright_gauss_blur_1_rd1_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd1_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd1_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd1_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd1_select_out;
  bright_gauss_blur_1_rd1_select selector_bright_gauss_blur_1_rd1_select(.clk(selector_bright_gauss_blur_1_rd1_select_clk), .rst(selector_bright_gauss_blur_1_rd1_select_rst), .d0(selector_bright_gauss_blur_1_rd1_select_d0), .d1(selector_bright_gauss_blur_1_rd1_select_d1), .out(selector_bright_gauss_blur_1_rd1_select_out));
  assign selector_bright_gauss_blur_1_rd1_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd1_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd1_select

  // selector_bright_gauss_blur_1_rd8_select
  logic [0:0] selector_bright_gauss_blur_1_rd8_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd8_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd8_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd8_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd8_select_out;
  bright_gauss_blur_1_rd8_select selector_bright_gauss_blur_1_rd8_select(.clk(selector_bright_gauss_blur_1_rd8_select_clk), .rst(selector_bright_gauss_blur_1_rd8_select_rst), .d0(selector_bright_gauss_blur_1_rd8_select_d0), .d1(selector_bright_gauss_blur_1_rd8_select_d1), .out(selector_bright_gauss_blur_1_rd8_select_out));
  assign selector_bright_gauss_blur_1_rd8_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd8_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd8_select

  // Bindings to bright_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_update_0_write_wdata;

  // selector_bright_laplace_diff_0_rd0_select
  logic [0:0] selector_bright_laplace_diff_0_rd0_select_clk;
  logic [0:0] selector_bright_laplace_diff_0_rd0_select_rst;
  logic [31:0] selector_bright_laplace_diff_0_rd0_select_d0;
  logic [31:0] selector_bright_laplace_diff_0_rd0_select_d1;
  logic [31:0] selector_bright_laplace_diff_0_rd0_select_out;
  bright_laplace_diff_0_rd0_select selector_bright_laplace_diff_0_rd0_select(.clk(selector_bright_laplace_diff_0_rd0_select_clk), .rst(selector_bright_laplace_diff_0_rd0_select_rst), .d0(selector_bright_laplace_diff_0_rd0_select_d0), .d1(selector_bright_laplace_diff_0_rd0_select_d1), .out(selector_bright_laplace_diff_0_rd0_select_out));
  assign selector_bright_laplace_diff_0_rd0_select_clk = clk;
  assign selector_bright_laplace_diff_0_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_diff_0_rd0_select

  // Bindings to bright_weights_update_0_read_dummy
    // rd_6
  assign rd_6 = bright_weights_update_0_read_dummy;

  // Bindings to bright_gauss_blur_1_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_gauss_blur_1_update_0_read_dummy;

  // selector_bright_gauss_blur_1_rd2_select
  logic [0:0] selector_bright_gauss_blur_1_rd2_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd2_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd2_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd2_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd2_select_out;
  bright_gauss_blur_1_rd2_select selector_bright_gauss_blur_1_rd2_select(.clk(selector_bright_gauss_blur_1_rd2_select_clk), .rst(selector_bright_gauss_blur_1_rd2_select_rst), .d0(selector_bright_gauss_blur_1_rd2_select_d0), .d1(selector_bright_gauss_blur_1_rd2_select_d1), .out(selector_bright_gauss_blur_1_rd2_select_out));
  assign selector_bright_gauss_blur_1_rd2_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd2_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd2_select

  // selector_bright_gauss_blur_1_rd3_select
  logic [0:0] selector_bright_gauss_blur_1_rd3_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd3_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd3_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd3_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd3_select_out;
  bright_gauss_blur_1_rd3_select selector_bright_gauss_blur_1_rd3_select(.clk(selector_bright_gauss_blur_1_rd3_select_clk), .rst(selector_bright_gauss_blur_1_rd3_select_rst), .d0(selector_bright_gauss_blur_1_rd3_select_d0), .d1(selector_bright_gauss_blur_1_rd3_select_d1), .out(selector_bright_gauss_blur_1_rd3_select_out));
  assign selector_bright_gauss_blur_1_rd3_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd3_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd3_select

  // Bindings to bright_update_0_write_wen
    // rd_0
  assign rd_0 = bright_update_0_write_wen;

  // selector_bright_gauss_blur_1_rd0_select
  logic [0:0] selector_bright_gauss_blur_1_rd0_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd0_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd0_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd0_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd0_select_out;
  bright_gauss_blur_1_rd0_select selector_bright_gauss_blur_1_rd0_select(.clk(selector_bright_gauss_blur_1_rd0_select_clk), .rst(selector_bright_gauss_blur_1_rd0_select_rst), .d0(selector_bright_gauss_blur_1_rd0_select_d0), .d1(selector_bright_gauss_blur_1_rd0_select_d1), .out(selector_bright_gauss_blur_1_rd0_select_out));
  assign selector_bright_gauss_blur_1_rd0_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd0_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd0_select

  // selector_bright_gauss_blur_1_rd4_select
  logic [0:0] selector_bright_gauss_blur_1_rd4_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd4_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd4_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd4_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd4_select_out;
  bright_gauss_blur_1_rd4_select selector_bright_gauss_blur_1_rd4_select(.clk(selector_bright_gauss_blur_1_rd4_select_clk), .rst(selector_bright_gauss_blur_1_rd4_select_rst), .d0(selector_bright_gauss_blur_1_rd4_select_d0), .d1(selector_bright_gauss_blur_1_rd4_select_d1), .out(selector_bright_gauss_blur_1_rd4_select_out));
  assign selector_bright_gauss_blur_1_rd4_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd4_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd4_select

  // selector_bright_gauss_blur_1_rd5_select
  logic [0:0] selector_bright_gauss_blur_1_rd5_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd5_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd5_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd5_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd5_select_out;
  bright_gauss_blur_1_rd5_select selector_bright_gauss_blur_1_rd5_select(.clk(selector_bright_gauss_blur_1_rd5_select_clk), .rst(selector_bright_gauss_blur_1_rd5_select_rst), .d0(selector_bright_gauss_blur_1_rd5_select_d0), .d1(selector_bright_gauss_blur_1_rd5_select_d1), .out(selector_bright_gauss_blur_1_rd5_select_out));
  assign selector_bright_gauss_blur_1_rd5_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd5_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd5_select

  // selector_bright_gauss_blur_1_rd6_select
  logic [0:0] selector_bright_gauss_blur_1_rd6_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd6_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd6_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd6_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd6_select_out;
  bright_gauss_blur_1_rd6_select selector_bright_gauss_blur_1_rd6_select(.clk(selector_bright_gauss_blur_1_rd6_select_clk), .rst(selector_bright_gauss_blur_1_rd6_select_rst), .d0(selector_bright_gauss_blur_1_rd6_select_d0), .d1(selector_bright_gauss_blur_1_rd6_select_d1), .out(selector_bright_gauss_blur_1_rd6_select_out));
  assign selector_bright_gauss_blur_1_rd6_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd6_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd6_select

  // selector_bright_gauss_blur_1_rd7_select
  logic [0:0] selector_bright_gauss_blur_1_rd7_select_clk;
  logic [0:0] selector_bright_gauss_blur_1_rd7_select_rst;
  logic [31:0] selector_bright_gauss_blur_1_rd7_select_d0;
  logic [31:0] selector_bright_gauss_blur_1_rd7_select_d1;
  logic [31:0] selector_bright_gauss_blur_1_rd7_select_out;
  bright_gauss_blur_1_rd7_select selector_bright_gauss_blur_1_rd7_select(.clk(selector_bright_gauss_blur_1_rd7_select_clk), .rst(selector_bright_gauss_blur_1_rd7_select_rst), .d0(selector_bright_gauss_blur_1_rd7_select_d0), .d1(selector_bright_gauss_blur_1_rd7_select_d1), .out(selector_bright_gauss_blur_1_rd7_select_out));
  assign selector_bright_gauss_blur_1_rd7_select_clk = clk;
  assign selector_bright_gauss_blur_1_rd7_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_1_rd7_select

  // Bindings to bright_gauss_blur_1_update_0_read_rdata
    // wr_3
  assign bright_gauss_blur_1_update_0_read_rdata = rd_2;

  // selector_bright_weights_rd0_select
  logic [0:0] selector_bright_weights_rd0_select_clk;
  logic [0:0] selector_bright_weights_rd0_select_rst;
  logic [31:0] selector_bright_weights_rd0_select_d0;
  logic [31:0] selector_bright_weights_rd0_select_d1;
  logic [31:0] selector_bright_weights_rd0_select_out;
  bright_weights_rd0_select selector_bright_weights_rd0_select(.clk(selector_bright_weights_rd0_select_clk), .rst(selector_bright_weights_rd0_select_rst), .d0(selector_bright_weights_rd0_select_d0), .d1(selector_bright_weights_rd0_select_d1), .out(selector_bright_weights_rd0_select_out));
  assign selector_bright_weights_rd0_select_clk = clk;
  assign selector_bright_weights_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_rd0_select

  // bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0
  logic [0:0] bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_clk;
  logic [0:0] bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_rst;
  logic [0:0] bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_start;
  logic [0:0] bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_done;
  bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0 bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0(.clk(bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_clk), .rst(bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_rst), .start(bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_start), .done(bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_done));
  assign bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_clk = clk;
  assign bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0_rst = rst;
  // Bindings to bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0

  // Bindings to bright_laplace_diff_0_update_0_read_dummy
    // rd_4
  assign rd_4 = bright_laplace_diff_0_update_0_read_dummy;

  // Bindings to bright_laplace_diff_0_update_0_read_rdata
    // wr_5
  assign bright_laplace_diff_0_update_0_read_rdata = rd_4;

  // Bindings to bright_weights_update_0_read_rdata
    // wr_7
  assign bright_weights_update_0_read_rdata = rd_6;

  // bright_bright_update_0_write0_merged_banks_10
  logic [0:0] bright_bright_update_0_write0_merged_banks_10_clk;
  logic [0:0] bright_bright_update_0_write0_merged_banks_10_rst;
  logic [0:0] bright_bright_update_0_write0_merged_banks_10_start;
  logic [0:0] bright_bright_update_0_write0_merged_banks_10_done;
  bright_bright_update_0_write0_merged_banks_10 bright_bright_update_0_write0_merged_banks_10(.clk(bright_bright_update_0_write0_merged_banks_10_clk), .rst(bright_bright_update_0_write0_merged_banks_10_rst), .start(bright_bright_update_0_write0_merged_banks_10_start), .done(bright_bright_update_0_write0_merged_banks_10_done));
  assign bright_bright_update_0_write0_merged_banks_10_clk = clk;
  assign bright_bright_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to bright_bright_update_0_write0_merged_banks_10



endmodule


module in_wire_bright_gauss_blur_1_update_0_read_dummy(output [287:0] bright_gauss_blur_1_update_0_read_dummy);

endmodule


module bright_gauss_blur_1_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2527;
    end
  end

endmodule


module bright_gauss_blur_1_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1264;
    end
  end

endmodule


module bright_gauss_blur_1_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module bright_gauss_blur_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2528;
    end
  end

endmodule


module bright_gauss_blur_1_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module in_wire_bright_update_0_write_wen(output [0:0] bright_update_0_write_wen);

endmodule


module bright_gauss_blur_1_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (1259 - d0 >= 0) ? (2526) : (-1260 + d0 == 0) ? (2526) : 0;
    end
  end

endmodule


module bright_gauss_blur_1_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module out_wire_bright_gauss_blur_1_update_0_read_rdata(input [287:0] bright_gauss_blur_1_update_0_read_rdata);

endmodule


module in_wire_bright_laplace_diff_0_update_0_read_dummy(output [31:0] bright_laplace_diff_0_update_0_read_dummy);

endmodule


module out_wire_bright_laplace_diff_0_update_0_read_rdata(input [31:0] bright_laplace_diff_0_update_0_read_rdata);

endmodule


module in_wire_bright_weights_update_0_read_dummy(output [31:0] bright_weights_update_0_read_dummy);

endmodule


module out_wire_bright_weights_update_0_read_rdata(input [31:0] bright_weights_update_0_read_rdata);

endmodule


module bright_gauss_blur_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] bright_gauss_ds_1_update_0_read_rdata, input [31:0] bright_gauss_ds_1_update_0_read_dummy, input [31:0] bright_gauss_blur_1_update_0_write_wdata, input [0:0] bright_gauss_blur_1_update_0_write_wen);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to bright_gauss_ds_1_update_0_read_rdata
    // wr_3
  assign bright_gauss_ds_1_update_0_read_rdata = rd_2;

  // Bindings to bright_gauss_ds_1_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_gauss_ds_1_update_0_read_dummy;

  // Bindings to bright_gauss_blur_1_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_gauss_blur_1_update_0_write_wdata;

  // bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1
  logic [0:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_done;
  bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1 bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1(.clk(bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_clk), .rst(bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_rst), .start(bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_start), .done(bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_done));
  assign bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_clk = clk;
  assign bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1

  // selector_bright_gauss_ds_1_rd0_select
  logic [0:0] selector_bright_gauss_ds_1_rd0_select_clk;
  logic [0:0] selector_bright_gauss_ds_1_rd0_select_rst;
  logic [31:0] selector_bright_gauss_ds_1_rd0_select_d0;
  logic [31:0] selector_bright_gauss_ds_1_rd0_select_d1;
  logic [31:0] selector_bright_gauss_ds_1_rd0_select_out;
  bright_gauss_ds_1_rd0_select selector_bright_gauss_ds_1_rd0_select(.clk(selector_bright_gauss_ds_1_rd0_select_clk), .rst(selector_bright_gauss_ds_1_rd0_select_rst), .d0(selector_bright_gauss_ds_1_rd0_select_d0), .d1(selector_bright_gauss_ds_1_rd0_select_d1), .out(selector_bright_gauss_ds_1_rd0_select_out));
  assign selector_bright_gauss_ds_1_rd0_select_clk = clk;
  assign selector_bright_gauss_ds_1_rd0_select_rst = rst;
  // Bindings to selector_bright_gauss_ds_1_rd0_select

  // Bindings to bright_gauss_blur_1_update_0_write_wen
    // rd_0
  assign rd_0 = bright_gauss_blur_1_update_0_write_wen;



endmodule


module bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268



endmodule


module in_wire_bright_gauss_ds_3_update_0_write_wen(output [0:0] bright_gauss_ds_3_update_0_write_wen);

endmodule


module bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module bright_laplace_us_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = ((-1 - d1) % 2 == 0 && 311 - d0 >= 0) ? ((156 - floord(2*d0, 4))) : 0;
    end
  end

endmodule


module in_wire_bright_weights_update_0_write_wen(output [0:0] bright_weights_update_0_write_wen);

endmodule


module in_wire_bright_weights_update_0_write_wdata(output [31:0] bright_weights_update_0_write_wdata);

endmodule


module in_wire_bright_weights_normed_update_0_read_dummy(output [31:0] bright_weights_normed_update_0_read_dummy);

endmodule


module out_wire_bright_weights_normed_update_0_read_rdata(input [31:0] bright_weights_normed_update_0_read_rdata);

endmodule


module in_wire_weight_sums_update_0_read_dummy(output [31:0] weight_sums_update_0_read_dummy);

endmodule


module out_wire_weight_sums_update_0_read_rdata(input [31:0] weight_sums_update_0_read_rdata);

endmodule


module bright_weights_normed_gauss_blur_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2528;
    end
  end

endmodule


module bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_1260 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_1260 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16



endmodule


module bright_weights_normed_gauss_blur_1_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (1259 - d0 >= 0) ? (2526) : (-1260 + d0 == 0) ? (2526) : 0;
    end
  end

endmodule


module bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_16431 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f314
  logic [0:0] f314_wen;
  logic [31:0] f314_wdata;
  logic [0:0] f314_clk;
  logic [0:0] f314_rst;
  logic [31:0] f314_rdata;
  sr_buffer_32_1 f314(.wen(f314_wen), .wdata(f314_wdata), .clk(f314_clk), .rst(f314_rst), .rdata(f314_rdata));
  assign f314_clk = clk;
  assign f314_rst = rst;
  // Bindings to f314

  // f316
  logic [0:0] f316_wen;
  logic [31:0] f316_wdata;
  logic [0:0] f316_clk;
  logic [0:0] f316_rst;
  logic [31:0] f316_rdata;
  sr_buffer_32_1 f316(.wen(f316_wen), .wdata(f316_wdata), .clk(f316_clk), .rst(f316_rst), .rdata(f316_rdata));
  assign f316_clk = clk;
  assign f316_rst = rst;
  // Bindings to f316

  // f318
  logic [0:0] f318_wen;
  logic [31:0] f318_wdata;
  logic [0:0] f318_clk;
  logic [0:0] f318_rst;
  logic [31:0] f318_rdata;
  sr_buffer_32_1 f318(.wen(f318_wen), .wdata(f318_wdata), .clk(f318_clk), .rst(f318_rst), .rdata(f318_rdata));
  assign f318_clk = clk;
  assign f318_rst = rst;
  // Bindings to f318

  // f320
  logic [0:0] f320_wen;
  logic [31:0] f320_wdata;
  logic [0:0] f320_clk;
  logic [0:0] f320_rst;
  logic [31:0] f320_rdata;
  sr_buffer_32_1 f320(.wen(f320_wen), .wdata(f320_wdata), .clk(f320_clk), .rst(f320_rst), .rdata(f320_rdata));
  assign f320_clk = clk;
  assign f320_rst = rst;
  // Bindings to f320

  // f322
  logic [0:0] f322_wen;
  logic [31:0] f322_wdata;
  logic [0:0] f322_clk;
  logic [0:0] f322_rst;
  logic [31:0] f322_rdata;
  sr_buffer_32_1 f322(.wen(f322_wen), .wdata(f322_wdata), .clk(f322_clk), .rst(f322_rst), .rdata(f322_rdata));
  assign f322_clk = clk;
  assign f322_rst = rst;
  // Bindings to f322

  // f324
  logic [0:0] f324_wen;
  logic [31:0] f324_wdata;
  logic [0:0] f324_clk;
  logic [0:0] f324_rst;
  logic [31:0] f324_rdata;
  sr_buffer_32_1 f324(.wen(f324_wen), .wdata(f324_wdata), .clk(f324_clk), .rst(f324_rst), .rdata(f324_rdata));
  assign f324_clk = clk;
  assign f324_rst = rst;
  // Bindings to f324

  // f326
  logic [0:0] f326_wen;
  logic [31:0] f326_wdata;
  logic [0:0] f326_clk;
  logic [0:0] f326_rst;
  logic [31:0] f326_rdata;
  sr_buffer_32_1 f326(.wen(f326_wen), .wdata(f326_wdata), .clk(f326_clk), .rst(f326_rst), .rdata(f326_rdata));
  assign f326_clk = clk;
  assign f326_rst = rst;
  // Bindings to f326

  // f328
  logic [0:0] f328_wen;
  logic [31:0] f328_wdata;
  logic [0:0] f328_clk;
  logic [0:0] f328_rst;
  logic [31:0] f328_rdata;
  sr_buffer_32_1 f328(.wen(f328_wen), .wdata(f328_wdata), .clk(f328_clk), .rst(f328_rst), .rdata(f328_rdata));
  assign f328_clk = clk;
  assign f328_rst = rst;
  // Bindings to f328

  // f330
  logic [0:0] f330_wen;
  logic [31:0] f330_wdata;
  logic [0:0] f330_clk;
  logic [0:0] f330_rst;
  logic [31:0] f330_rdata;
  sr_buffer_32_1 f330(.wen(f330_wen), .wdata(f330_wdata), .clk(f330_clk), .rst(f330_rst), .rdata(f330_rdata));
  assign f330_clk = clk;
  assign f330_rst = rst;
  // Bindings to f330

  // f332
  logic [0:0] f332_wen;
  logic [31:0] f332_wdata;
  logic [0:0] f332_clk;
  logic [0:0] f332_rst;
  logic [31:0] f332_rdata;
  sr_buffer_32_1 f332(.wen(f332_wen), .wdata(f332_wdata), .clk(f332_clk), .rst(f332_rst), .rdata(f332_rdata));
  assign f332_clk = clk;
  assign f332_rst = rst;
  // Bindings to f332

  // f334
  logic [0:0] f334_wen;
  logic [31:0] f334_wdata;
  logic [0:0] f334_clk;
  logic [0:0] f334_rst;
  logic [31:0] f334_rdata;
  sr_buffer_32_1 f334(.wen(f334_wen), .wdata(f334_wdata), .clk(f334_clk), .rst(f334_rst), .rdata(f334_rdata));
  assign f334_clk = clk;
  assign f334_rst = rst;
  // Bindings to f334

  // f336
  logic [0:0] f336_wen;
  logic [31:0] f336_wdata;
  logic [0:0] f336_clk;
  logic [0:0] f336_rst;
  logic [31:0] f336_rdata;
  sr_buffer_32_1 f336(.wen(f336_wen), .wdata(f336_wdata), .clk(f336_clk), .rst(f336_rst), .rdata(f336_rdata));
  assign f336_clk = clk;
  assign f336_rst = rst;
  // Bindings to f336

  // f338
  logic [0:0] f338_wen;
  logic [31:0] f338_wdata;
  logic [0:0] f338_clk;
  logic [0:0] f338_rst;
  logic [31:0] f338_rdata;
  sr_buffer_32_1 f338(.wen(f338_wen), .wdata(f338_wdata), .clk(f338_clk), .rst(f338_rst), .rdata(f338_rdata));
  assign f338_clk = clk;
  assign f338_rst = rst;
  // Bindings to f338

  // f340
  logic [0:0] f340_wen;
  logic [31:0] f340_wdata;
  logic [0:0] f340_clk;
  logic [0:0] f340_rst;
  logic [31:0] f340_rdata;
  sr_buffer_32_1 f340(.wen(f340_wen), .wdata(f340_wdata), .clk(f340_clk), .rst(f340_rst), .rdata(f340_rdata));
  assign f340_clk = clk;
  assign f340_rst = rst;
  // Bindings to f340

  // f342
  logic [0:0] f342_wen;
  logic [31:0] f342_wdata;
  logic [0:0] f342_clk;
  logic [0:0] f342_rst;
  logic [31:0] f342_rdata;
  sr_buffer_32_1 f342(.wen(f342_wen), .wdata(f342_wdata), .clk(f342_clk), .rst(f342_rst), .rdata(f342_rdata));
  assign f342_clk = clk;
  assign f342_rst = rst;
  // Bindings to f342

  // f344
  logic [0:0] f344_wen;
  logic [31:0] f344_wdata;
  logic [0:0] f344_clk;
  logic [0:0] f344_rst;
  logic [31:0] f344_rdata;
  sr_buffer_32_1 f344(.wen(f344_wen), .wdata(f344_wdata), .clk(f344_clk), .rst(f344_rst), .rdata(f344_rdata));
  assign f344_clk = clk;
  assign f344_rst = rst;
  // Bindings to f344

  // f346
  logic [0:0] f346_wen;
  logic [31:0] f346_wdata;
  logic [0:0] f346_clk;
  logic [0:0] f346_rst;
  logic [31:0] f346_rdata;
  sr_buffer_32_1 f346(.wen(f346_wen), .wdata(f346_wdata), .clk(f346_clk), .rst(f346_rst), .rdata(f346_rdata));
  assign f346_clk = clk;
  assign f346_rst = rst;
  // Bindings to f346

  // f348
  logic [0:0] f348_wen;
  logic [31:0] f348_wdata;
  logic [0:0] f348_clk;
  logic [0:0] f348_rst;
  logic [31:0] f348_rdata;
  sr_buffer_32_1 f348(.wen(f348_wen), .wdata(f348_wdata), .clk(f348_clk), .rst(f348_rst), .rdata(f348_rdata));
  assign f348_clk = clk;
  assign f348_rst = rst;
  // Bindings to f348

  // f350
  logic [0:0] f350_wen;
  logic [31:0] f350_wdata;
  logic [0:0] f350_clk;
  logic [0:0] f350_rst;
  logic [31:0] f350_rdata;
  sr_buffer_32_1 f350(.wen(f350_wen), .wdata(f350_wdata), .clk(f350_clk), .rst(f350_rst), .rdata(f350_rdata));
  assign f350_clk = clk;
  assign f350_rst = rst;
  // Bindings to f350

  // f352
  logic [0:0] f352_wen;
  logic [31:0] f352_wdata;
  logic [0:0] f352_clk;
  logic [0:0] f352_rst;
  logic [31:0] f352_rdata;
  sr_buffer_32_1 f352(.wen(f352_wen), .wdata(f352_wdata), .clk(f352_clk), .rst(f352_rst), .rdata(f352_rdata));
  assign f352_clk = clk;
  assign f352_rst = rst;
  // Bindings to f352

  // f354
  logic [0:0] f354_wen;
  logic [31:0] f354_wdata;
  logic [0:0] f354_clk;
  logic [0:0] f354_rst;
  logic [31:0] f354_rdata;
  sr_buffer_32_1 f354(.wen(f354_wen), .wdata(f354_wdata), .clk(f354_clk), .rst(f354_rst), .rdata(f354_rdata));
  assign f354_clk = clk;
  assign f354_rst = rst;
  // Bindings to f354

  // f356
  logic [0:0] f356_wen;
  logic [31:0] f356_wdata;
  logic [0:0] f356_clk;
  logic [0:0] f356_rst;
  logic [31:0] f356_rdata;
  sr_buffer_32_1 f356(.wen(f356_wen), .wdata(f356_wdata), .clk(f356_clk), .rst(f356_rst), .rdata(f356_rdata));
  assign f356_clk = clk;
  assign f356_rst = rst;
  // Bindings to f356

  // f358
  logic [0:0] f358_wen;
  logic [31:0] f358_wdata;
  logic [0:0] f358_clk;
  logic [0:0] f358_rst;
  logic [31:0] f358_rdata;
  sr_buffer_32_1 f358(.wen(f358_wen), .wdata(f358_wdata), .clk(f358_clk), .rst(f358_rst), .rdata(f358_rdata));
  assign f358_clk = clk;
  assign f358_rst = rst;
  // Bindings to f358

  // f360
  logic [0:0] f360_wen;
  logic [31:0] f360_wdata;
  logic [0:0] f360_clk;
  logic [0:0] f360_rst;
  logic [31:0] f360_rdata;
  sr_buffer_32_1 f360(.wen(f360_wen), .wdata(f360_wdata), .clk(f360_clk), .rst(f360_rst), .rdata(f360_rdata));
  assign f360_clk = clk;
  assign f360_rst = rst;
  // Bindings to f360

  // f362
  logic [0:0] f362_wen;
  logic [31:0] f362_wdata;
  logic [0:0] f362_clk;
  logic [0:0] f362_rst;
  logic [31:0] f362_rdata;
  sr_buffer_32_1 f362(.wen(f362_wen), .wdata(f362_wdata), .clk(f362_clk), .rst(f362_rst), .rdata(f362_rdata));
  assign f362_clk = clk;
  assign f362_rst = rst;
  // Bindings to f362

  // f364
  logic [0:0] f364_wen;
  logic [31:0] f364_wdata;
  logic [0:0] f364_clk;
  logic [0:0] f364_rst;
  logic [31:0] f364_rdata;
  sr_buffer_32_1 f364(.wen(f364_wen), .wdata(f364_wdata), .clk(f364_clk), .rst(f364_rst), .rdata(f364_rdata));
  assign f364_clk = clk;
  assign f364_rst = rst;
  // Bindings to f364

  // f366
  logic [0:0] f366_wen;
  logic [31:0] f366_wdata;
  logic [0:0] f366_clk;
  logic [0:0] f366_rst;
  logic [31:0] f366_rdata;
  sr_buffer_32_1 f366(.wen(f366_wen), .wdata(f366_wdata), .clk(f366_clk), .rst(f366_rst), .rdata(f366_rdata));
  assign f366_clk = clk;
  assign f366_rst = rst;
  // Bindings to f366

  // f368
  logic [0:0] f368_wen;
  logic [31:0] f368_wdata;
  logic [0:0] f368_clk;
  logic [0:0] f368_rst;
  logic [31:0] f368_rdata;
  sr_buffer_32_1 f368(.wen(f368_wen), .wdata(f368_wdata), .clk(f368_clk), .rst(f368_rst), .rdata(f368_rdata));
  assign f368_clk = clk;
  assign f368_rst = rst;
  // Bindings to f368

  // f370
  logic [0:0] f370_wen;
  logic [31:0] f370_wdata;
  logic [0:0] f370_clk;
  logic [0:0] f370_rst;
  logic [31:0] f370_rdata;
  sr_buffer_32_1 f370(.wen(f370_wen), .wdata(f370_wdata), .clk(f370_clk), .rst(f370_rst), .rdata(f370_rdata));
  assign f370_clk = clk;
  assign f370_rst = rst;
  // Bindings to f370

  // f372
  logic [0:0] f372_wen;
  logic [31:0] f372_wdata;
  logic [0:0] f372_clk;
  logic [0:0] f372_rst;
  logic [31:0] f372_rdata;
  sr_buffer_32_1 f372(.wen(f372_wen), .wdata(f372_wdata), .clk(f372_clk), .rst(f372_rst), .rdata(f372_rdata));
  assign f372_clk = clk;
  assign f372_rst = rst;
  // Bindings to f372

  // f374
  logic [0:0] f374_wen;
  logic [31:0] f374_wdata;
  logic [0:0] f374_clk;
  logic [0:0] f374_rst;
  logic [31:0] f374_rdata;
  sr_buffer_32_1 f374(.wen(f374_wen), .wdata(f374_wdata), .clk(f374_clk), .rst(f374_rst), .rdata(f374_rdata));
  assign f374_clk = clk;
  assign f374_rst = rst;
  // Bindings to f374

  // f376
  logic [0:0] f376_wen;
  logic [31:0] f376_wdata;
  logic [0:0] f376_clk;
  logic [0:0] f376_rst;
  logic [31:0] f376_rdata;
  sr_buffer_32_1 f376(.wen(f376_wen), .wdata(f376_wdata), .clk(f376_clk), .rst(f376_rst), .rdata(f376_rdata));
  assign f376_clk = clk;
  assign f376_rst = rst;
  // Bindings to f376

  // f378
  logic [0:0] f378_wen;
  logic [31:0] f378_wdata;
  logic [0:0] f378_clk;
  logic [0:0] f378_rst;
  logic [31:0] f378_rdata;
  sr_buffer_32_1 f378(.wen(f378_wen), .wdata(f378_wdata), .clk(f378_clk), .rst(f378_rst), .rdata(f378_rdata));
  assign f378_clk = clk;
  assign f378_rst = rst;
  // Bindings to f378

  // f380
  logic [0:0] f380_wen;
  logic [31:0] f380_wdata;
  logic [0:0] f380_clk;
  logic [0:0] f380_rst;
  logic [31:0] f380_rdata;
  sr_buffer_32_1 f380(.wen(f380_wen), .wdata(f380_wdata), .clk(f380_clk), .rst(f380_rst), .rdata(f380_rdata));
  assign f380_clk = clk;
  assign f380_rst = rst;
  // Bindings to f380

  // f382
  logic [0:0] f382_wen;
  logic [31:0] f382_wdata;
  logic [0:0] f382_clk;
  logic [0:0] f382_rst;
  logic [31:0] f382_rdata;
  sr_buffer_32_1 f382(.wen(f382_wen), .wdata(f382_wdata), .clk(f382_clk), .rst(f382_rst), .rdata(f382_rdata));
  assign f382_clk = clk;
  assign f382_rst = rst;
  // Bindings to f382

  // f384
  logic [0:0] f384_wen;
  logic [31:0] f384_wdata;
  logic [0:0] f384_clk;
  logic [0:0] f384_rst;
  logic [31:0] f384_rdata;
  sr_buffer_32_1 f384(.wen(f384_wen), .wdata(f384_wdata), .clk(f384_clk), .rst(f384_rst), .rdata(f384_rdata));
  assign f384_clk = clk;
  assign f384_rst = rst;
  // Bindings to f384

  // f386
  logic [0:0] f386_wen;
  logic [31:0] f386_wdata;
  logic [0:0] f386_clk;
  logic [0:0] f386_rst;
  logic [31:0] f386_rdata;
  sr_buffer_32_1 f386(.wen(f386_wen), .wdata(f386_wdata), .clk(f386_clk), .rst(f386_rst), .rdata(f386_rdata));
  assign f386_clk = clk;
  assign f386_rst = rst;
  // Bindings to f386

  // f388
  logic [0:0] f388_wen;
  logic [31:0] f388_wdata;
  logic [0:0] f388_clk;
  logic [0:0] f388_rst;
  logic [31:0] f388_rdata;
  sr_buffer_32_1 f388(.wen(f388_wen), .wdata(f388_wdata), .clk(f388_clk), .rst(f388_rst), .rdata(f388_rdata));
  assign f388_clk = clk;
  assign f388_rst = rst;
  // Bindings to f388

  // f390
  logic [0:0] f390_wen;
  logic [31:0] f390_wdata;
  logic [0:0] f390_clk;
  logic [0:0] f390_rst;
  logic [31:0] f390_rdata;
  sr_buffer_32_1 f390(.wen(f390_wen), .wdata(f390_wdata), .clk(f390_clk), .rst(f390_rst), .rdata(f390_rdata));
  assign f390_clk = clk;
  assign f390_rst = rst;
  // Bindings to f390

  // f392
  logic [0:0] f392_wen;
  logic [31:0] f392_wdata;
  logic [0:0] f392_clk;
  logic [0:0] f392_rst;
  logic [31:0] f392_rdata;
  sr_buffer_32_1 f392(.wen(f392_wen), .wdata(f392_wdata), .clk(f392_clk), .rst(f392_rst), .rdata(f392_rdata));
  assign f392_clk = clk;
  assign f392_rst = rst;
  // Bindings to f392

  // f394
  logic [0:0] f394_wen;
  logic [31:0] f394_wdata;
  logic [0:0] f394_clk;
  logic [0:0] f394_rst;
  logic [31:0] f394_rdata;
  sr_buffer_32_1 f394(.wen(f394_wen), .wdata(f394_wdata), .clk(f394_clk), .rst(f394_rst), .rdata(f394_rdata));
  assign f394_clk = clk;
  assign f394_rst = rst;
  // Bindings to f394

  // f396
  logic [0:0] f396_wen;
  logic [31:0] f396_wdata;
  logic [0:0] f396_clk;
  logic [0:0] f396_rst;
  logic [31:0] f396_rdata;
  sr_buffer_32_1 f396(.wen(f396_wen), .wdata(f396_wdata), .clk(f396_clk), .rst(f396_rst), .rdata(f396_rdata));
  assign f396_clk = clk;
  assign f396_rst = rst;
  // Bindings to f396

  // f398
  logic [0:0] f398_wen;
  logic [31:0] f398_wdata;
  logic [0:0] f398_clk;
  logic [0:0] f398_rst;
  logic [31:0] f398_rdata;
  sr_buffer_32_1 f398(.wen(f398_wen), .wdata(f398_wdata), .clk(f398_clk), .rst(f398_rst), .rdata(f398_rdata));
  assign f398_clk = clk;
  assign f398_rst = rst;
  // Bindings to f398

  // f400
  logic [0:0] f400_wen;
  logic [31:0] f400_wdata;
  logic [0:0] f400_clk;
  logic [0:0] f400_rst;
  logic [31:0] f400_rdata;
  sr_buffer_32_1 f400(.wen(f400_wen), .wdata(f400_wdata), .clk(f400_clk), .rst(f400_rst), .rdata(f400_rdata));
  assign f400_clk = clk;
  assign f400_rst = rst;
  // Bindings to f400

  // f402
  logic [0:0] f402_wen;
  logic [31:0] f402_wdata;
  logic [0:0] f402_clk;
  logic [0:0] f402_rst;
  logic [31:0] f402_rdata;
  sr_buffer_32_1 f402(.wen(f402_wen), .wdata(f402_wdata), .clk(f402_clk), .rst(f402_rst), .rdata(f402_rdata));
  assign f402_clk = clk;
  assign f402_rst = rst;
  // Bindings to f402

  // f404
  logic [0:0] f404_wen;
  logic [31:0] f404_wdata;
  logic [0:0] f404_clk;
  logic [0:0] f404_rst;
  logic [31:0] f404_rdata;
  sr_buffer_32_1 f404(.wen(f404_wen), .wdata(f404_wdata), .clk(f404_clk), .rst(f404_rst), .rdata(f404_rdata));
  assign f404_clk = clk;
  assign f404_rst = rst;
  // Bindings to f404

  // f406
  logic [0:0] f406_wen;
  logic [31:0] f406_wdata;
  logic [0:0] f406_clk;
  logic [0:0] f406_rst;
  logic [31:0] f406_rdata;
  sr_buffer_32_1 f406(.wen(f406_wen), .wdata(f406_wdata), .clk(f406_clk), .rst(f406_rst), .rdata(f406_rdata));
  assign f406_clk = clk;
  assign f406_rst = rst;
  // Bindings to f406

  // f408
  logic [0:0] f408_wen;
  logic [31:0] f408_wdata;
  logic [0:0] f408_clk;
  logic [0:0] f408_rst;
  logic [31:0] f408_rdata;
  sr_buffer_32_1 f408(.wen(f408_wen), .wdata(f408_wdata), .clk(f408_clk), .rst(f408_rst), .rdata(f408_rdata));
  assign f408_clk = clk;
  assign f408_rst = rst;
  // Bindings to f408

  // f410
  logic [0:0] f410_wen;
  logic [31:0] f410_wdata;
  logic [0:0] f410_clk;
  logic [0:0] f410_rst;
  logic [31:0] f410_rdata;
  sr_buffer_32_1 f410(.wen(f410_wen), .wdata(f410_wdata), .clk(f410_clk), .rst(f410_rst), .rdata(f410_rdata));
  assign f410_clk = clk;
  assign f410_rst = rst;
  // Bindings to f410

  // f412
  logic [0:0] f412_wen;
  logic [31:0] f412_wdata;
  logic [0:0] f412_clk;
  logic [0:0] f412_rst;
  logic [31:0] f412_rdata;
  sr_buffer_32_1 f412(.wen(f412_wen), .wdata(f412_wdata), .clk(f412_clk), .rst(f412_rst), .rdata(f412_rdata));
  assign f412_clk = clk;
  assign f412_rst = rst;
  // Bindings to f412

  // f414
  logic [0:0] f414_wen;
  logic [31:0] f414_wdata;
  logic [0:0] f414_clk;
  logic [0:0] f414_rst;
  logic [31:0] f414_rdata;
  sr_buffer_32_1 f414(.wen(f414_wen), .wdata(f414_wdata), .clk(f414_clk), .rst(f414_rst), .rdata(f414_rdata));
  assign f414_clk = clk;
  assign f414_rst = rst;
  // Bindings to f414

  // f416
  logic [0:0] f416_wen;
  logic [31:0] f416_wdata;
  logic [0:0] f416_clk;
  logic [0:0] f416_rst;
  logic [31:0] f416_rdata;
  sr_buffer_32_1 f416(.wen(f416_wen), .wdata(f416_wdata), .clk(f416_clk), .rst(f416_rst), .rdata(f416_rdata));
  assign f416_clk = clk;
  assign f416_rst = rst;
  // Bindings to f416

  // f418
  logic [0:0] f418_wen;
  logic [31:0] f418_wdata;
  logic [0:0] f418_clk;
  logic [0:0] f418_rst;
  logic [31:0] f418_rdata;
  sr_buffer_32_1 f418(.wen(f418_wen), .wdata(f418_wdata), .clk(f418_clk), .rst(f418_rst), .rdata(f418_rdata));
  assign f418_clk = clk;
  assign f418_rst = rst;
  // Bindings to f418

  // f420
  logic [0:0] f420_wen;
  logic [31:0] f420_wdata;
  logic [0:0] f420_clk;
  logic [0:0] f420_rst;
  logic [31:0] f420_rdata;
  sr_buffer_32_1 f420(.wen(f420_wen), .wdata(f420_wdata), .clk(f420_clk), .rst(f420_rst), .rdata(f420_rdata));
  assign f420_clk = clk;
  assign f420_rst = rst;
  // Bindings to f420

  // f422
  logic [0:0] f422_wen;
  logic [31:0] f422_wdata;
  logic [0:0] f422_clk;
  logic [0:0] f422_rst;
  logic [31:0] f422_rdata;
  sr_buffer_32_1 f422(.wen(f422_wen), .wdata(f422_wdata), .clk(f422_clk), .rst(f422_rst), .rdata(f422_rdata));
  assign f422_clk = clk;
  assign f422_rst = rst;
  // Bindings to f422

  // f424
  logic [0:0] f424_wen;
  logic [31:0] f424_wdata;
  logic [0:0] f424_clk;
  logic [0:0] f424_rst;
  logic [31:0] f424_rdata;
  sr_buffer_32_1 f424(.wen(f424_wen), .wdata(f424_wdata), .clk(f424_clk), .rst(f424_rst), .rdata(f424_rdata));
  assign f424_clk = clk;
  assign f424_rst = rst;
  // Bindings to f424

  // f426
  logic [0:0] f426_wen;
  logic [31:0] f426_wdata;
  logic [0:0] f426_clk;
  logic [0:0] f426_rst;
  logic [31:0] f426_rdata;
  sr_buffer_32_1 f426(.wen(f426_wen), .wdata(f426_wdata), .clk(f426_clk), .rst(f426_rst), .rdata(f426_rdata));
  assign f426_clk = clk;
  assign f426_rst = rst;
  // Bindings to f426

  // f428
  logic [0:0] f428_wen;
  logic [31:0] f428_wdata;
  logic [0:0] f428_clk;
  logic [0:0] f428_rst;
  logic [31:0] f428_rdata;
  sr_buffer_32_1 f428(.wen(f428_wen), .wdata(f428_wdata), .clk(f428_clk), .rst(f428_rst), .rdata(f428_rdata));
  assign f428_clk = clk;
  assign f428_rst = rst;
  // Bindings to f428

  // f430
  logic [0:0] f430_wen;
  logic [31:0] f430_wdata;
  logic [0:0] f430_clk;
  logic [0:0] f430_rst;
  logic [31:0] f430_rdata;
  sr_buffer_32_1 f430(.wen(f430_wen), .wdata(f430_wdata), .clk(f430_clk), .rst(f430_rst), .rdata(f430_rdata));
  assign f430_clk = clk;
  assign f430_rst = rst;
  // Bindings to f430

  // f432
  logic [0:0] f432_wen;
  logic [31:0] f432_wdata;
  logic [0:0] f432_clk;
  logic [0:0] f432_rst;
  logic [31:0] f432_rdata;
  sr_buffer_32_1 f432(.wen(f432_wen), .wdata(f432_wdata), .clk(f432_clk), .rst(f432_rst), .rdata(f432_rdata));
  assign f432_clk = clk;
  assign f432_rst = rst;
  // Bindings to f432

  // f434
  logic [0:0] f434_wen;
  logic [31:0] f434_wdata;
  logic [0:0] f434_clk;
  logic [0:0] f434_rst;
  logic [31:0] f434_rdata;
  sr_buffer_32_1 f434(.wen(f434_wen), .wdata(f434_wdata), .clk(f434_clk), .rst(f434_rst), .rdata(f434_rdata));
  assign f434_clk = clk;
  assign f434_rst = rst;
  // Bindings to f434

  // f436
  logic [0:0] f436_wen;
  logic [31:0] f436_wdata;
  logic [0:0] f436_clk;
  logic [0:0] f436_rst;
  logic [31:0] f436_rdata;
  sr_buffer_32_1 f436(.wen(f436_wen), .wdata(f436_wdata), .clk(f436_clk), .rst(f436_rst), .rdata(f436_rdata));
  assign f436_clk = clk;
  assign f436_rst = rst;
  // Bindings to f436

  // f438
  logic [0:0] f438_wen;
  logic [31:0] f438_wdata;
  logic [0:0] f438_clk;
  logic [0:0] f438_rst;
  logic [31:0] f438_rdata;
  sr_buffer_32_1 f438(.wen(f438_wen), .wdata(f438_wdata), .clk(f438_clk), .rst(f438_rst), .rdata(f438_rdata));
  assign f438_clk = clk;
  assign f438_rst = rst;
  // Bindings to f438

  // f440
  logic [0:0] f440_wen;
  logic [31:0] f440_wdata;
  logic [0:0] f440_clk;
  logic [0:0] f440_rst;
  logic [31:0] f440_rdata;
  sr_buffer_32_1 f440(.wen(f440_wen), .wdata(f440_wdata), .clk(f440_clk), .rst(f440_rst), .rdata(f440_rdata));
  assign f440_clk = clk;
  assign f440_rst = rst;
  // Bindings to f440

  // f442
  logic [0:0] f442_wen;
  logic [31:0] f442_wdata;
  logic [0:0] f442_clk;
  logic [0:0] f442_rst;
  logic [31:0] f442_rdata;
  sr_buffer_32_1 f442(.wen(f442_wen), .wdata(f442_wdata), .clk(f442_clk), .rst(f442_rst), .rdata(f442_rdata));
  assign f442_clk = clk;
  assign f442_rst = rst;
  // Bindings to f442

  // f444
  logic [0:0] f444_wen;
  logic [31:0] f444_wdata;
  logic [0:0] f444_clk;
  logic [0:0] f444_rst;
  logic [31:0] f444_rdata;
  sr_buffer_32_1 f444(.wen(f444_wen), .wdata(f444_wdata), .clk(f444_clk), .rst(f444_rst), .rdata(f444_rdata));
  assign f444_clk = clk;
  assign f444_rst = rst;
  // Bindings to f444

  // f446
  logic [0:0] f446_wen;
  logic [31:0] f446_wdata;
  logic [0:0] f446_clk;
  logic [0:0] f446_rst;
  logic [31:0] f446_rdata;
  sr_buffer_32_1 f446(.wen(f446_wen), .wdata(f446_wdata), .clk(f446_clk), .rst(f446_rst), .rdata(f446_rdata));
  assign f446_clk = clk;
  assign f446_rst = rst;
  // Bindings to f446

  // f448
  logic [0:0] f448_wen;
  logic [31:0] f448_wdata;
  logic [0:0] f448_clk;
  logic [0:0] f448_rst;
  logic [31:0] f448_rdata;
  sr_buffer_32_1 f448(.wen(f448_wen), .wdata(f448_wdata), .clk(f448_clk), .rst(f448_rst), .rdata(f448_rdata));
  assign f448_clk = clk;
  assign f448_rst = rst;
  // Bindings to f448

  // f450
  logic [0:0] f450_wen;
  logic [31:0] f450_wdata;
  logic [0:0] f450_clk;
  logic [0:0] f450_rst;
  logic [31:0] f450_rdata;
  sr_buffer_32_1 f450(.wen(f450_wen), .wdata(f450_wdata), .clk(f450_clk), .rst(f450_rst), .rdata(f450_rdata));
  assign f450_clk = clk;
  assign f450_rst = rst;
  // Bindings to f450

  // f452
  logic [0:0] f452_wen;
  logic [31:0] f452_wdata;
  logic [0:0] f452_clk;
  logic [0:0] f452_rst;
  logic [31:0] f452_rdata;
  sr_buffer_32_1 f452(.wen(f452_wen), .wdata(f452_wdata), .clk(f452_clk), .rst(f452_rst), .rdata(f452_rdata));
  assign f452_clk = clk;
  assign f452_rst = rst;
  // Bindings to f452

  // f454
  logic [0:0] f454_wen;
  logic [31:0] f454_wdata;
  logic [0:0] f454_clk;
  logic [0:0] f454_rst;
  logic [31:0] f454_rdata;
  sr_buffer_32_1 f454(.wen(f454_wen), .wdata(f454_wdata), .clk(f454_clk), .rst(f454_rst), .rdata(f454_rdata));
  assign f454_clk = clk;
  assign f454_rst = rst;
  // Bindings to f454

  // f456
  logic [0:0] f456_wen;
  logic [31:0] f456_wdata;
  logic [0:0] f456_clk;
  logic [0:0] f456_rst;
  logic [31:0] f456_rdata;
  sr_buffer_32_1 f456(.wen(f456_wen), .wdata(f456_wdata), .clk(f456_clk), .rst(f456_rst), .rdata(f456_rdata));
  assign f456_clk = clk;
  assign f456_rst = rst;
  // Bindings to f456

  // f458
  logic [0:0] f458_wen;
  logic [31:0] f458_wdata;
  logic [0:0] f458_clk;
  logic [0:0] f458_rst;
  logic [31:0] f458_rdata;
  sr_buffer_32_1 f458(.wen(f458_wen), .wdata(f458_wdata), .clk(f458_clk), .rst(f458_rst), .rdata(f458_rdata));
  assign f458_clk = clk;
  assign f458_rst = rst;
  // Bindings to f458

  // f460
  logic [0:0] f460_wen;
  logic [31:0] f460_wdata;
  logic [0:0] f460_clk;
  logic [0:0] f460_rst;
  logic [31:0] f460_rdata;
  sr_buffer_32_1 f460(.wen(f460_wen), .wdata(f460_wdata), .clk(f460_clk), .rst(f460_rst), .rdata(f460_rdata));
  assign f460_clk = clk;
  assign f460_rst = rst;
  // Bindings to f460

  // f462
  logic [0:0] f462_wen;
  logic [31:0] f462_wdata;
  logic [0:0] f462_clk;
  logic [0:0] f462_rst;
  logic [31:0] f462_rdata;
  sr_buffer_32_1 f462(.wen(f462_wen), .wdata(f462_wdata), .clk(f462_clk), .rst(f462_rst), .rdata(f462_rdata));
  assign f462_clk = clk;
  assign f462_rst = rst;
  // Bindings to f462

  // f464
  logic [0:0] f464_wen;
  logic [31:0] f464_wdata;
  logic [0:0] f464_clk;
  logic [0:0] f464_rst;
  logic [31:0] f464_rdata;
  sr_buffer_32_1 f464(.wen(f464_wen), .wdata(f464_wdata), .clk(f464_clk), .rst(f464_rst), .rdata(f464_rdata));
  assign f464_clk = clk;
  assign f464_rst = rst;
  // Bindings to f464

  // f466
  logic [0:0] f466_wen;
  logic [31:0] f466_wdata;
  logic [0:0] f466_clk;
  logic [0:0] f466_rst;
  logic [31:0] f466_rdata;
  sr_buffer_32_1 f466(.wen(f466_wen), .wdata(f466_wdata), .clk(f466_clk), .rst(f466_rst), .rdata(f466_rdata));
  assign f466_clk = clk;
  assign f466_rst = rst;
  // Bindings to f466

  // f468
  logic [0:0] f468_wen;
  logic [31:0] f468_wdata;
  logic [0:0] f468_clk;
  logic [0:0] f468_rst;
  logic [31:0] f468_rdata;
  sr_buffer_32_1 f468(.wen(f468_wen), .wdata(f468_wdata), .clk(f468_clk), .rst(f468_rst), .rdata(f468_rdata));
  assign f468_clk = clk;
  assign f468_rst = rst;
  // Bindings to f468

  // f470
  logic [0:0] f470_wen;
  logic [31:0] f470_wdata;
  logic [0:0] f470_clk;
  logic [0:0] f470_rst;
  logic [31:0] f470_rdata;
  sr_buffer_32_1 f470(.wen(f470_wen), .wdata(f470_wdata), .clk(f470_clk), .rst(f470_rst), .rdata(f470_rdata));
  assign f470_clk = clk;
  assign f470_rst = rst;
  // Bindings to f470

  // f472
  logic [0:0] f472_wen;
  logic [31:0] f472_wdata;
  logic [0:0] f472_clk;
  logic [0:0] f472_rst;
  logic [31:0] f472_rdata;
  sr_buffer_32_1 f472(.wen(f472_wen), .wdata(f472_wdata), .clk(f472_clk), .rst(f472_rst), .rdata(f472_rdata));
  assign f472_clk = clk;
  assign f472_rst = rst;
  // Bindings to f472

  // f474
  logic [0:0] f474_wen;
  logic [31:0] f474_wdata;
  logic [0:0] f474_clk;
  logic [0:0] f474_rst;
  logic [31:0] f474_rdata;
  sr_buffer_32_1 f474(.wen(f474_wen), .wdata(f474_wdata), .clk(f474_clk), .rst(f474_rst), .rdata(f474_rdata));
  assign f474_clk = clk;
  assign f474_rst = rst;
  // Bindings to f474

  // f476
  logic [0:0] f476_wen;
  logic [31:0] f476_wdata;
  logic [0:0] f476_clk;
  logic [0:0] f476_rst;
  logic [31:0] f476_rdata;
  sr_buffer_32_1 f476(.wen(f476_wen), .wdata(f476_wdata), .clk(f476_clk), .rst(f476_rst), .rdata(f476_rdata));
  assign f476_clk = clk;
  assign f476_rst = rst;
  // Bindings to f476

  // f478
  logic [0:0] f478_wen;
  logic [31:0] f478_wdata;
  logic [0:0] f478_clk;
  logic [0:0] f478_rst;
  logic [31:0] f478_rdata;
  sr_buffer_32_1 f478(.wen(f478_wen), .wdata(f478_wdata), .clk(f478_clk), .rst(f478_rst), .rdata(f478_rdata));
  assign f478_clk = clk;
  assign f478_rst = rst;
  // Bindings to f478

  // f480
  logic [0:0] f480_wen;
  logic [31:0] f480_wdata;
  logic [0:0] f480_clk;
  logic [0:0] f480_rst;
  logic [31:0] f480_rdata;
  sr_buffer_32_1 f480(.wen(f480_wen), .wdata(f480_wdata), .clk(f480_clk), .rst(f480_rst), .rdata(f480_rdata));
  assign f480_clk = clk;
  assign f480_rst = rst;
  // Bindings to f480

  // f482
  logic [0:0] f482_wen;
  logic [31:0] f482_wdata;
  logic [0:0] f482_clk;
  logic [0:0] f482_rst;
  logic [31:0] f482_rdata;
  sr_buffer_32_1 f482(.wen(f482_wen), .wdata(f482_wdata), .clk(f482_clk), .rst(f482_rst), .rdata(f482_rdata));
  assign f482_clk = clk;
  assign f482_rst = rst;
  // Bindings to f482

  // f484
  logic [0:0] f484_wen;
  logic [31:0] f484_wdata;
  logic [0:0] f484_clk;
  logic [0:0] f484_rst;
  logic [31:0] f484_rdata;
  sr_buffer_32_1 f484(.wen(f484_wen), .wdata(f484_wdata), .clk(f484_clk), .rst(f484_rst), .rdata(f484_rdata));
  assign f484_clk = clk;
  assign f484_rst = rst;
  // Bindings to f484

  // f486
  logic [0:0] f486_wen;
  logic [31:0] f486_wdata;
  logic [0:0] f486_clk;
  logic [0:0] f486_rst;
  logic [31:0] f486_rdata;
  sr_buffer_32_1 f486(.wen(f486_wen), .wdata(f486_wdata), .clk(f486_clk), .rst(f486_rst), .rdata(f486_rdata));
  assign f486_clk = clk;
  assign f486_rst = rst;
  // Bindings to f486

  // f488
  logic [0:0] f488_wen;
  logic [31:0] f488_wdata;
  logic [0:0] f488_clk;
  logic [0:0] f488_rst;
  logic [31:0] f488_rdata;
  sr_buffer_32_1 f488(.wen(f488_wen), .wdata(f488_wdata), .clk(f488_clk), .rst(f488_rst), .rdata(f488_rdata));
  assign f488_clk = clk;
  assign f488_rst = rst;
  // Bindings to f488

  // f490
  logic [0:0] f490_wen;
  logic [31:0] f490_wdata;
  logic [0:0] f490_clk;
  logic [0:0] f490_rst;
  logic [31:0] f490_rdata;
  sr_buffer_32_1 f490(.wen(f490_wen), .wdata(f490_wdata), .clk(f490_clk), .rst(f490_rst), .rdata(f490_rdata));
  assign f490_clk = clk;
  assign f490_rst = rst;
  // Bindings to f490

  // f492
  logic [0:0] f492_wen;
  logic [31:0] f492_wdata;
  logic [0:0] f492_clk;
  logic [0:0] f492_rst;
  logic [31:0] f492_rdata;
  sr_buffer_32_1 f492(.wen(f492_wen), .wdata(f492_wdata), .clk(f492_clk), .rst(f492_rst), .rdata(f492_rdata));
  assign f492_clk = clk;
  assign f492_rst = rst;
  // Bindings to f492

  // f494
  logic [0:0] f494_wen;
  logic [31:0] f494_wdata;
  logic [0:0] f494_clk;
  logic [0:0] f494_rst;
  logic [31:0] f494_rdata;
  sr_buffer_32_1 f494(.wen(f494_wen), .wdata(f494_wdata), .clk(f494_clk), .rst(f494_rst), .rdata(f494_rdata));
  assign f494_clk = clk;
  assign f494_rst = rst;
  // Bindings to f494

  // f496
  logic [0:0] f496_wen;
  logic [31:0] f496_wdata;
  logic [0:0] f496_clk;
  logic [0:0] f496_rst;
  logic [31:0] f496_rdata;
  sr_buffer_32_1 f496(.wen(f496_wen), .wdata(f496_wdata), .clk(f496_clk), .rst(f496_rst), .rdata(f496_rdata));
  assign f496_clk = clk;
  assign f496_rst = rst;
  // Bindings to f496

  // f498
  logic [0:0] f498_wen;
  logic [31:0] f498_wdata;
  logic [0:0] f498_clk;
  logic [0:0] f498_rst;
  logic [31:0] f498_rdata;
  sr_buffer_32_1 f498(.wen(f498_wen), .wdata(f498_wdata), .clk(f498_clk), .rst(f498_rst), .rdata(f498_rdata));
  assign f498_clk = clk;
  assign f498_rst = rst;
  // Bindings to f498

  // f500
  logic [0:0] f500_wen;
  logic [31:0] f500_wdata;
  logic [0:0] f500_clk;
  logic [0:0] f500_rst;
  logic [31:0] f500_rdata;
  sr_buffer_32_1 f500(.wen(f500_wen), .wdata(f500_wdata), .clk(f500_clk), .rst(f500_rst), .rdata(f500_rdata));
  assign f500_clk = clk;
  assign f500_rst = rst;
  // Bindings to f500

  // f502
  logic [0:0] f502_wen;
  logic [31:0] f502_wdata;
  logic [0:0] f502_clk;
  logic [0:0] f502_rst;
  logic [31:0] f502_rdata;
  sr_buffer_32_1 f502(.wen(f502_wen), .wdata(f502_wdata), .clk(f502_clk), .rst(f502_rst), .rdata(f502_rdata));
  assign f502_clk = clk;
  assign f502_rst = rst;
  // Bindings to f502

  // f504
  logic [0:0] f504_wen;
  logic [31:0] f504_wdata;
  logic [0:0] f504_clk;
  logic [0:0] f504_rst;
  logic [31:0] f504_rdata;
  sr_buffer_32_1 f504(.wen(f504_wen), .wdata(f504_wdata), .clk(f504_clk), .rst(f504_rst), .rdata(f504_rdata));
  assign f504_clk = clk;
  assign f504_rst = rst;
  // Bindings to f504

  // f506
  logic [0:0] f506_wen;
  logic [31:0] f506_wdata;
  logic [0:0] f506_clk;
  logic [0:0] f506_rst;
  logic [31:0] f506_rdata;
  sr_buffer_32_1 f506(.wen(f506_wen), .wdata(f506_wdata), .clk(f506_clk), .rst(f506_rst), .rdata(f506_rdata));
  assign f506_clk = clk;
  assign f506_rst = rst;
  // Bindings to f506

  // f508
  logic [0:0] f508_wen;
  logic [31:0] f508_wdata;
  logic [0:0] f508_clk;
  logic [0:0] f508_rst;
  logic [31:0] f508_rdata;
  sr_buffer_32_1 f508(.wen(f508_wen), .wdata(f508_wdata), .clk(f508_clk), .rst(f508_rst), .rdata(f508_rdata));
  assign f508_clk = clk;
  assign f508_rst = rst;
  // Bindings to f508

  // f510
  logic [0:0] f510_wen;
  logic [31:0] f510_wdata;
  logic [0:0] f510_clk;
  logic [0:0] f510_rst;
  logic [31:0] f510_rdata;
  sr_buffer_32_1 f510(.wen(f510_wen), .wdata(f510_wdata), .clk(f510_clk), .rst(f510_rst), .rdata(f510_rdata));
  assign f510_clk = clk;
  assign f510_rst = rst;
  // Bindings to f510

  // f512
  logic [0:0] f512_wen;
  logic [31:0] f512_wdata;
  logic [0:0] f512_clk;
  logic [0:0] f512_rst;
  logic [31:0] f512_rdata;
  sr_buffer_32_1 f512(.wen(f512_wen), .wdata(f512_wdata), .clk(f512_clk), .rst(f512_rst), .rdata(f512_rdata));
  assign f512_clk = clk;
  assign f512_rst = rst;
  // Bindings to f512

  // f514
  logic [0:0] f514_wen;
  logic [31:0] f514_wdata;
  logic [0:0] f514_clk;
  logic [0:0] f514_rst;
  logic [31:0] f514_rdata;
  sr_buffer_32_1 f514(.wen(f514_wen), .wdata(f514_wdata), .clk(f514_clk), .rst(f514_rst), .rdata(f514_rdata));
  assign f514_clk = clk;
  assign f514_rst = rst;
  // Bindings to f514

  // f516
  logic [0:0] f516_wen;
  logic [31:0] f516_wdata;
  logic [0:0] f516_clk;
  logic [0:0] f516_rst;
  logic [31:0] f516_rdata;
  sr_buffer_32_1 f516(.wen(f516_wen), .wdata(f516_wdata), .clk(f516_clk), .rst(f516_rst), .rdata(f516_rdata));
  assign f516_clk = clk;
  assign f516_rst = rst;
  // Bindings to f516

  // f518
  logic [0:0] f518_wen;
  logic [31:0] f518_wdata;
  logic [0:0] f518_clk;
  logic [0:0] f518_rst;
  logic [31:0] f518_rdata;
  sr_buffer_32_1 f518(.wen(f518_wen), .wdata(f518_wdata), .clk(f518_clk), .rst(f518_rst), .rdata(f518_rdata));
  assign f518_clk = clk;
  assign f518_rst = rst;
  // Bindings to f518

  // f520
  logic [0:0] f520_wen;
  logic [31:0] f520_wdata;
  logic [0:0] f520_clk;
  logic [0:0] f520_rst;
  logic [31:0] f520_rdata;
  sr_buffer_32_1 f520(.wen(f520_wen), .wdata(f520_wdata), .clk(f520_clk), .rst(f520_rst), .rdata(f520_rdata));
  assign f520_clk = clk;
  assign f520_rst = rst;
  // Bindings to f520

  // f522
  logic [0:0] f522_wen;
  logic [31:0] f522_wdata;
  logic [0:0] f522_clk;
  logic [0:0] f522_rst;
  logic [31:0] f522_rdata;
  sr_buffer_32_1 f522(.wen(f522_wen), .wdata(f522_wdata), .clk(f522_clk), .rst(f522_rst), .rdata(f522_rdata));
  assign f522_clk = clk;
  assign f522_rst = rst;
  // Bindings to f522

  // f524
  logic [0:0] f524_wen;
  logic [31:0] f524_wdata;
  logic [0:0] f524_clk;
  logic [0:0] f524_rst;
  logic [31:0] f524_rdata;
  sr_buffer_32_1 f524(.wen(f524_wen), .wdata(f524_wdata), .clk(f524_clk), .rst(f524_rst), .rdata(f524_rdata));
  assign f524_clk = clk;
  assign f524_rst = rst;
  // Bindings to f524

  // f526
  logic [0:0] f526_wen;
  logic [31:0] f526_wdata;
  logic [0:0] f526_clk;
  logic [0:0] f526_rst;
  logic [31:0] f526_rdata;
  sr_buffer_32_1 f526(.wen(f526_wen), .wdata(f526_wdata), .clk(f526_clk), .rst(f526_rst), .rdata(f526_rdata));
  assign f526_clk = clk;
  assign f526_rst = rst;
  // Bindings to f526

  // f528
  logic [0:0] f528_wen;
  logic [31:0] f528_wdata;
  logic [0:0] f528_clk;
  logic [0:0] f528_rst;
  logic [31:0] f528_rdata;
  sr_buffer_32_1 f528(.wen(f528_wen), .wdata(f528_wdata), .clk(f528_clk), .rst(f528_rst), .rdata(f528_rdata));
  assign f528_clk = clk;
  assign f528_rst = rst;
  // Bindings to f528

  // f530
  logic [0:0] f530_wen;
  logic [31:0] f530_wdata;
  logic [0:0] f530_clk;
  logic [0:0] f530_rst;
  logic [31:0] f530_rdata;
  sr_buffer_32_1 f530(.wen(f530_wen), .wdata(f530_wdata), .clk(f530_clk), .rst(f530_rst), .rdata(f530_rdata));
  assign f530_clk = clk;
  assign f530_rst = rst;
  // Bindings to f530

  // f532
  logic [0:0] f532_wen;
  logic [31:0] f532_wdata;
  logic [0:0] f532_clk;
  logic [0:0] f532_rst;
  logic [31:0] f532_rdata;
  sr_buffer_32_1 f532(.wen(f532_wen), .wdata(f532_wdata), .clk(f532_clk), .rst(f532_rst), .rdata(f532_rdata));
  assign f532_clk = clk;
  assign f532_rst = rst;
  // Bindings to f532

  // f534
  logic [0:0] f534_wen;
  logic [31:0] f534_wdata;
  logic [0:0] f534_clk;
  logic [0:0] f534_rst;
  logic [31:0] f534_rdata;
  sr_buffer_32_1 f534(.wen(f534_wen), .wdata(f534_wdata), .clk(f534_clk), .rst(f534_rst), .rdata(f534_rdata));
  assign f534_clk = clk;
  assign f534_rst = rst;
  // Bindings to f534

  // f536
  logic [0:0] f536_wen;
  logic [31:0] f536_wdata;
  logic [0:0] f536_clk;
  logic [0:0] f536_rst;
  logic [31:0] f536_rdata;
  sr_buffer_32_1 f536(.wen(f536_wen), .wdata(f536_wdata), .clk(f536_clk), .rst(f536_rst), .rdata(f536_rdata));
  assign f536_clk = clk;
  assign f536_rst = rst;
  // Bindings to f536

  // f538
  logic [0:0] f538_wen;
  logic [31:0] f538_wdata;
  logic [0:0] f538_clk;
  logic [0:0] f538_rst;
  logic [31:0] f538_rdata;
  sr_buffer_32_1 f538(.wen(f538_wen), .wdata(f538_wdata), .clk(f538_clk), .rst(f538_rst), .rdata(f538_rdata));
  assign f538_clk = clk;
  assign f538_rst = rst;
  // Bindings to f538

  // f540
  logic [0:0] f540_wen;
  logic [31:0] f540_wdata;
  logic [0:0] f540_clk;
  logic [0:0] f540_rst;
  logic [31:0] f540_rdata;
  sr_buffer_32_1 f540(.wen(f540_wen), .wdata(f540_wdata), .clk(f540_clk), .rst(f540_rst), .rdata(f540_rdata));
  assign f540_clk = clk;
  assign f540_rst = rst;
  // Bindings to f540

  // f542
  logic [0:0] f542_wen;
  logic [31:0] f542_wdata;
  logic [0:0] f542_clk;
  logic [0:0] f542_rst;
  logic [31:0] f542_rdata;
  sr_buffer_32_1 f542(.wen(f542_wen), .wdata(f542_wdata), .clk(f542_clk), .rst(f542_rst), .rdata(f542_rdata));
  assign f542_clk = clk;
  assign f542_rst = rst;
  // Bindings to f542

  // f544
  logic [0:0] f544_wen;
  logic [31:0] f544_wdata;
  logic [0:0] f544_clk;
  logic [0:0] f544_rst;
  logic [31:0] f544_rdata;
  sr_buffer_32_1 f544(.wen(f544_wen), .wdata(f544_wdata), .clk(f544_clk), .rst(f544_rst), .rdata(f544_rdata));
  assign f544_clk = clk;
  assign f544_rst = rst;
  // Bindings to f544

  // f546
  logic [0:0] f546_wen;
  logic [31:0] f546_wdata;
  logic [0:0] f546_clk;
  logic [0:0] f546_rst;
  logic [31:0] f546_rdata;
  sr_buffer_32_1 f546(.wen(f546_wen), .wdata(f546_wdata), .clk(f546_clk), .rst(f546_rst), .rdata(f546_rdata));
  assign f546_clk = clk;
  assign f546_rst = rst;
  // Bindings to f546

  // f548
  logic [0:0] f548_wen;
  logic [31:0] f548_wdata;
  logic [0:0] f548_clk;
  logic [0:0] f548_rst;
  logic [31:0] f548_rdata;
  sr_buffer_32_1 f548(.wen(f548_wen), .wdata(f548_wdata), .clk(f548_clk), .rst(f548_rst), .rdata(f548_rdata));
  assign f548_clk = clk;
  assign f548_rst = rst;
  // Bindings to f548

  // f550
  logic [0:0] f550_wen;
  logic [31:0] f550_wdata;
  logic [0:0] f550_clk;
  logic [0:0] f550_rst;
  logic [31:0] f550_rdata;
  sr_buffer_32_1 f550(.wen(f550_wen), .wdata(f550_wdata), .clk(f550_clk), .rst(f550_rst), .rdata(f550_rdata));
  assign f550_clk = clk;
  assign f550_rst = rst;
  // Bindings to f550

  // f552
  logic [0:0] f552_wen;
  logic [31:0] f552_wdata;
  logic [0:0] f552_clk;
  logic [0:0] f552_rst;
  logic [31:0] f552_rdata;
  sr_buffer_32_1 f552(.wen(f552_wen), .wdata(f552_wdata), .clk(f552_clk), .rst(f552_rst), .rdata(f552_rdata));
  assign f552_clk = clk;
  assign f552_rst = rst;
  // Bindings to f552

  // f554
  logic [0:0] f554_wen;
  logic [31:0] f554_wdata;
  logic [0:0] f554_clk;
  logic [0:0] f554_rst;
  logic [31:0] f554_rdata;
  sr_buffer_32_1 f554(.wen(f554_wen), .wdata(f554_wdata), .clk(f554_clk), .rst(f554_rst), .rdata(f554_rdata));
  assign f554_clk = clk;
  assign f554_rst = rst;
  // Bindings to f554

  // f556
  logic [0:0] f556_wen;
  logic [31:0] f556_wdata;
  logic [0:0] f556_clk;
  logic [0:0] f556_rst;
  logic [31:0] f556_rdata;
  sr_buffer_32_1 f556(.wen(f556_wen), .wdata(f556_wdata), .clk(f556_clk), .rst(f556_rst), .rdata(f556_rdata));
  assign f556_clk = clk;
  assign f556_rst = rst;
  // Bindings to f556

  // f558
  logic [0:0] f558_wen;
  logic [31:0] f558_wdata;
  logic [0:0] f558_clk;
  logic [0:0] f558_rst;
  logic [31:0] f558_rdata;
  sr_buffer_32_1 f558(.wen(f558_wen), .wdata(f558_wdata), .clk(f558_clk), .rst(f558_rst), .rdata(f558_rdata));
  assign f558_clk = clk;
  assign f558_rst = rst;
  // Bindings to f558

  // f560
  logic [0:0] f560_wen;
  logic [31:0] f560_wdata;
  logic [0:0] f560_clk;
  logic [0:0] f560_rst;
  logic [31:0] f560_rdata;
  sr_buffer_32_1 f560(.wen(f560_wen), .wdata(f560_wdata), .clk(f560_clk), .rst(f560_rst), .rdata(f560_rdata));
  assign f560_clk = clk;
  assign f560_rst = rst;
  // Bindings to f560

  // f562
  logic [0:0] f562_wen;
  logic [31:0] f562_wdata;
  logic [0:0] f562_clk;
  logic [0:0] f562_rst;
  logic [31:0] f562_rdata;
  sr_buffer_32_1 f562(.wen(f562_wen), .wdata(f562_wdata), .clk(f562_clk), .rst(f562_rst), .rdata(f562_rdata));
  assign f562_clk = clk;
  assign f562_rst = rst;
  // Bindings to f562

  // f564
  logic [0:0] f564_wen;
  logic [31:0] f564_wdata;
  logic [0:0] f564_clk;
  logic [0:0] f564_rst;
  logic [31:0] f564_rdata;
  sr_buffer_32_1 f564(.wen(f564_wen), .wdata(f564_wdata), .clk(f564_clk), .rst(f564_rst), .rdata(f564_rdata));
  assign f564_clk = clk;
  assign f564_rst = rst;
  // Bindings to f564

  // f566
  logic [0:0] f566_wen;
  logic [31:0] f566_wdata;
  logic [0:0] f566_clk;
  logic [0:0] f566_rst;
  logic [31:0] f566_rdata;
  sr_buffer_32_1 f566(.wen(f566_wen), .wdata(f566_wdata), .clk(f566_clk), .rst(f566_rst), .rdata(f566_rdata));
  assign f566_clk = clk;
  assign f566_rst = rst;
  // Bindings to f566

  // f568
  logic [0:0] f568_wen;
  logic [31:0] f568_wdata;
  logic [0:0] f568_clk;
  logic [0:0] f568_rst;
  logic [31:0] f568_rdata;
  sr_buffer_32_1 f568(.wen(f568_wen), .wdata(f568_wdata), .clk(f568_clk), .rst(f568_rst), .rdata(f568_rdata));
  assign f568_clk = clk;
  assign f568_rst = rst;
  // Bindings to f568

  // f570
  logic [0:0] f570_wen;
  logic [31:0] f570_wdata;
  logic [0:0] f570_clk;
  logic [0:0] f570_rst;
  logic [31:0] f570_rdata;
  sr_buffer_32_1 f570(.wen(f570_wen), .wdata(f570_wdata), .clk(f570_clk), .rst(f570_rst), .rdata(f570_rdata));
  assign f570_clk = clk;
  assign f570_rst = rst;
  // Bindings to f570

  // f572
  logic [0:0] f572_wen;
  logic [31:0] f572_wdata;
  logic [0:0] f572_clk;
  logic [0:0] f572_rst;
  logic [31:0] f572_rdata;
  sr_buffer_32_1 f572(.wen(f572_wen), .wdata(f572_wdata), .clk(f572_clk), .rst(f572_rst), .rdata(f572_rdata));
  assign f572_clk = clk;
  assign f572_rst = rst;
  // Bindings to f572

  // f574
  logic [0:0] f574_wen;
  logic [31:0] f574_wdata;
  logic [0:0] f574_clk;
  logic [0:0] f574_rst;
  logic [31:0] f574_rdata;
  sr_buffer_32_1 f574(.wen(f574_wen), .wdata(f574_wdata), .clk(f574_clk), .rst(f574_rst), .rdata(f574_rdata));
  assign f574_clk = clk;
  assign f574_rst = rst;
  // Bindings to f574

  // f576
  logic [0:0] f576_wen;
  logic [31:0] f576_wdata;
  logic [0:0] f576_clk;
  logic [0:0] f576_rst;
  logic [31:0] f576_rdata;
  sr_buffer_32_1 f576(.wen(f576_wen), .wdata(f576_wdata), .clk(f576_clk), .rst(f576_rst), .rdata(f576_rdata));
  assign f576_clk = clk;
  assign f576_rst = rst;
  // Bindings to f576

  // f578
  logic [0:0] f578_wen;
  logic [31:0] f578_wdata;
  logic [0:0] f578_clk;
  logic [0:0] f578_rst;
  logic [31:0] f578_rdata;
  sr_buffer_32_1 f578(.wen(f578_wen), .wdata(f578_wdata), .clk(f578_clk), .rst(f578_rst), .rdata(f578_rdata));
  assign f578_clk = clk;
  assign f578_rst = rst;
  // Bindings to f578

  // f580
  logic [0:0] f580_wen;
  logic [31:0] f580_wdata;
  logic [0:0] f580_clk;
  logic [0:0] f580_rst;
  logic [31:0] f580_rdata;
  sr_buffer_32_1 f580(.wen(f580_wen), .wdata(f580_wdata), .clk(f580_clk), .rst(f580_rst), .rdata(f580_rdata));
  assign f580_clk = clk;
  assign f580_rst = rst;
  // Bindings to f580

  // f582
  logic [0:0] f582_wen;
  logic [31:0] f582_wdata;
  logic [0:0] f582_clk;
  logic [0:0] f582_rst;
  logic [31:0] f582_rdata;
  sr_buffer_32_1 f582(.wen(f582_wen), .wdata(f582_wdata), .clk(f582_clk), .rst(f582_rst), .rdata(f582_rdata));
  assign f582_clk = clk;
  assign f582_rst = rst;
  // Bindings to f582

  // f584
  logic [0:0] f584_wen;
  logic [31:0] f584_wdata;
  logic [0:0] f584_clk;
  logic [0:0] f584_rst;
  logic [31:0] f584_rdata;
  sr_buffer_32_1 f584(.wen(f584_wen), .wdata(f584_wdata), .clk(f584_clk), .rst(f584_rst), .rdata(f584_rdata));
  assign f584_clk = clk;
  assign f584_rst = rst;
  // Bindings to f584

  // f586
  logic [0:0] f586_wen;
  logic [31:0] f586_wdata;
  logic [0:0] f586_clk;
  logic [0:0] f586_rst;
  logic [31:0] f586_rdata;
  sr_buffer_32_1 f586(.wen(f586_wen), .wdata(f586_wdata), .clk(f586_clk), .rst(f586_rst), .rdata(f586_rdata));
  assign f586_clk = clk;
  assign f586_rst = rst;
  // Bindings to f586

  // f588
  logic [0:0] f588_wen;
  logic [31:0] f588_wdata;
  logic [0:0] f588_clk;
  logic [0:0] f588_rst;
  logic [31:0] f588_rdata;
  sr_buffer_32_1 f588(.wen(f588_wen), .wdata(f588_wdata), .clk(f588_clk), .rst(f588_rst), .rdata(f588_rdata));
  assign f588_clk = clk;
  assign f588_rst = rst;
  // Bindings to f588

  // f590
  logic [0:0] f590_wen;
  logic [31:0] f590_wdata;
  logic [0:0] f590_clk;
  logic [0:0] f590_rst;
  logic [31:0] f590_rdata;
  sr_buffer_32_1 f590(.wen(f590_wen), .wdata(f590_wdata), .clk(f590_clk), .rst(f590_rst), .rdata(f590_rdata));
  assign f590_clk = clk;
  assign f590_rst = rst;
  // Bindings to f590

  // f592
  logic [0:0] f592_wen;
  logic [31:0] f592_wdata;
  logic [0:0] f592_clk;
  logic [0:0] f592_rst;
  logic [31:0] f592_rdata;
  sr_buffer_32_1 f592(.wen(f592_wen), .wdata(f592_wdata), .clk(f592_clk), .rst(f592_rst), .rdata(f592_rdata));
  assign f592_clk = clk;
  assign f592_rst = rst;
  // Bindings to f592

  // f594
  logic [0:0] f594_wen;
  logic [31:0] f594_wdata;
  logic [0:0] f594_clk;
  logic [0:0] f594_rst;
  logic [31:0] f594_rdata;
  sr_buffer_32_1 f594(.wen(f594_wen), .wdata(f594_wdata), .clk(f594_clk), .rst(f594_rst), .rdata(f594_rdata));
  assign f594_clk = clk;
  assign f594_rst = rst;
  // Bindings to f594

  // f596
  logic [0:0] f596_wen;
  logic [31:0] f596_wdata;
  logic [0:0] f596_clk;
  logic [0:0] f596_rst;
  logic [31:0] f596_rdata;
  sr_buffer_32_1 f596(.wen(f596_wen), .wdata(f596_wdata), .clk(f596_clk), .rst(f596_rst), .rdata(f596_rdata));
  assign f596_clk = clk;
  assign f596_rst = rst;
  // Bindings to f596

  // f598
  logic [0:0] f598_wen;
  logic [31:0] f598_wdata;
  logic [0:0] f598_clk;
  logic [0:0] f598_rst;
  logic [31:0] f598_rdata;
  sr_buffer_32_1 f598(.wen(f598_wen), .wdata(f598_wdata), .clk(f598_clk), .rst(f598_rst), .rdata(f598_rdata));
  assign f598_clk = clk;
  assign f598_rst = rst;
  // Bindings to f598

  // f600
  logic [0:0] f600_wen;
  logic [31:0] f600_wdata;
  logic [0:0] f600_clk;
  logic [0:0] f600_rst;
  logic [31:0] f600_rdata;
  sr_buffer_32_1 f600(.wen(f600_wen), .wdata(f600_wdata), .clk(f600_clk), .rst(f600_rst), .rdata(f600_rdata));
  assign f600_clk = clk;
  assign f600_rst = rst;
  // Bindings to f600

  // f602
  logic [0:0] f602_wen;
  logic [31:0] f602_wdata;
  logic [0:0] f602_clk;
  logic [0:0] f602_rst;
  logic [31:0] f602_rdata;
  sr_buffer_32_1 f602(.wen(f602_wen), .wdata(f602_wdata), .clk(f602_clk), .rst(f602_rst), .rdata(f602_rdata));
  assign f602_clk = clk;
  assign f602_rst = rst;
  // Bindings to f602

  // f604
  logic [0:0] f604_wen;
  logic [31:0] f604_wdata;
  logic [0:0] f604_clk;
  logic [0:0] f604_rst;
  logic [31:0] f604_rdata;
  sr_buffer_32_1 f604(.wen(f604_wen), .wdata(f604_wdata), .clk(f604_clk), .rst(f604_rst), .rdata(f604_rdata));
  assign f604_clk = clk;
  assign f604_rst = rst;
  // Bindings to f604

  // f606
  logic [0:0] f606_wen;
  logic [31:0] f606_wdata;
  logic [0:0] f606_clk;
  logic [0:0] f606_rst;
  logic [31:0] f606_rdata;
  sr_buffer_32_1 f606(.wen(f606_wen), .wdata(f606_wdata), .clk(f606_clk), .rst(f606_rst), .rdata(f606_rdata));
  assign f606_clk = clk;
  assign f606_rst = rst;
  // Bindings to f606

  // f608
  logic [0:0] f608_wen;
  logic [31:0] f608_wdata;
  logic [0:0] f608_clk;
  logic [0:0] f608_rst;
  logic [31:0] f608_rdata;
  sr_buffer_32_1 f608(.wen(f608_wen), .wdata(f608_wdata), .clk(f608_clk), .rst(f608_rst), .rdata(f608_rdata));
  assign f608_clk = clk;
  assign f608_rst = rst;
  // Bindings to f608

  // f610
  logic [0:0] f610_wen;
  logic [31:0] f610_wdata;
  logic [0:0] f610_clk;
  logic [0:0] f610_rst;
  logic [31:0] f610_rdata;
  sr_buffer_32_1 f610(.wen(f610_wen), .wdata(f610_wdata), .clk(f610_clk), .rst(f610_rst), .rdata(f610_rdata));
  assign f610_clk = clk;
  assign f610_rst = rst;
  // Bindings to f610

  // f612
  logic [0:0] f612_wen;
  logic [31:0] f612_wdata;
  logic [0:0] f612_clk;
  logic [0:0] f612_rst;
  logic [31:0] f612_rdata;
  sr_buffer_32_1 f612(.wen(f612_wen), .wdata(f612_wdata), .clk(f612_clk), .rst(f612_rst), .rdata(f612_rdata));
  assign f612_clk = clk;
  assign f612_rst = rst;
  // Bindings to f612

  // f614
  logic [0:0] f614_wen;
  logic [31:0] f614_wdata;
  logic [0:0] f614_clk;
  logic [0:0] f614_rst;
  logic [31:0] f614_rdata;
  sr_buffer_32_1 f614(.wen(f614_wen), .wdata(f614_wdata), .clk(f614_clk), .rst(f614_rst), .rdata(f614_rdata));
  assign f614_clk = clk;
  assign f614_rst = rst;
  // Bindings to f614

  // f616
  logic [0:0] f616_wen;
  logic [31:0] f616_wdata;
  logic [0:0] f616_clk;
  logic [0:0] f616_rst;
  logic [31:0] f616_rdata;
  sr_buffer_32_1 f616(.wen(f616_wen), .wdata(f616_wdata), .clk(f616_clk), .rst(f616_rst), .rdata(f616_rdata));
  assign f616_clk = clk;
  assign f616_rst = rst;
  // Bindings to f616

  // f618
  logic [0:0] f618_wen;
  logic [31:0] f618_wdata;
  logic [0:0] f618_clk;
  logic [0:0] f618_rst;
  logic [31:0] f618_rdata;
  sr_buffer_32_1 f618(.wen(f618_wen), .wdata(f618_wdata), .clk(f618_clk), .rst(f618_rst), .rdata(f618_rdata));
  assign f618_clk = clk;
  assign f618_rst = rst;
  // Bindings to f618

  // f620
  logic [0:0] f620_wen;
  logic [31:0] f620_wdata;
  logic [0:0] f620_clk;
  logic [0:0] f620_rst;
  logic [31:0] f620_rdata;
  sr_buffer_32_1 f620(.wen(f620_wen), .wdata(f620_wdata), .clk(f620_clk), .rst(f620_rst), .rdata(f620_rdata));
  assign f620_clk = clk;
  assign f620_rst = rst;
  // Bindings to f620

  // f622
  logic [0:0] f622_wen;
  logic [31:0] f622_wdata;
  logic [0:0] f622_clk;
  logic [0:0] f622_rst;
  logic [31:0] f622_rdata;
  sr_buffer_32_1 f622(.wen(f622_wen), .wdata(f622_wdata), .clk(f622_clk), .rst(f622_rst), .rdata(f622_rdata));
  assign f622_clk = clk;
  assign f622_rst = rst;
  // Bindings to f622

  // f624
  logic [0:0] f624_wen;
  logic [31:0] f624_wdata;
  logic [0:0] f624_clk;
  logic [0:0] f624_rst;
  logic [31:0] f624_rdata;
  sr_buffer_32_1 f624(.wen(f624_wen), .wdata(f624_wdata), .clk(f624_clk), .rst(f624_rst), .rdata(f624_rdata));
  assign f624_clk = clk;
  assign f624_rst = rst;
  // Bindings to f624

  // f626
  logic [0:0] f626_wen;
  logic [31:0] f626_wdata;
  logic [0:0] f626_clk;
  logic [0:0] f626_rst;
  logic [31:0] f626_rdata;
  sr_buffer_32_1 f626(.wen(f626_wen), .wdata(f626_wdata), .clk(f626_clk), .rst(f626_rst), .rdata(f626_rdata));
  assign f626_clk = clk;
  assign f626_rst = rst;
  // Bindings to f626

  // f628
  logic [0:0] f628_wen;
  logic [31:0] f628_wdata;
  logic [0:0] f628_clk;
  logic [0:0] f628_rst;
  logic [31:0] f628_rdata;
  sr_buffer_32_1 f628(.wen(f628_wen), .wdata(f628_wdata), .clk(f628_clk), .rst(f628_rst), .rdata(f628_rdata));
  assign f628_clk = clk;
  assign f628_rst = rst;
  // Bindings to f628

  // f630
  logic [0:0] f630_wen;
  logic [31:0] f630_wdata;
  logic [0:0] f630_clk;
  logic [0:0] f630_rst;
  logic [31:0] f630_rdata;
  sr_buffer_32_1 f630(.wen(f630_wen), .wdata(f630_wdata), .clk(f630_clk), .rst(f630_rst), .rdata(f630_rdata));
  assign f630_clk = clk;
  assign f630_rst = rst;
  // Bindings to f630

  // f632
  logic [0:0] f632_wen;
  logic [31:0] f632_wdata;
  logic [0:0] f632_clk;
  logic [0:0] f632_rst;
  logic [31:0] f632_rdata;
  sr_buffer_32_1 f632(.wen(f632_wen), .wdata(f632_wdata), .clk(f632_clk), .rst(f632_rst), .rdata(f632_rdata));
  assign f632_clk = clk;
  assign f632_rst = rst;
  // Bindings to f632

  // f634
  logic [0:0] f634_wen;
  logic [31:0] f634_wdata;
  logic [0:0] f634_clk;
  logic [0:0] f634_rst;
  logic [31:0] f634_rdata;
  sr_buffer_32_1 f634(.wen(f634_wen), .wdata(f634_wdata), .clk(f634_clk), .rst(f634_rst), .rdata(f634_rdata));
  assign f634_clk = clk;
  assign f634_rst = rst;
  // Bindings to f634

  // f636
  logic [0:0] f636_wen;
  logic [31:0] f636_wdata;
  logic [0:0] f636_clk;
  logic [0:0] f636_rst;
  logic [31:0] f636_rdata;
  sr_buffer_32_1 f636(.wen(f636_wen), .wdata(f636_wdata), .clk(f636_clk), .rst(f636_rst), .rdata(f636_rdata));
  assign f636_clk = clk;
  assign f636_rst = rst;
  // Bindings to f636

  // f638
  logic [0:0] f638_wen;
  logic [31:0] f638_wdata;
  logic [0:0] f638_clk;
  logic [0:0] f638_rst;
  logic [31:0] f638_rdata;
  sr_buffer_32_1 f638(.wen(f638_wen), .wdata(f638_wdata), .clk(f638_clk), .rst(f638_rst), .rdata(f638_rdata));
  assign f638_clk = clk;
  assign f638_rst = rst;
  // Bindings to f638

  // f640
  logic [0:0] f640_wen;
  logic [31:0] f640_wdata;
  logic [0:0] f640_clk;
  logic [0:0] f640_rst;
  logic [31:0] f640_rdata;
  sr_buffer_32_1 f640(.wen(f640_wen), .wdata(f640_wdata), .clk(f640_clk), .rst(f640_rst), .rdata(f640_rdata));
  assign f640_clk = clk;
  assign f640_rst = rst;
  // Bindings to f640

  // f642
  logic [0:0] f642_wen;
  logic [31:0] f642_wdata;
  logic [0:0] f642_clk;
  logic [0:0] f642_rst;
  logic [31:0] f642_rdata;
  sr_buffer_32_1 f642(.wen(f642_wen), .wdata(f642_wdata), .clk(f642_clk), .rst(f642_rst), .rdata(f642_rdata));
  assign f642_clk = clk;
  assign f642_rst = rst;
  // Bindings to f642

  // f644
  logic [0:0] f644_wen;
  logic [31:0] f644_wdata;
  logic [0:0] f644_clk;
  logic [0:0] f644_rst;
  logic [31:0] f644_rdata;
  sr_buffer_32_1 f644(.wen(f644_wen), .wdata(f644_wdata), .clk(f644_clk), .rst(f644_rst), .rdata(f644_rdata));
  assign f644_clk = clk;
  assign f644_rst = rst;
  // Bindings to f644

  // f646
  logic [0:0] f646_wen;
  logic [31:0] f646_wdata;
  logic [0:0] f646_clk;
  logic [0:0] f646_rst;
  logic [31:0] f646_rdata;
  sr_buffer_32_1 f646(.wen(f646_wen), .wdata(f646_wdata), .clk(f646_clk), .rst(f646_rst), .rdata(f646_rdata));
  assign f646_clk = clk;
  assign f646_rst = rst;
  // Bindings to f646

  // f648
  logic [0:0] f648_wen;
  logic [31:0] f648_wdata;
  logic [0:0] f648_clk;
  logic [0:0] f648_rst;
  logic [31:0] f648_rdata;
  sr_buffer_32_1 f648(.wen(f648_wen), .wdata(f648_wdata), .clk(f648_clk), .rst(f648_rst), .rdata(f648_rdata));
  assign f648_clk = clk;
  assign f648_rst = rst;
  // Bindings to f648

  // f650
  logic [0:0] f650_wen;
  logic [31:0] f650_wdata;
  logic [0:0] f650_clk;
  logic [0:0] f650_rst;
  logic [31:0] f650_rdata;
  sr_buffer_32_1 f650(.wen(f650_wen), .wdata(f650_wdata), .clk(f650_clk), .rst(f650_rst), .rdata(f650_rdata));
  assign f650_clk = clk;
  assign f650_rst = rst;
  // Bindings to f650

  // f652
  logic [0:0] f652_wen;
  logic [31:0] f652_wdata;
  logic [0:0] f652_clk;
  logic [0:0] f652_rst;
  logic [31:0] f652_rdata;
  sr_buffer_32_1 f652(.wen(f652_wen), .wdata(f652_wdata), .clk(f652_clk), .rst(f652_rst), .rdata(f652_rdata));
  assign f652_clk = clk;
  assign f652_rst = rst;
  // Bindings to f652

  // f654
  logic [0:0] f654_wen;
  logic [31:0] f654_wdata;
  logic [0:0] f654_clk;
  logic [0:0] f654_rst;
  logic [31:0] f654_rdata;
  sr_buffer_32_1 f654(.wen(f654_wen), .wdata(f654_wdata), .clk(f654_clk), .rst(f654_rst), .rdata(f654_rdata));
  assign f654_clk = clk;
  assign f654_rst = rst;
  // Bindings to f654

  // f656
  logic [0:0] f656_wen;
  logic [31:0] f656_wdata;
  logic [0:0] f656_clk;
  logic [0:0] f656_rst;
  logic [31:0] f656_rdata;
  sr_buffer_32_1 f656(.wen(f656_wen), .wdata(f656_wdata), .clk(f656_clk), .rst(f656_rst), .rdata(f656_rdata));
  assign f656_clk = clk;
  assign f656_rst = rst;
  // Bindings to f656

  // f658
  logic [0:0] f658_wen;
  logic [31:0] f658_wdata;
  logic [0:0] f658_clk;
  logic [0:0] f658_rst;
  logic [31:0] f658_rdata;
  sr_buffer_32_1 f658(.wen(f658_wen), .wdata(f658_wdata), .clk(f658_clk), .rst(f658_rst), .rdata(f658_rdata));
  assign f658_clk = clk;
  assign f658_rst = rst;
  // Bindings to f658

  // f660
  logic [0:0] f660_wen;
  logic [31:0] f660_wdata;
  logic [0:0] f660_clk;
  logic [0:0] f660_rst;
  logic [31:0] f660_rdata;
  sr_buffer_32_1 f660(.wen(f660_wen), .wdata(f660_wdata), .clk(f660_clk), .rst(f660_rst), .rdata(f660_rdata));
  assign f660_clk = clk;
  assign f660_rst = rst;
  // Bindings to f660

  // f662
  logic [0:0] f662_wen;
  logic [31:0] f662_wdata;
  logic [0:0] f662_clk;
  logic [0:0] f662_rst;
  logic [31:0] f662_rdata;
  sr_buffer_32_1 f662(.wen(f662_wen), .wdata(f662_wdata), .clk(f662_clk), .rst(f662_rst), .rdata(f662_rdata));
  assign f662_clk = clk;
  assign f662_rst = rst;
  // Bindings to f662

  // f664
  logic [0:0] f664_wen;
  logic [31:0] f664_wdata;
  logic [0:0] f664_clk;
  logic [0:0] f664_rst;
  logic [31:0] f664_rdata;
  sr_buffer_32_1 f664(.wen(f664_wen), .wdata(f664_wdata), .clk(f664_clk), .rst(f664_rst), .rdata(f664_rdata));
  assign f664_clk = clk;
  assign f664_rst = rst;
  // Bindings to f664

  // f666
  logic [0:0] f666_wen;
  logic [31:0] f666_wdata;
  logic [0:0] f666_clk;
  logic [0:0] f666_rst;
  logic [31:0] f666_rdata;
  sr_buffer_32_1 f666(.wen(f666_wen), .wdata(f666_wdata), .clk(f666_clk), .rst(f666_rst), .rdata(f666_rdata));
  assign f666_clk = clk;
  assign f666_rst = rst;
  // Bindings to f666

  // f668
  logic [0:0] f668_wen;
  logic [31:0] f668_wdata;
  logic [0:0] f668_clk;
  logic [0:0] f668_rst;
  logic [31:0] f668_rdata;
  sr_buffer_32_1 f668(.wen(f668_wen), .wdata(f668_wdata), .clk(f668_clk), .rst(f668_rst), .rdata(f668_rdata));
  assign f668_clk = clk;
  assign f668_rst = rst;
  // Bindings to f668

  // f670
  logic [0:0] f670_wen;
  logic [31:0] f670_wdata;
  logic [0:0] f670_clk;
  logic [0:0] f670_rst;
  logic [31:0] f670_rdata;
  sr_buffer_32_1 f670(.wen(f670_wen), .wdata(f670_wdata), .clk(f670_clk), .rst(f670_rst), .rdata(f670_rdata));
  assign f670_clk = clk;
  assign f670_rst = rst;
  // Bindings to f670

  // f672
  logic [0:0] f672_wen;
  logic [31:0] f672_wdata;
  logic [0:0] f672_clk;
  logic [0:0] f672_rst;
  logic [31:0] f672_rdata;
  sr_buffer_32_1 f672(.wen(f672_wen), .wdata(f672_wdata), .clk(f672_clk), .rst(f672_rst), .rdata(f672_rdata));
  assign f672_clk = clk;
  assign f672_rst = rst;
  // Bindings to f672

  // f674
  logic [0:0] f674_wen;
  logic [31:0] f674_wdata;
  logic [0:0] f674_clk;
  logic [0:0] f674_rst;
  logic [31:0] f674_rdata;
  sr_buffer_32_1 f674(.wen(f674_wen), .wdata(f674_wdata), .clk(f674_clk), .rst(f674_rst), .rdata(f674_rdata));
  assign f674_clk = clk;
  assign f674_rst = rst;
  // Bindings to f674

  // f676
  logic [0:0] f676_wen;
  logic [31:0] f676_wdata;
  logic [0:0] f676_clk;
  logic [0:0] f676_rst;
  logic [31:0] f676_rdata;
  sr_buffer_32_1 f676(.wen(f676_wen), .wdata(f676_wdata), .clk(f676_clk), .rst(f676_rst), .rdata(f676_rdata));
  assign f676_clk = clk;
  assign f676_rst = rst;
  // Bindings to f676

  // f678
  logic [0:0] f678_wen;
  logic [31:0] f678_wdata;
  logic [0:0] f678_clk;
  logic [0:0] f678_rst;
  logic [31:0] f678_rdata;
  sr_buffer_32_1 f678(.wen(f678_wen), .wdata(f678_wdata), .clk(f678_clk), .rst(f678_rst), .rdata(f678_rdata));
  assign f678_clk = clk;
  assign f678_rst = rst;
  // Bindings to f678

  // f680
  logic [0:0] f680_wen;
  logic [31:0] f680_wdata;
  logic [0:0] f680_clk;
  logic [0:0] f680_rst;
  logic [31:0] f680_rdata;
  sr_buffer_32_1 f680(.wen(f680_wen), .wdata(f680_wdata), .clk(f680_clk), .rst(f680_rst), .rdata(f680_rdata));
  assign f680_clk = clk;
  assign f680_rst = rst;
  // Bindings to f680

  // f682
  logic [0:0] f682_wen;
  logic [31:0] f682_wdata;
  logic [0:0] f682_clk;
  logic [0:0] f682_rst;
  logic [31:0] f682_rdata;
  sr_buffer_32_1 f682(.wen(f682_wen), .wdata(f682_wdata), .clk(f682_clk), .rst(f682_rst), .rdata(f682_rdata));
  assign f682_clk = clk;
  assign f682_rst = rst;
  // Bindings to f682

  // f684
  logic [0:0] f684_wen;
  logic [31:0] f684_wdata;
  logic [0:0] f684_clk;
  logic [0:0] f684_rst;
  logic [31:0] f684_rdata;
  sr_buffer_32_1 f684(.wen(f684_wen), .wdata(f684_wdata), .clk(f684_clk), .rst(f684_rst), .rdata(f684_rdata));
  assign f684_clk = clk;
  assign f684_rst = rst;
  // Bindings to f684

  // f686
  logic [0:0] f686_wen;
  logic [31:0] f686_wdata;
  logic [0:0] f686_clk;
  logic [0:0] f686_rst;
  logic [31:0] f686_rdata;
  sr_buffer_32_1 f686(.wen(f686_wen), .wdata(f686_wdata), .clk(f686_clk), .rst(f686_rst), .rdata(f686_rdata));
  assign f686_clk = clk;
  assign f686_rst = rst;
  // Bindings to f686

  // f688
  logic [0:0] f688_wen;
  logic [31:0] f688_wdata;
  logic [0:0] f688_clk;
  logic [0:0] f688_rst;
  logic [31:0] f688_rdata;
  sr_buffer_32_1 f688(.wen(f688_wen), .wdata(f688_wdata), .clk(f688_clk), .rst(f688_rst), .rdata(f688_rdata));
  assign f688_clk = clk;
  assign f688_rst = rst;
  // Bindings to f688

  // f690
  logic [0:0] f690_wen;
  logic [31:0] f690_wdata;
  logic [0:0] f690_clk;
  logic [0:0] f690_rst;
  logic [31:0] f690_rdata;
  sr_buffer_32_1 f690(.wen(f690_wen), .wdata(f690_wdata), .clk(f690_clk), .rst(f690_rst), .rdata(f690_rdata));
  assign f690_clk = clk;
  assign f690_rst = rst;
  // Bindings to f690

  // f692
  logic [0:0] f692_wen;
  logic [31:0] f692_wdata;
  logic [0:0] f692_clk;
  logic [0:0] f692_rst;
  logic [31:0] f692_rdata;
  sr_buffer_32_1 f692(.wen(f692_wen), .wdata(f692_wdata), .clk(f692_clk), .rst(f692_rst), .rdata(f692_rdata));
  assign f692_clk = clk;
  assign f692_rst = rst;
  // Bindings to f692

  // f694
  logic [0:0] f694_wen;
  logic [31:0] f694_wdata;
  logic [0:0] f694_clk;
  logic [0:0] f694_rst;
  logic [31:0] f694_rdata;
  sr_buffer_32_1 f694(.wen(f694_wen), .wdata(f694_wdata), .clk(f694_clk), .rst(f694_rst), .rdata(f694_rdata));
  assign f694_clk = clk;
  assign f694_rst = rst;
  // Bindings to f694

  // f696
  logic [0:0] f696_wen;
  logic [31:0] f696_wdata;
  logic [0:0] f696_clk;
  logic [0:0] f696_rst;
  logic [31:0] f696_rdata;
  sr_buffer_32_1 f696(.wen(f696_wen), .wdata(f696_wdata), .clk(f696_clk), .rst(f696_rst), .rdata(f696_rdata));
  assign f696_clk = clk;
  assign f696_rst = rst;
  // Bindings to f696

  // f698
  logic [0:0] f698_wen;
  logic [31:0] f698_wdata;
  logic [0:0] f698_clk;
  logic [0:0] f698_rst;
  logic [31:0] f698_rdata;
  sr_buffer_32_1 f698(.wen(f698_wen), .wdata(f698_wdata), .clk(f698_clk), .rst(f698_rst), .rdata(f698_rdata));
  assign f698_clk = clk;
  assign f698_rst = rst;
  // Bindings to f698

  // f700
  logic [0:0] f700_wen;
  logic [31:0] f700_wdata;
  logic [0:0] f700_clk;
  logic [0:0] f700_rst;
  logic [31:0] f700_rdata;
  sr_buffer_32_1 f700(.wen(f700_wen), .wdata(f700_wdata), .clk(f700_clk), .rst(f700_rst), .rdata(f700_rdata));
  assign f700_clk = clk;
  assign f700_rst = rst;
  // Bindings to f700

  // f702
  logic [0:0] f702_wen;
  logic [31:0] f702_wdata;
  logic [0:0] f702_clk;
  logic [0:0] f702_rst;
  logic [31:0] f702_rdata;
  sr_buffer_32_1 f702(.wen(f702_wen), .wdata(f702_wdata), .clk(f702_clk), .rst(f702_rst), .rdata(f702_rdata));
  assign f702_clk = clk;
  assign f702_rst = rst;
  // Bindings to f702

  // f704
  logic [0:0] f704_wen;
  logic [31:0] f704_wdata;
  logic [0:0] f704_clk;
  logic [0:0] f704_rst;
  logic [31:0] f704_rdata;
  sr_buffer_32_1 f704(.wen(f704_wen), .wdata(f704_wdata), .clk(f704_clk), .rst(f704_rst), .rdata(f704_rdata));
  assign f704_clk = clk;
  assign f704_rst = rst;
  // Bindings to f704

  // f706
  logic [0:0] f706_wen;
  logic [31:0] f706_wdata;
  logic [0:0] f706_clk;
  logic [0:0] f706_rst;
  logic [31:0] f706_rdata;
  sr_buffer_32_1 f706(.wen(f706_wen), .wdata(f706_wdata), .clk(f706_clk), .rst(f706_rst), .rdata(f706_rdata));
  assign f706_clk = clk;
  assign f706_rst = rst;
  // Bindings to f706

  // f804
  logic [0:0] f804_wen;
  logic [31:0] f804_wdata;
  logic [0:0] f804_clk;
  logic [0:0] f804_rst;
  logic [31:0] f804_rdata;
  sr_buffer_32_1 f804(.wen(f804_wen), .wdata(f804_wdata), .clk(f804_clk), .rst(f804_rst), .rdata(f804_rdata));
  assign f804_clk = clk;
  assign f804_rst = rst;
  // Bindings to f804

  // f838
  logic [0:0] f838_wen;
  logic [31:0] f838_wdata;
  logic [0:0] f838_clk;
  logic [0:0] f838_rst;
  logic [31:0] f838_rdata;
  sr_buffer_32_1 f838(.wen(f838_wen), .wdata(f838_wdata), .clk(f838_clk), .rst(f838_rst), .rdata(f838_rdata));
  assign f838_clk = clk;
  assign f838_rst = rst;
  // Bindings to f838

  // f940
  logic [0:0] f940_wen;
  logic [31:0] f940_wdata;
  logic [0:0] f940_clk;
  logic [0:0] f940_rst;
  logic [31:0] f940_rdata;
  sr_buffer_32_1 f940(.wen(f940_wen), .wdata(f940_wdata), .clk(f940_clk), .rst(f940_rst), .rdata(f940_rdata));
  assign f940_clk = clk;
  assign f940_rst = rst;
  // Bindings to f940

  // f942
  logic [0:0] f942_wen;
  logic [31:0] f942_wdata;
  logic [0:0] f942_clk;
  logic [0:0] f942_rst;
  logic [31:0] f942_rdata;
  sr_buffer_32_1 f942(.wen(f942_wen), .wdata(f942_wdata), .clk(f942_clk), .rst(f942_rst), .rdata(f942_rdata));
  assign f942_clk = clk;
  assign f942_rst = rst;
  // Bindings to f942

  // f944
  logic [0:0] f944_wen;
  logic [31:0] f944_wdata;
  logic [0:0] f944_clk;
  logic [0:0] f944_rst;
  logic [31:0] f944_rdata;
  sr_buffer_32_1 f944(.wen(f944_wen), .wdata(f944_wdata), .clk(f944_clk), .rst(f944_rst), .rdata(f944_rdata));
  assign f944_clk = clk;
  assign f944_rst = rst;
  // Bindings to f944

  // f946
  logic [0:0] f946_wen;
  logic [31:0] f946_wdata;
  logic [0:0] f946_clk;
  logic [0:0] f946_rst;
  logic [31:0] f946_rdata;
  sr_buffer_32_1 f946(.wen(f946_wen), .wdata(f946_wdata), .clk(f946_clk), .rst(f946_rst), .rdata(f946_rdata));
  assign f946_clk = clk;
  assign f946_rst = rst;
  // Bindings to f946

  // f948
  logic [0:0] f948_wen;
  logic [31:0] f948_wdata;
  logic [0:0] f948_clk;
  logic [0:0] f948_rst;
  logic [31:0] f948_rdata;
  sr_buffer_32_1 f948(.wen(f948_wen), .wdata(f948_wdata), .clk(f948_clk), .rst(f948_rst), .rdata(f948_rdata));
  assign f948_clk = clk;
  assign f948_rst = rst;
  // Bindings to f948

  // f950
  logic [0:0] f950_wen;
  logic [31:0] f950_wdata;
  logic [0:0] f950_clk;
  logic [0:0] f950_rst;
  logic [31:0] f950_rdata;
  sr_buffer_32_1 f950(.wen(f950_wen), .wdata(f950_wdata), .clk(f950_clk), .rst(f950_rst), .rdata(f950_rdata));
  assign f950_clk = clk;
  assign f950_rst = rst;
  // Bindings to f950

  // f952
  logic [0:0] f952_wen;
  logic [31:0] f952_wdata;
  logic [0:0] f952_clk;
  logic [0:0] f952_rst;
  logic [31:0] f952_rdata;
  sr_buffer_32_1 f952(.wen(f952_wen), .wdata(f952_wdata), .clk(f952_clk), .rst(f952_rst), .rdata(f952_rdata));
  assign f952_clk = clk;
  assign f952_rst = rst;
  // Bindings to f952

  // f954
  logic [0:0] f954_wen;
  logic [31:0] f954_wdata;
  logic [0:0] f954_clk;
  logic [0:0] f954_rst;
  logic [31:0] f954_rdata;
  sr_buffer_32_1 f954(.wen(f954_wen), .wdata(f954_wdata), .clk(f954_clk), .rst(f954_rst), .rdata(f954_rdata));
  assign f954_clk = clk;
  assign f954_rst = rst;
  // Bindings to f954

  // f956
  logic [0:0] f956_wen;
  logic [31:0] f956_wdata;
  logic [0:0] f956_clk;
  logic [0:0] f956_rst;
  logic [31:0] f956_rdata;
  sr_buffer_32_1 f956(.wen(f956_wen), .wdata(f956_wdata), .clk(f956_clk), .rst(f956_rst), .rdata(f956_rdata));
  assign f956_clk = clk;
  assign f956_rst = rst;
  // Bindings to f956

  // f958
  logic [0:0] f958_wen;
  logic [31:0] f958_wdata;
  logic [0:0] f958_clk;
  logic [0:0] f958_rst;
  logic [31:0] f958_rdata;
  sr_buffer_32_1 f958(.wen(f958_wen), .wdata(f958_wdata), .clk(f958_clk), .rst(f958_rst), .rdata(f958_rdata));
  assign f958_clk = clk;
  assign f958_rst = rst;
  // Bindings to f958

  // f960
  logic [0:0] f960_wen;
  logic [31:0] f960_wdata;
  logic [0:0] f960_clk;
  logic [0:0] f960_rst;
  logic [31:0] f960_rdata;
  sr_buffer_32_1 f960(.wen(f960_wen), .wdata(f960_wdata), .clk(f960_clk), .rst(f960_rst), .rdata(f960_rdata));
  assign f960_clk = clk;
  assign f960_rst = rst;
  // Bindings to f960

  // f962
  logic [0:0] f962_wen;
  logic [31:0] f962_wdata;
  logic [0:0] f962_clk;
  logic [0:0] f962_rst;
  logic [31:0] f962_rdata;
  sr_buffer_32_1 f962(.wen(f962_wen), .wdata(f962_wdata), .clk(f962_clk), .rst(f962_rst), .rdata(f962_rdata));
  assign f962_clk = clk;
  assign f962_rst = rst;
  // Bindings to f962

  // f964
  logic [0:0] f964_wen;
  logic [31:0] f964_wdata;
  logic [0:0] f964_clk;
  logic [0:0] f964_rst;
  logic [31:0] f964_rdata;
  sr_buffer_32_1 f964(.wen(f964_wen), .wdata(f964_wdata), .clk(f964_clk), .rst(f964_rst), .rdata(f964_rdata));
  assign f964_clk = clk;
  assign f964_rst = rst;
  // Bindings to f964

  // f966
  logic [0:0] f966_wen;
  logic [31:0] f966_wdata;
  logic [0:0] f966_clk;
  logic [0:0] f966_rst;
  logic [31:0] f966_rdata;
  sr_buffer_32_1 f966(.wen(f966_wen), .wdata(f966_wdata), .clk(f966_clk), .rst(f966_rst), .rdata(f966_rdata));
  assign f966_clk = clk;
  assign f966_rst = rst;
  // Bindings to f966

  // f968
  logic [0:0] f968_wen;
  logic [31:0] f968_wdata;
  logic [0:0] f968_clk;
  logic [0:0] f968_rst;
  logic [31:0] f968_rdata;
  sr_buffer_32_1 f968(.wen(f968_wen), .wdata(f968_wdata), .clk(f968_clk), .rst(f968_rst), .rdata(f968_rdata));
  assign f968_clk = clk;
  assign f968_rst = rst;
  // Bindings to f968

  // f970
  logic [0:0] f970_wen;
  logic [31:0] f970_wdata;
  logic [0:0] f970_clk;
  logic [0:0] f970_rst;
  logic [31:0] f970_rdata;
  sr_buffer_32_1 f970(.wen(f970_wen), .wdata(f970_wdata), .clk(f970_clk), .rst(f970_rst), .rdata(f970_rdata));
  assign f970_clk = clk;
  assign f970_rst = rst;
  // Bindings to f970

  // f972
  logic [0:0] f972_wen;
  logic [31:0] f972_wdata;
  logic [0:0] f972_clk;
  logic [0:0] f972_rst;
  logic [31:0] f972_rdata;
  sr_buffer_32_1 f972(.wen(f972_wen), .wdata(f972_wdata), .clk(f972_clk), .rst(f972_rst), .rdata(f972_rdata));
  assign f972_clk = clk;
  assign f972_rst = rst;
  // Bindings to f972

  // f974
  logic [0:0] f974_wen;
  logic [31:0] f974_wdata;
  logic [0:0] f974_clk;
  logic [0:0] f974_rst;
  logic [31:0] f974_rdata;
  sr_buffer_32_1 f974(.wen(f974_wen), .wdata(f974_wdata), .clk(f974_clk), .rst(f974_rst), .rdata(f974_rdata));
  assign f974_clk = clk;
  assign f974_rst = rst;
  // Bindings to f974

  // f976
  logic [0:0] f976_wen;
  logic [31:0] f976_wdata;
  logic [0:0] f976_clk;
  logic [0:0] f976_rst;
  logic [31:0] f976_rdata;
  sr_buffer_32_1 f976(.wen(f976_wen), .wdata(f976_wdata), .clk(f976_clk), .rst(f976_rst), .rdata(f976_rdata));
  assign f976_clk = clk;
  assign f976_rst = rst;
  // Bindings to f976

  // f978
  logic [0:0] f978_wen;
  logic [31:0] f978_wdata;
  logic [0:0] f978_clk;
  logic [0:0] f978_rst;
  logic [31:0] f978_rdata;
  sr_buffer_32_1 f978(.wen(f978_wen), .wdata(f978_wdata), .clk(f978_clk), .rst(f978_rst), .rdata(f978_rdata));
  assign f978_clk = clk;
  assign f978_rst = rst;
  // Bindings to f978

  // f980
  logic [0:0] f980_wen;
  logic [31:0] f980_wdata;
  logic [0:0] f980_clk;
  logic [0:0] f980_rst;
  logic [31:0] f980_rdata;
  sr_buffer_32_1 f980(.wen(f980_wen), .wdata(f980_wdata), .clk(f980_clk), .rst(f980_rst), .rdata(f980_rdata));
  assign f980_clk = clk;
  assign f980_rst = rst;
  // Bindings to f980

  // f982
  logic [0:0] f982_wen;
  logic [31:0] f982_wdata;
  logic [0:0] f982_clk;
  logic [0:0] f982_rst;
  logic [31:0] f982_rdata;
  sr_buffer_32_1 f982(.wen(f982_wen), .wdata(f982_wdata), .clk(f982_clk), .rst(f982_rst), .rdata(f982_rdata));
  assign f982_clk = clk;
  assign f982_rst = rst;
  // Bindings to f982

  // f984
  logic [0:0] f984_wen;
  logic [31:0] f984_wdata;
  logic [0:0] f984_clk;
  logic [0:0] f984_rst;
  logic [31:0] f984_rdata;
  sr_buffer_32_1 f984(.wen(f984_wen), .wdata(f984_wdata), .clk(f984_clk), .rst(f984_rst), .rdata(f984_rdata));
  assign f984_clk = clk;
  assign f984_rst = rst;
  // Bindings to f984

  // f986
  logic [0:0] f986_wen;
  logic [31:0] f986_wdata;
  logic [0:0] f986_clk;
  logic [0:0] f986_rst;
  logic [31:0] f986_rdata;
  sr_buffer_32_1 f986(.wen(f986_wen), .wdata(f986_wdata), .clk(f986_clk), .rst(f986_rst), .rdata(f986_rdata));
  assign f986_clk = clk;
  assign f986_rst = rst;
  // Bindings to f986

  // f988
  logic [0:0] f988_wen;
  logic [31:0] f988_wdata;
  logic [0:0] f988_clk;
  logic [0:0] f988_rst;
  logic [31:0] f988_rdata;
  sr_buffer_32_1 f988(.wen(f988_wen), .wdata(f988_wdata), .clk(f988_clk), .rst(f988_rst), .rdata(f988_rdata));
  assign f988_clk = clk;
  assign f988_rst = rst;
  // Bindings to f988

  // f990
  logic [0:0] f990_wen;
  logic [31:0] f990_wdata;
  logic [0:0] f990_clk;
  logic [0:0] f990_rst;
  logic [31:0] f990_rdata;
  sr_buffer_32_1 f990(.wen(f990_wen), .wdata(f990_wdata), .clk(f990_clk), .rst(f990_rst), .rdata(f990_rdata));
  assign f990_clk = clk;
  assign f990_rst = rst;
  // Bindings to f990

  // f992
  logic [0:0] f992_wen;
  logic [31:0] f992_wdata;
  logic [0:0] f992_clk;
  logic [0:0] f992_rst;
  logic [31:0] f992_rdata;
  sr_buffer_32_1 f992(.wen(f992_wen), .wdata(f992_wdata), .clk(f992_clk), .rst(f992_rst), .rdata(f992_rdata));
  assign f992_clk = clk;
  assign f992_rst = rst;
  // Bindings to f992

  // f994
  logic [0:0] f994_wen;
  logic [31:0] f994_wdata;
  logic [0:0] f994_clk;
  logic [0:0] f994_rst;
  logic [31:0] f994_rdata;
  sr_buffer_32_1 f994(.wen(f994_wen), .wdata(f994_wdata), .clk(f994_clk), .rst(f994_rst), .rdata(f994_rdata));
  assign f994_clk = clk;
  assign f994_rst = rst;
  // Bindings to f994

  // f996
  logic [0:0] f996_wen;
  logic [31:0] f996_wdata;
  logic [0:0] f996_clk;
  logic [0:0] f996_rst;
  logic [31:0] f996_rdata;
  sr_buffer_32_1 f996(.wen(f996_wen), .wdata(f996_wdata), .clk(f996_clk), .rst(f996_rst), .rdata(f996_rdata));
  assign f996_clk = clk;
  assign f996_rst = rst;
  // Bindings to f996

  // f998
  logic [0:0] f998_wen;
  logic [31:0] f998_wdata;
  logic [0:0] f998_clk;
  logic [0:0] f998_rst;
  logic [31:0] f998_rdata;
  sr_buffer_32_1 f998(.wen(f998_wen), .wdata(f998_wdata), .clk(f998_clk), .rst(f998_rst), .rdata(f998_rdata));
  assign f998_clk = clk;
  assign f998_rst = rst;
  // Bindings to f998

  // f1000
  logic [0:0] f1000_wen;
  logic [31:0] f1000_wdata;
  logic [0:0] f1000_clk;
  logic [0:0] f1000_rst;
  logic [31:0] f1000_rdata;
  sr_buffer_32_1 f1000(.wen(f1000_wen), .wdata(f1000_wdata), .clk(f1000_clk), .rst(f1000_rst), .rdata(f1000_rdata));
  assign f1000_clk = clk;
  assign f1000_rst = rst;
  // Bindings to f1000

  // f1002
  logic [0:0] f1002_wen;
  logic [31:0] f1002_wdata;
  logic [0:0] f1002_clk;
  logic [0:0] f1002_rst;
  logic [31:0] f1002_rdata;
  sr_buffer_32_1 f1002(.wen(f1002_wen), .wdata(f1002_wdata), .clk(f1002_clk), .rst(f1002_rst), .rdata(f1002_rdata));
  assign f1002_clk = clk;
  assign f1002_rst = rst;
  // Bindings to f1002

  // f1004
  logic [0:0] f1004_wen;
  logic [31:0] f1004_wdata;
  logic [0:0] f1004_clk;
  logic [0:0] f1004_rst;
  logic [31:0] f1004_rdata;
  sr_buffer_32_1 f1004(.wen(f1004_wen), .wdata(f1004_wdata), .clk(f1004_clk), .rst(f1004_rst), .rdata(f1004_rdata));
  assign f1004_clk = clk;
  assign f1004_rst = rst;
  // Bindings to f1004

  // f1006
  logic [0:0] f1006_wen;
  logic [31:0] f1006_wdata;
  logic [0:0] f1006_clk;
  logic [0:0] f1006_rst;
  logic [31:0] f1006_rdata;
  sr_buffer_32_1 f1006(.wen(f1006_wen), .wdata(f1006_wdata), .clk(f1006_clk), .rst(f1006_rst), .rdata(f1006_rdata));
  assign f1006_clk = clk;
  assign f1006_rst = rst;
  // Bindings to f1006

  // f1008
  logic [0:0] f1008_wen;
  logic [31:0] f1008_wdata;
  logic [0:0] f1008_clk;
  logic [0:0] f1008_rst;
  logic [31:0] f1008_rdata;
  sr_buffer_32_1 f1008(.wen(f1008_wen), .wdata(f1008_wdata), .clk(f1008_clk), .rst(f1008_rst), .rdata(f1008_rdata));
  assign f1008_clk = clk;
  assign f1008_rst = rst;
  // Bindings to f1008

  // f1010
  logic [0:0] f1010_wen;
  logic [31:0] f1010_wdata;
  logic [0:0] f1010_clk;
  logic [0:0] f1010_rst;
  logic [31:0] f1010_rdata;
  sr_buffer_32_1 f1010(.wen(f1010_wen), .wdata(f1010_wdata), .clk(f1010_clk), .rst(f1010_rst), .rdata(f1010_rdata));
  assign f1010_clk = clk;
  assign f1010_rst = rst;
  // Bindings to f1010

  // f1012
  logic [0:0] f1012_wen;
  logic [31:0] f1012_wdata;
  logic [0:0] f1012_clk;
  logic [0:0] f1012_rst;
  logic [31:0] f1012_rdata;
  sr_buffer_32_1 f1012(.wen(f1012_wen), .wdata(f1012_wdata), .clk(f1012_clk), .rst(f1012_rst), .rdata(f1012_rdata));
  assign f1012_clk = clk;
  assign f1012_rst = rst;
  // Bindings to f1012

  // f1014
  logic [0:0] f1014_wen;
  logic [31:0] f1014_wdata;
  logic [0:0] f1014_clk;
  logic [0:0] f1014_rst;
  logic [31:0] f1014_rdata;
  sr_buffer_32_1 f1014(.wen(f1014_wen), .wdata(f1014_wdata), .clk(f1014_clk), .rst(f1014_rst), .rdata(f1014_rdata));
  assign f1014_clk = clk;
  assign f1014_rst = rst;
  // Bindings to f1014

  // f1016
  logic [0:0] f1016_wen;
  logic [31:0] f1016_wdata;
  logic [0:0] f1016_clk;
  logic [0:0] f1016_rst;
  logic [31:0] f1016_rdata;
  sr_buffer_32_1 f1016(.wen(f1016_wen), .wdata(f1016_wdata), .clk(f1016_clk), .rst(f1016_rst), .rdata(f1016_rdata));
  assign f1016_clk = clk;
  assign f1016_rst = rst;
  // Bindings to f1016

  // f1018
  logic [0:0] f1018_wen;
  logic [31:0] f1018_wdata;
  logic [0:0] f1018_clk;
  logic [0:0] f1018_rst;
  logic [31:0] f1018_rdata;
  sr_buffer_32_1 f1018(.wen(f1018_wen), .wdata(f1018_wdata), .clk(f1018_clk), .rst(f1018_rst), .rdata(f1018_rdata));
  assign f1018_clk = clk;
  assign f1018_rst = rst;
  // Bindings to f1018

  // f1020
  logic [0:0] f1020_wen;
  logic [31:0] f1020_wdata;
  logic [0:0] f1020_clk;
  logic [0:0] f1020_rst;
  logic [31:0] f1020_rdata;
  sr_buffer_32_1 f1020(.wen(f1020_wen), .wdata(f1020_wdata), .clk(f1020_clk), .rst(f1020_rst), .rdata(f1020_rdata));
  assign f1020_clk = clk;
  assign f1020_rst = rst;
  // Bindings to f1020

  // f1022
  logic [0:0] f1022_wen;
  logic [31:0] f1022_wdata;
  logic [0:0] f1022_clk;
  logic [0:0] f1022_rst;
  logic [31:0] f1022_rdata;
  sr_buffer_32_1 f1022(.wen(f1022_wen), .wdata(f1022_wdata), .clk(f1022_clk), .rst(f1022_rst), .rdata(f1022_rdata));
  assign f1022_clk = clk;
  assign f1022_rst = rst;
  // Bindings to f1022

  // f1024
  logic [0:0] f1024_wen;
  logic [31:0] f1024_wdata;
  logic [0:0] f1024_clk;
  logic [0:0] f1024_rst;
  logic [31:0] f1024_rdata;
  sr_buffer_32_1 f1024(.wen(f1024_wen), .wdata(f1024_wdata), .clk(f1024_clk), .rst(f1024_rst), .rdata(f1024_rdata));
  assign f1024_clk = clk;
  assign f1024_rst = rst;
  // Bindings to f1024

  // f1026
  logic [0:0] f1026_wen;
  logic [31:0] f1026_wdata;
  logic [0:0] f1026_clk;
  logic [0:0] f1026_rst;
  logic [31:0] f1026_rdata;
  sr_buffer_32_1 f1026(.wen(f1026_wen), .wdata(f1026_wdata), .clk(f1026_clk), .rst(f1026_rst), .rdata(f1026_rdata));
  assign f1026_clk = clk;
  assign f1026_rst = rst;
  // Bindings to f1026

  // f1028
  logic [0:0] f1028_wen;
  logic [31:0] f1028_wdata;
  logic [0:0] f1028_clk;
  logic [0:0] f1028_rst;
  logic [31:0] f1028_rdata;
  sr_buffer_32_1 f1028(.wen(f1028_wen), .wdata(f1028_wdata), .clk(f1028_clk), .rst(f1028_rst), .rdata(f1028_rdata));
  assign f1028_clk = clk;
  assign f1028_rst = rst;
  // Bindings to f1028

  // f1030
  logic [0:0] f1030_wen;
  logic [31:0] f1030_wdata;
  logic [0:0] f1030_clk;
  logic [0:0] f1030_rst;
  logic [31:0] f1030_rdata;
  sr_buffer_32_1 f1030(.wen(f1030_wen), .wdata(f1030_wdata), .clk(f1030_clk), .rst(f1030_rst), .rdata(f1030_rdata));
  assign f1030_clk = clk;
  assign f1030_rst = rst;
  // Bindings to f1030

  // f1032
  logic [0:0] f1032_wen;
  logic [31:0] f1032_wdata;
  logic [0:0] f1032_clk;
  logic [0:0] f1032_rst;
  logic [31:0] f1032_rdata;
  sr_buffer_32_1 f1032(.wen(f1032_wen), .wdata(f1032_wdata), .clk(f1032_clk), .rst(f1032_rst), .rdata(f1032_rdata));
  assign f1032_clk = clk;
  assign f1032_rst = rst;
  // Bindings to f1032

  // f1034
  logic [0:0] f1034_wen;
  logic [31:0] f1034_wdata;
  logic [0:0] f1034_clk;
  logic [0:0] f1034_rst;
  logic [31:0] f1034_rdata;
  sr_buffer_32_1 f1034(.wen(f1034_wen), .wdata(f1034_wdata), .clk(f1034_clk), .rst(f1034_rst), .rdata(f1034_rdata));
  assign f1034_clk = clk;
  assign f1034_rst = rst;
  // Bindings to f1034

  // f1036
  logic [0:0] f1036_wen;
  logic [31:0] f1036_wdata;
  logic [0:0] f1036_clk;
  logic [0:0] f1036_rst;
  logic [31:0] f1036_rdata;
  sr_buffer_32_1 f1036(.wen(f1036_wen), .wdata(f1036_wdata), .clk(f1036_clk), .rst(f1036_rst), .rdata(f1036_rdata));
  assign f1036_clk = clk;
  assign f1036_rst = rst;
  // Bindings to f1036

  // f1038
  logic [0:0] f1038_wen;
  logic [31:0] f1038_wdata;
  logic [0:0] f1038_clk;
  logic [0:0] f1038_rst;
  logic [31:0] f1038_rdata;
  sr_buffer_32_1 f1038(.wen(f1038_wen), .wdata(f1038_wdata), .clk(f1038_clk), .rst(f1038_rst), .rdata(f1038_rdata));
  assign f1038_clk = clk;
  assign f1038_rst = rst;
  // Bindings to f1038

  // f1040
  logic [0:0] f1040_wen;
  logic [31:0] f1040_wdata;
  logic [0:0] f1040_clk;
  logic [0:0] f1040_rst;
  logic [31:0] f1040_rdata;
  sr_buffer_32_1 f1040(.wen(f1040_wen), .wdata(f1040_wdata), .clk(f1040_clk), .rst(f1040_rst), .rdata(f1040_rdata));
  assign f1040_clk = clk;
  assign f1040_rst = rst;
  // Bindings to f1040

  // f1042
  logic [0:0] f1042_wen;
  logic [31:0] f1042_wdata;
  logic [0:0] f1042_clk;
  logic [0:0] f1042_rst;
  logic [31:0] f1042_rdata;
  sr_buffer_32_1 f1042(.wen(f1042_wen), .wdata(f1042_wdata), .clk(f1042_clk), .rst(f1042_rst), .rdata(f1042_rdata));
  assign f1042_clk = clk;
  assign f1042_rst = rst;
  // Bindings to f1042

  // f1044
  logic [0:0] f1044_wen;
  logic [31:0] f1044_wdata;
  logic [0:0] f1044_clk;
  logic [0:0] f1044_rst;
  logic [31:0] f1044_rdata;
  sr_buffer_32_1 f1044(.wen(f1044_wen), .wdata(f1044_wdata), .clk(f1044_clk), .rst(f1044_rst), .rdata(f1044_rdata));
  assign f1044_clk = clk;
  assign f1044_rst = rst;
  // Bindings to f1044

  // f1046
  logic [0:0] f1046_wen;
  logic [31:0] f1046_wdata;
  logic [0:0] f1046_clk;
  logic [0:0] f1046_rst;
  logic [31:0] f1046_rdata;
  sr_buffer_32_1 f1046(.wen(f1046_wen), .wdata(f1046_wdata), .clk(f1046_clk), .rst(f1046_rst), .rdata(f1046_rdata));
  assign f1046_clk = clk;
  assign f1046_rst = rst;
  // Bindings to f1046

  // f1048
  logic [0:0] f1048_wen;
  logic [31:0] f1048_wdata;
  logic [0:0] f1048_clk;
  logic [0:0] f1048_rst;
  logic [31:0] f1048_rdata;
  sr_buffer_32_1 f1048(.wen(f1048_wen), .wdata(f1048_wdata), .clk(f1048_clk), .rst(f1048_rst), .rdata(f1048_rdata));
  assign f1048_clk = clk;
  assign f1048_rst = rst;
  // Bindings to f1048

  // f1050
  logic [0:0] f1050_wen;
  logic [31:0] f1050_wdata;
  logic [0:0] f1050_clk;
  logic [0:0] f1050_rst;
  logic [31:0] f1050_rdata;
  sr_buffer_32_1 f1050(.wen(f1050_wen), .wdata(f1050_wdata), .clk(f1050_clk), .rst(f1050_rst), .rdata(f1050_rdata));
  assign f1050_clk = clk;
  assign f1050_rst = rst;
  // Bindings to f1050

  // f1052
  logic [0:0] f1052_wen;
  logic [31:0] f1052_wdata;
  logic [0:0] f1052_clk;
  logic [0:0] f1052_rst;
  logic [31:0] f1052_rdata;
  sr_buffer_32_1 f1052(.wen(f1052_wen), .wdata(f1052_wdata), .clk(f1052_clk), .rst(f1052_rst), .rdata(f1052_rdata));
  assign f1052_clk = clk;
  assign f1052_rst = rst;
  // Bindings to f1052

  // f1054
  logic [0:0] f1054_wen;
  logic [31:0] f1054_wdata;
  logic [0:0] f1054_clk;
  logic [0:0] f1054_rst;
  logic [31:0] f1054_rdata;
  sr_buffer_32_1 f1054(.wen(f1054_wen), .wdata(f1054_wdata), .clk(f1054_clk), .rst(f1054_rst), .rdata(f1054_rdata));
  assign f1054_clk = clk;
  assign f1054_rst = rst;
  // Bindings to f1054

  // f1056
  logic [0:0] f1056_wen;
  logic [31:0] f1056_wdata;
  logic [0:0] f1056_clk;
  logic [0:0] f1056_rst;
  logic [31:0] f1056_rdata;
  sr_buffer_32_1 f1056(.wen(f1056_wen), .wdata(f1056_wdata), .clk(f1056_clk), .rst(f1056_rst), .rdata(f1056_rdata));
  assign f1056_clk = clk;
  assign f1056_rst = rst;
  // Bindings to f1056

  // f1058
  logic [0:0] f1058_wen;
  logic [31:0] f1058_wdata;
  logic [0:0] f1058_clk;
  logic [0:0] f1058_rst;
  logic [31:0] f1058_rdata;
  sr_buffer_32_1 f1058(.wen(f1058_wen), .wdata(f1058_wdata), .clk(f1058_clk), .rst(f1058_rst), .rdata(f1058_rdata));
  assign f1058_clk = clk;
  assign f1058_rst = rst;
  // Bindings to f1058

  // f1060
  logic [0:0] f1060_wen;
  logic [31:0] f1060_wdata;
  logic [0:0] f1060_clk;
  logic [0:0] f1060_rst;
  logic [31:0] f1060_rdata;
  sr_buffer_32_1 f1060(.wen(f1060_wen), .wdata(f1060_wdata), .clk(f1060_clk), .rst(f1060_rst), .rdata(f1060_rdata));
  assign f1060_clk = clk;
  assign f1060_rst = rst;
  // Bindings to f1060

  // f1062
  logic [0:0] f1062_wen;
  logic [31:0] f1062_wdata;
  logic [0:0] f1062_clk;
  logic [0:0] f1062_rst;
  logic [31:0] f1062_rdata;
  sr_buffer_32_1 f1062(.wen(f1062_wen), .wdata(f1062_wdata), .clk(f1062_clk), .rst(f1062_rst), .rdata(f1062_rdata));
  assign f1062_clk = clk;
  assign f1062_rst = rst;
  // Bindings to f1062

  // f1064
  logic [0:0] f1064_wen;
  logic [31:0] f1064_wdata;
  logic [0:0] f1064_clk;
  logic [0:0] f1064_rst;
  logic [31:0] f1064_rdata;
  sr_buffer_32_1 f1064(.wen(f1064_wen), .wdata(f1064_wdata), .clk(f1064_clk), .rst(f1064_rst), .rdata(f1064_rdata));
  assign f1064_clk = clk;
  assign f1064_rst = rst;
  // Bindings to f1064

  // f1066
  logic [0:0] f1066_wen;
  logic [31:0] f1066_wdata;
  logic [0:0] f1066_clk;
  logic [0:0] f1066_rst;
  logic [31:0] f1066_rdata;
  sr_buffer_32_1 f1066(.wen(f1066_wen), .wdata(f1066_wdata), .clk(f1066_clk), .rst(f1066_rst), .rdata(f1066_rdata));
  assign f1066_clk = clk;
  assign f1066_rst = rst;
  // Bindings to f1066

  // f1068
  logic [0:0] f1068_wen;
  logic [31:0] f1068_wdata;
  logic [0:0] f1068_clk;
  logic [0:0] f1068_rst;
  logic [31:0] f1068_rdata;
  sr_buffer_32_1 f1068(.wen(f1068_wen), .wdata(f1068_wdata), .clk(f1068_clk), .rst(f1068_rst), .rdata(f1068_rdata));
  assign f1068_clk = clk;
  assign f1068_rst = rst;
  // Bindings to f1068

  // f1070
  logic [0:0] f1070_wen;
  logic [31:0] f1070_wdata;
  logic [0:0] f1070_clk;
  logic [0:0] f1070_rst;
  logic [31:0] f1070_rdata;
  sr_buffer_32_1 f1070(.wen(f1070_wen), .wdata(f1070_wdata), .clk(f1070_clk), .rst(f1070_rst), .rdata(f1070_rdata));
  assign f1070_clk = clk;
  assign f1070_rst = rst;
  // Bindings to f1070

  // f1072
  logic [0:0] f1072_wen;
  logic [31:0] f1072_wdata;
  logic [0:0] f1072_clk;
  logic [0:0] f1072_rst;
  logic [31:0] f1072_rdata;
  sr_buffer_32_1 f1072(.wen(f1072_wen), .wdata(f1072_wdata), .clk(f1072_clk), .rst(f1072_rst), .rdata(f1072_rdata));
  assign f1072_clk = clk;
  assign f1072_rst = rst;
  // Bindings to f1072

  // f1074
  logic [0:0] f1074_wen;
  logic [31:0] f1074_wdata;
  logic [0:0] f1074_clk;
  logic [0:0] f1074_rst;
  logic [31:0] f1074_rdata;
  sr_buffer_32_1 f1074(.wen(f1074_wen), .wdata(f1074_wdata), .clk(f1074_clk), .rst(f1074_rst), .rdata(f1074_rdata));
  assign f1074_clk = clk;
  assign f1074_rst = rst;
  // Bindings to f1074

  // f1076
  logic [0:0] f1076_wen;
  logic [31:0] f1076_wdata;
  logic [0:0] f1076_clk;
  logic [0:0] f1076_rst;
  logic [31:0] f1076_rdata;
  sr_buffer_32_1 f1076(.wen(f1076_wen), .wdata(f1076_wdata), .clk(f1076_clk), .rst(f1076_rst), .rdata(f1076_rdata));
  assign f1076_clk = clk;
  assign f1076_rst = rst;
  // Bindings to f1076

  // f1078
  logic [0:0] f1078_wen;
  logic [31:0] f1078_wdata;
  logic [0:0] f1078_clk;
  logic [0:0] f1078_rst;
  logic [31:0] f1078_rdata;
  sr_buffer_32_1 f1078(.wen(f1078_wen), .wdata(f1078_wdata), .clk(f1078_clk), .rst(f1078_rst), .rdata(f1078_rdata));
  assign f1078_clk = clk;
  assign f1078_rst = rst;
  // Bindings to f1078

  // f1080
  logic [0:0] f1080_wen;
  logic [31:0] f1080_wdata;
  logic [0:0] f1080_clk;
  logic [0:0] f1080_rst;
  logic [31:0] f1080_rdata;
  sr_buffer_32_1 f1080(.wen(f1080_wen), .wdata(f1080_wdata), .clk(f1080_clk), .rst(f1080_rst), .rdata(f1080_rdata));
  assign f1080_clk = clk;
  assign f1080_rst = rst;
  // Bindings to f1080

  // f1082
  logic [0:0] f1082_wen;
  logic [31:0] f1082_wdata;
  logic [0:0] f1082_clk;
  logic [0:0] f1082_rst;
  logic [31:0] f1082_rdata;
  sr_buffer_32_1 f1082(.wen(f1082_wen), .wdata(f1082_wdata), .clk(f1082_clk), .rst(f1082_rst), .rdata(f1082_rdata));
  assign f1082_clk = clk;
  assign f1082_rst = rst;
  // Bindings to f1082

  // f1084
  logic [0:0] f1084_wen;
  logic [31:0] f1084_wdata;
  logic [0:0] f1084_clk;
  logic [0:0] f1084_rst;
  logic [31:0] f1084_rdata;
  sr_buffer_32_1 f1084(.wen(f1084_wen), .wdata(f1084_wdata), .clk(f1084_clk), .rst(f1084_rst), .rdata(f1084_rdata));
  assign f1084_clk = clk;
  assign f1084_rst = rst;
  // Bindings to f1084

  // f1086
  logic [0:0] f1086_wen;
  logic [31:0] f1086_wdata;
  logic [0:0] f1086_clk;
  logic [0:0] f1086_rst;
  logic [31:0] f1086_rdata;
  sr_buffer_32_1 f1086(.wen(f1086_wen), .wdata(f1086_wdata), .clk(f1086_clk), .rst(f1086_rst), .rdata(f1086_rdata));
  assign f1086_clk = clk;
  assign f1086_rst = rst;
  // Bindings to f1086

  // f1088
  logic [0:0] f1088_wen;
  logic [31:0] f1088_wdata;
  logic [0:0] f1088_clk;
  logic [0:0] f1088_rst;
  logic [31:0] f1088_rdata;
  sr_buffer_32_1 f1088(.wen(f1088_wen), .wdata(f1088_wdata), .clk(f1088_clk), .rst(f1088_rst), .rdata(f1088_rdata));
  assign f1088_clk = clk;
  assign f1088_rst = rst;
  // Bindings to f1088

  // f1090
  logic [0:0] f1090_wen;
  logic [31:0] f1090_wdata;
  logic [0:0] f1090_clk;
  logic [0:0] f1090_rst;
  logic [31:0] f1090_rdata;
  sr_buffer_32_1 f1090(.wen(f1090_wen), .wdata(f1090_wdata), .clk(f1090_clk), .rst(f1090_rst), .rdata(f1090_rdata));
  assign f1090_clk = clk;
  assign f1090_rst = rst;
  // Bindings to f1090

  // f1092
  logic [0:0] f1092_wen;
  logic [31:0] f1092_wdata;
  logic [0:0] f1092_clk;
  logic [0:0] f1092_rst;
  logic [31:0] f1092_rdata;
  sr_buffer_32_1 f1092(.wen(f1092_wen), .wdata(f1092_wdata), .clk(f1092_clk), .rst(f1092_rst), .rdata(f1092_rdata));
  assign f1092_clk = clk;
  assign f1092_rst = rst;
  // Bindings to f1092

  // f1094
  logic [0:0] f1094_wen;
  logic [31:0] f1094_wdata;
  logic [0:0] f1094_clk;
  logic [0:0] f1094_rst;
  logic [31:0] f1094_rdata;
  sr_buffer_32_1 f1094(.wen(f1094_wen), .wdata(f1094_wdata), .clk(f1094_clk), .rst(f1094_rst), .rdata(f1094_rdata));
  assign f1094_clk = clk;
  assign f1094_rst = rst;
  // Bindings to f1094

  // f1096
  logic [0:0] f1096_wen;
  logic [31:0] f1096_wdata;
  logic [0:0] f1096_clk;
  logic [0:0] f1096_rst;
  logic [31:0] f1096_rdata;
  sr_buffer_32_1 f1096(.wen(f1096_wen), .wdata(f1096_wdata), .clk(f1096_clk), .rst(f1096_rst), .rdata(f1096_rdata));
  assign f1096_clk = clk;
  assign f1096_rst = rst;
  // Bindings to f1096

  // f1098
  logic [0:0] f1098_wen;
  logic [31:0] f1098_wdata;
  logic [0:0] f1098_clk;
  logic [0:0] f1098_rst;
  logic [31:0] f1098_rdata;
  sr_buffer_32_1 f1098(.wen(f1098_wen), .wdata(f1098_wdata), .clk(f1098_clk), .rst(f1098_rst), .rdata(f1098_rdata));
  assign f1098_clk = clk;
  assign f1098_rst = rst;
  // Bindings to f1098

  // f1100
  logic [0:0] f1100_wen;
  logic [31:0] f1100_wdata;
  logic [0:0] f1100_clk;
  logic [0:0] f1100_rst;
  logic [31:0] f1100_rdata;
  sr_buffer_32_1 f1100(.wen(f1100_wen), .wdata(f1100_wdata), .clk(f1100_clk), .rst(f1100_rst), .rdata(f1100_rdata));
  assign f1100_clk = clk;
  assign f1100_rst = rst;
  // Bindings to f1100

  // f1102
  logic [0:0] f1102_wen;
  logic [31:0] f1102_wdata;
  logic [0:0] f1102_clk;
  logic [0:0] f1102_rst;
  logic [31:0] f1102_rdata;
  sr_buffer_32_1 f1102(.wen(f1102_wen), .wdata(f1102_wdata), .clk(f1102_clk), .rst(f1102_rst), .rdata(f1102_rdata));
  assign f1102_clk = clk;
  assign f1102_rst = rst;
  // Bindings to f1102

  // f1104
  logic [0:0] f1104_wen;
  logic [31:0] f1104_wdata;
  logic [0:0] f1104_clk;
  logic [0:0] f1104_rst;
  logic [31:0] f1104_rdata;
  sr_buffer_32_1 f1104(.wen(f1104_wen), .wdata(f1104_wdata), .clk(f1104_clk), .rst(f1104_rst), .rdata(f1104_rdata));
  assign f1104_clk = clk;
  assign f1104_rst = rst;
  // Bindings to f1104

  // f1106
  logic [0:0] f1106_wen;
  logic [31:0] f1106_wdata;
  logic [0:0] f1106_clk;
  logic [0:0] f1106_rst;
  logic [31:0] f1106_rdata;
  sr_buffer_32_1 f1106(.wen(f1106_wen), .wdata(f1106_wdata), .clk(f1106_clk), .rst(f1106_rst), .rdata(f1106_rdata));
  assign f1106_clk = clk;
  assign f1106_rst = rst;
  // Bindings to f1106

  // f1108
  logic [0:0] f1108_wen;
  logic [31:0] f1108_wdata;
  logic [0:0] f1108_clk;
  logic [0:0] f1108_rst;
  logic [31:0] f1108_rdata;
  sr_buffer_32_1 f1108(.wen(f1108_wen), .wdata(f1108_wdata), .clk(f1108_clk), .rst(f1108_rst), .rdata(f1108_rdata));
  assign f1108_clk = clk;
  assign f1108_rst = rst;
  // Bindings to f1108

  // f1110
  logic [0:0] f1110_wen;
  logic [31:0] f1110_wdata;
  logic [0:0] f1110_clk;
  logic [0:0] f1110_rst;
  logic [31:0] f1110_rdata;
  sr_buffer_32_1 f1110(.wen(f1110_wen), .wdata(f1110_wdata), .clk(f1110_clk), .rst(f1110_rst), .rdata(f1110_rdata));
  assign f1110_clk = clk;
  assign f1110_rst = rst;
  // Bindings to f1110

  // f1112
  logic [0:0] f1112_wen;
  logic [31:0] f1112_wdata;
  logic [0:0] f1112_clk;
  logic [0:0] f1112_rst;
  logic [31:0] f1112_rdata;
  sr_buffer_32_1 f1112(.wen(f1112_wen), .wdata(f1112_wdata), .clk(f1112_clk), .rst(f1112_rst), .rdata(f1112_rdata));
  assign f1112_clk = clk;
  assign f1112_rst = rst;
  // Bindings to f1112

  // f1114
  logic [0:0] f1114_wen;
  logic [31:0] f1114_wdata;
  logic [0:0] f1114_clk;
  logic [0:0] f1114_rst;
  logic [31:0] f1114_rdata;
  sr_buffer_32_1 f1114(.wen(f1114_wen), .wdata(f1114_wdata), .clk(f1114_clk), .rst(f1114_rst), .rdata(f1114_rdata));
  assign f1114_clk = clk;
  assign f1114_rst = rst;
  // Bindings to f1114

  // f1116
  logic [0:0] f1116_wen;
  logic [31:0] f1116_wdata;
  logic [0:0] f1116_clk;
  logic [0:0] f1116_rst;
  logic [31:0] f1116_rdata;
  sr_buffer_32_1 f1116(.wen(f1116_wen), .wdata(f1116_wdata), .clk(f1116_clk), .rst(f1116_rst), .rdata(f1116_rdata));
  assign f1116_clk = clk;
  assign f1116_rst = rst;
  // Bindings to f1116

  // f1118
  logic [0:0] f1118_wen;
  logic [31:0] f1118_wdata;
  logic [0:0] f1118_clk;
  logic [0:0] f1118_rst;
  logic [31:0] f1118_rdata;
  sr_buffer_32_1 f1118(.wen(f1118_wen), .wdata(f1118_wdata), .clk(f1118_clk), .rst(f1118_rst), .rdata(f1118_rdata));
  assign f1118_clk = clk;
  assign f1118_rst = rst;
  // Bindings to f1118

  // f1120
  logic [0:0] f1120_wen;
  logic [31:0] f1120_wdata;
  logic [0:0] f1120_clk;
  logic [0:0] f1120_rst;
  logic [31:0] f1120_rdata;
  sr_buffer_32_1 f1120(.wen(f1120_wen), .wdata(f1120_wdata), .clk(f1120_clk), .rst(f1120_rst), .rdata(f1120_rdata));
  assign f1120_clk = clk;
  assign f1120_rst = rst;
  // Bindings to f1120

  // f1122
  logic [0:0] f1122_wen;
  logic [31:0] f1122_wdata;
  logic [0:0] f1122_clk;
  logic [0:0] f1122_rst;
  logic [31:0] f1122_rdata;
  sr_buffer_32_1 f1122(.wen(f1122_wen), .wdata(f1122_wdata), .clk(f1122_clk), .rst(f1122_rst), .rdata(f1122_rdata));
  assign f1122_clk = clk;
  assign f1122_rst = rst;
  // Bindings to f1122

  // f1124
  logic [0:0] f1124_wen;
  logic [31:0] f1124_wdata;
  logic [0:0] f1124_clk;
  logic [0:0] f1124_rst;
  logic [31:0] f1124_rdata;
  sr_buffer_32_1 f1124(.wen(f1124_wen), .wdata(f1124_wdata), .clk(f1124_clk), .rst(f1124_rst), .rdata(f1124_rdata));
  assign f1124_clk = clk;
  assign f1124_rst = rst;
  // Bindings to f1124

  // f1126
  logic [0:0] f1126_wen;
  logic [31:0] f1126_wdata;
  logic [0:0] f1126_clk;
  logic [0:0] f1126_rst;
  logic [31:0] f1126_rdata;
  sr_buffer_32_1 f1126(.wen(f1126_wen), .wdata(f1126_wdata), .clk(f1126_clk), .rst(f1126_rst), .rdata(f1126_rdata));
  assign f1126_clk = clk;
  assign f1126_rst = rst;
  // Bindings to f1126

  // f1128
  logic [0:0] f1128_wen;
  logic [31:0] f1128_wdata;
  logic [0:0] f1128_clk;
  logic [0:0] f1128_rst;
  logic [31:0] f1128_rdata;
  sr_buffer_32_1 f1128(.wen(f1128_wen), .wdata(f1128_wdata), .clk(f1128_clk), .rst(f1128_rst), .rdata(f1128_rdata));
  assign f1128_clk = clk;
  assign f1128_rst = rst;
  // Bindings to f1128

  // f1130
  logic [0:0] f1130_wen;
  logic [31:0] f1130_wdata;
  logic [0:0] f1130_clk;
  logic [0:0] f1130_rst;
  logic [31:0] f1130_rdata;
  sr_buffer_32_1 f1130(.wen(f1130_wen), .wdata(f1130_wdata), .clk(f1130_clk), .rst(f1130_rst), .rdata(f1130_rdata));
  assign f1130_clk = clk;
  assign f1130_rst = rst;
  // Bindings to f1130

  // f1132
  logic [0:0] f1132_wen;
  logic [31:0] f1132_wdata;
  logic [0:0] f1132_clk;
  logic [0:0] f1132_rst;
  logic [31:0] f1132_rdata;
  sr_buffer_32_1 f1132(.wen(f1132_wen), .wdata(f1132_wdata), .clk(f1132_clk), .rst(f1132_rst), .rdata(f1132_rdata));
  assign f1132_clk = clk;
  assign f1132_rst = rst;
  // Bindings to f1132

  // f1134
  logic [0:0] f1134_wen;
  logic [31:0] f1134_wdata;
  logic [0:0] f1134_clk;
  logic [0:0] f1134_rst;
  logic [31:0] f1134_rdata;
  sr_buffer_32_1 f1134(.wen(f1134_wen), .wdata(f1134_wdata), .clk(f1134_clk), .rst(f1134_rst), .rdata(f1134_rdata));
  assign f1134_clk = clk;
  assign f1134_rst = rst;
  // Bindings to f1134

  // f1136
  logic [0:0] f1136_wen;
  logic [31:0] f1136_wdata;
  logic [0:0] f1136_clk;
  logic [0:0] f1136_rst;
  logic [31:0] f1136_rdata;
  sr_buffer_32_1 f1136(.wen(f1136_wen), .wdata(f1136_wdata), .clk(f1136_clk), .rst(f1136_rst), .rdata(f1136_rdata));
  assign f1136_clk = clk;
  assign f1136_rst = rst;
  // Bindings to f1136

  // f1138
  logic [0:0] f1138_wen;
  logic [31:0] f1138_wdata;
  logic [0:0] f1138_clk;
  logic [0:0] f1138_rst;
  logic [31:0] f1138_rdata;
  sr_buffer_32_1 f1138(.wen(f1138_wen), .wdata(f1138_wdata), .clk(f1138_clk), .rst(f1138_rst), .rdata(f1138_rdata));
  assign f1138_clk = clk;
  assign f1138_rst = rst;
  // Bindings to f1138

  // f1140
  logic [0:0] f1140_wen;
  logic [31:0] f1140_wdata;
  logic [0:0] f1140_clk;
  logic [0:0] f1140_rst;
  logic [31:0] f1140_rdata;
  sr_buffer_32_1 f1140(.wen(f1140_wen), .wdata(f1140_wdata), .clk(f1140_clk), .rst(f1140_rst), .rdata(f1140_rdata));
  assign f1140_clk = clk;
  assign f1140_rst = rst;
  // Bindings to f1140

  // f1142
  logic [0:0] f1142_wen;
  logic [31:0] f1142_wdata;
  logic [0:0] f1142_clk;
  logic [0:0] f1142_rst;
  logic [31:0] f1142_rdata;
  sr_buffer_32_1 f1142(.wen(f1142_wen), .wdata(f1142_wdata), .clk(f1142_clk), .rst(f1142_rst), .rdata(f1142_rdata));
  assign f1142_clk = clk;
  assign f1142_rst = rst;
  // Bindings to f1142

  // f1144
  logic [0:0] f1144_wen;
  logic [31:0] f1144_wdata;
  logic [0:0] f1144_clk;
  logic [0:0] f1144_rst;
  logic [31:0] f1144_rdata;
  sr_buffer_32_1 f1144(.wen(f1144_wen), .wdata(f1144_wdata), .clk(f1144_clk), .rst(f1144_rst), .rdata(f1144_rdata));
  assign f1144_clk = clk;
  assign f1144_rst = rst;
  // Bindings to f1144

  // f1146
  logic [0:0] f1146_wen;
  logic [31:0] f1146_wdata;
  logic [0:0] f1146_clk;
  logic [0:0] f1146_rst;
  logic [31:0] f1146_rdata;
  sr_buffer_32_1 f1146(.wen(f1146_wen), .wdata(f1146_wdata), .clk(f1146_clk), .rst(f1146_rst), .rdata(f1146_rdata));
  assign f1146_clk = clk;
  assign f1146_rst = rst;
  // Bindings to f1146

  // f1148
  logic [0:0] f1148_wen;
  logic [31:0] f1148_wdata;
  logic [0:0] f1148_clk;
  logic [0:0] f1148_rst;
  logic [31:0] f1148_rdata;
  sr_buffer_32_1 f1148(.wen(f1148_wen), .wdata(f1148_wdata), .clk(f1148_clk), .rst(f1148_rst), .rdata(f1148_rdata));
  assign f1148_clk = clk;
  assign f1148_rst = rst;
  // Bindings to f1148

  // f1150
  logic [0:0] f1150_wen;
  logic [31:0] f1150_wdata;
  logic [0:0] f1150_clk;
  logic [0:0] f1150_rst;
  logic [31:0] f1150_rdata;
  sr_buffer_32_1 f1150(.wen(f1150_wen), .wdata(f1150_wdata), .clk(f1150_clk), .rst(f1150_rst), .rdata(f1150_rdata));
  assign f1150_clk = clk;
  assign f1150_rst = rst;
  // Bindings to f1150

  // f1152
  logic [0:0] f1152_wen;
  logic [31:0] f1152_wdata;
  logic [0:0] f1152_clk;
  logic [0:0] f1152_rst;
  logic [31:0] f1152_rdata;
  sr_buffer_32_1 f1152(.wen(f1152_wen), .wdata(f1152_wdata), .clk(f1152_clk), .rst(f1152_rst), .rdata(f1152_rdata));
  assign f1152_clk = clk;
  assign f1152_rst = rst;
  // Bindings to f1152

  // f1154
  logic [0:0] f1154_wen;
  logic [31:0] f1154_wdata;
  logic [0:0] f1154_clk;
  logic [0:0] f1154_rst;
  logic [31:0] f1154_rdata;
  sr_buffer_32_1 f1154(.wen(f1154_wen), .wdata(f1154_wdata), .clk(f1154_clk), .rst(f1154_rst), .rdata(f1154_rdata));
  assign f1154_clk = clk;
  assign f1154_rst = rst;
  // Bindings to f1154

  // f1156
  logic [0:0] f1156_wen;
  logic [31:0] f1156_wdata;
  logic [0:0] f1156_clk;
  logic [0:0] f1156_rst;
  logic [31:0] f1156_rdata;
  sr_buffer_32_1 f1156(.wen(f1156_wen), .wdata(f1156_wdata), .clk(f1156_clk), .rst(f1156_rst), .rdata(f1156_rdata));
  assign f1156_clk = clk;
  assign f1156_rst = rst;
  // Bindings to f1156

  // f1158
  logic [0:0] f1158_wen;
  logic [31:0] f1158_wdata;
  logic [0:0] f1158_clk;
  logic [0:0] f1158_rst;
  logic [31:0] f1158_rdata;
  sr_buffer_32_1 f1158(.wen(f1158_wen), .wdata(f1158_wdata), .clk(f1158_clk), .rst(f1158_rst), .rdata(f1158_rdata));
  assign f1158_clk = clk;
  assign f1158_rst = rst;
  // Bindings to f1158

  // f1160
  logic [0:0] f1160_wen;
  logic [31:0] f1160_wdata;
  logic [0:0] f1160_clk;
  logic [0:0] f1160_rst;
  logic [31:0] f1160_rdata;
  sr_buffer_32_1 f1160(.wen(f1160_wen), .wdata(f1160_wdata), .clk(f1160_clk), .rst(f1160_rst), .rdata(f1160_rdata));
  assign f1160_clk = clk;
  assign f1160_rst = rst;
  // Bindings to f1160

  // f1162
  logic [0:0] f1162_wen;
  logic [31:0] f1162_wdata;
  logic [0:0] f1162_clk;
  logic [0:0] f1162_rst;
  logic [31:0] f1162_rdata;
  sr_buffer_32_1 f1162(.wen(f1162_wen), .wdata(f1162_wdata), .clk(f1162_clk), .rst(f1162_rst), .rdata(f1162_rdata));
  assign f1162_clk = clk;
  assign f1162_rst = rst;
  // Bindings to f1162

  // f1164
  logic [0:0] f1164_wen;
  logic [31:0] f1164_wdata;
  logic [0:0] f1164_clk;
  logic [0:0] f1164_rst;
  logic [31:0] f1164_rdata;
  sr_buffer_32_1 f1164(.wen(f1164_wen), .wdata(f1164_wdata), .clk(f1164_clk), .rst(f1164_rst), .rdata(f1164_rdata));
  assign f1164_clk = clk;
  assign f1164_rst = rst;
  // Bindings to f1164

  // f1166
  logic [0:0] f1166_wen;
  logic [31:0] f1166_wdata;
  logic [0:0] f1166_clk;
  logic [0:0] f1166_rst;
  logic [31:0] f1166_rdata;
  sr_buffer_32_1 f1166(.wen(f1166_wen), .wdata(f1166_wdata), .clk(f1166_clk), .rst(f1166_rst), .rdata(f1166_rdata));
  assign f1166_clk = clk;
  assign f1166_rst = rst;
  // Bindings to f1166

  // f1168
  logic [0:0] f1168_wen;
  logic [31:0] f1168_wdata;
  logic [0:0] f1168_clk;
  logic [0:0] f1168_rst;
  logic [31:0] f1168_rdata;
  sr_buffer_32_1 f1168(.wen(f1168_wen), .wdata(f1168_wdata), .clk(f1168_clk), .rst(f1168_rst), .rdata(f1168_rdata));
  assign f1168_clk = clk;
  assign f1168_rst = rst;
  // Bindings to f1168

  // f1170
  logic [0:0] f1170_wen;
  logic [31:0] f1170_wdata;
  logic [0:0] f1170_clk;
  logic [0:0] f1170_rst;
  logic [31:0] f1170_rdata;
  sr_buffer_32_1 f1170(.wen(f1170_wen), .wdata(f1170_wdata), .clk(f1170_clk), .rst(f1170_rst), .rdata(f1170_rdata));
  assign f1170_clk = clk;
  assign f1170_rst = rst;
  // Bindings to f1170

  // f1172
  logic [0:0] f1172_wen;
  logic [31:0] f1172_wdata;
  logic [0:0] f1172_clk;
  logic [0:0] f1172_rst;
  logic [31:0] f1172_rdata;
  sr_buffer_32_1 f1172(.wen(f1172_wen), .wdata(f1172_wdata), .clk(f1172_clk), .rst(f1172_rst), .rdata(f1172_rdata));
  assign f1172_clk = clk;
  assign f1172_rst = rst;
  // Bindings to f1172

  // f1174
  logic [0:0] f1174_wen;
  logic [31:0] f1174_wdata;
  logic [0:0] f1174_clk;
  logic [0:0] f1174_rst;
  logic [31:0] f1174_rdata;
  sr_buffer_32_1 f1174(.wen(f1174_wen), .wdata(f1174_wdata), .clk(f1174_clk), .rst(f1174_rst), .rdata(f1174_rdata));
  assign f1174_clk = clk;
  assign f1174_rst = rst;
  // Bindings to f1174

  // f1176
  logic [0:0] f1176_wen;
  logic [31:0] f1176_wdata;
  logic [0:0] f1176_clk;
  logic [0:0] f1176_rst;
  logic [31:0] f1176_rdata;
  sr_buffer_32_1 f1176(.wen(f1176_wen), .wdata(f1176_wdata), .clk(f1176_clk), .rst(f1176_rst), .rdata(f1176_rdata));
  assign f1176_clk = clk;
  assign f1176_rst = rst;
  // Bindings to f1176

  // f1178
  logic [0:0] f1178_wen;
  logic [31:0] f1178_wdata;
  logic [0:0] f1178_clk;
  logic [0:0] f1178_rst;
  logic [31:0] f1178_rdata;
  sr_buffer_32_1 f1178(.wen(f1178_wen), .wdata(f1178_wdata), .clk(f1178_clk), .rst(f1178_rst), .rdata(f1178_rdata));
  assign f1178_clk = clk;
  assign f1178_rst = rst;
  // Bindings to f1178

  // f1180
  logic [0:0] f1180_wen;
  logic [31:0] f1180_wdata;
  logic [0:0] f1180_clk;
  logic [0:0] f1180_rst;
  logic [31:0] f1180_rdata;
  sr_buffer_32_1 f1180(.wen(f1180_wen), .wdata(f1180_wdata), .clk(f1180_clk), .rst(f1180_rst), .rdata(f1180_rdata));
  assign f1180_clk = clk;
  assign f1180_rst = rst;
  // Bindings to f1180

  // f1182
  logic [0:0] f1182_wen;
  logic [31:0] f1182_wdata;
  logic [0:0] f1182_clk;
  logic [0:0] f1182_rst;
  logic [31:0] f1182_rdata;
  sr_buffer_32_1 f1182(.wen(f1182_wen), .wdata(f1182_wdata), .clk(f1182_clk), .rst(f1182_rst), .rdata(f1182_rdata));
  assign f1182_clk = clk;
  assign f1182_rst = rst;
  // Bindings to f1182

  // f1184
  logic [0:0] f1184_wen;
  logic [31:0] f1184_wdata;
  logic [0:0] f1184_clk;
  logic [0:0] f1184_rst;
  logic [31:0] f1184_rdata;
  sr_buffer_32_1 f1184(.wen(f1184_wen), .wdata(f1184_wdata), .clk(f1184_clk), .rst(f1184_rst), .rdata(f1184_rdata));
  assign f1184_clk = clk;
  assign f1184_rst = rst;
  // Bindings to f1184

  // f1186
  logic [0:0] f1186_wen;
  logic [31:0] f1186_wdata;
  logic [0:0] f1186_clk;
  logic [0:0] f1186_rst;
  logic [31:0] f1186_rdata;
  sr_buffer_32_1 f1186(.wen(f1186_wen), .wdata(f1186_wdata), .clk(f1186_clk), .rst(f1186_rst), .rdata(f1186_rdata));
  assign f1186_clk = clk;
  assign f1186_rst = rst;
  // Bindings to f1186

  // f1188
  logic [0:0] f1188_wen;
  logic [31:0] f1188_wdata;
  logic [0:0] f1188_clk;
  logic [0:0] f1188_rst;
  logic [31:0] f1188_rdata;
  sr_buffer_32_1 f1188(.wen(f1188_wen), .wdata(f1188_wdata), .clk(f1188_clk), .rst(f1188_rst), .rdata(f1188_rdata));
  assign f1188_clk = clk;
  assign f1188_rst = rst;
  // Bindings to f1188

  // f1190
  logic [0:0] f1190_wen;
  logic [31:0] f1190_wdata;
  logic [0:0] f1190_clk;
  logic [0:0] f1190_rst;
  logic [31:0] f1190_rdata;
  sr_buffer_32_1 f1190(.wen(f1190_wen), .wdata(f1190_wdata), .clk(f1190_clk), .rst(f1190_rst), .rdata(f1190_rdata));
  assign f1190_clk = clk;
  assign f1190_rst = rst;
  // Bindings to f1190

  // f1192
  logic [0:0] f1192_wen;
  logic [31:0] f1192_wdata;
  logic [0:0] f1192_clk;
  logic [0:0] f1192_rst;
  logic [31:0] f1192_rdata;
  sr_buffer_32_1 f1192(.wen(f1192_wen), .wdata(f1192_wdata), .clk(f1192_clk), .rst(f1192_rst), .rdata(f1192_rdata));
  assign f1192_clk = clk;
  assign f1192_rst = rst;
  // Bindings to f1192

  // f1194
  logic [0:0] f1194_wen;
  logic [31:0] f1194_wdata;
  logic [0:0] f1194_clk;
  logic [0:0] f1194_rst;
  logic [31:0] f1194_rdata;
  sr_buffer_32_1 f1194(.wen(f1194_wen), .wdata(f1194_wdata), .clk(f1194_clk), .rst(f1194_rst), .rdata(f1194_rdata));
  assign f1194_clk = clk;
  assign f1194_rst = rst;
  // Bindings to f1194

  // f1196
  logic [0:0] f1196_wen;
  logic [31:0] f1196_wdata;
  logic [0:0] f1196_clk;
  logic [0:0] f1196_rst;
  logic [31:0] f1196_rdata;
  sr_buffer_32_1 f1196(.wen(f1196_wen), .wdata(f1196_wdata), .clk(f1196_clk), .rst(f1196_rst), .rdata(f1196_rdata));
  assign f1196_clk = clk;
  assign f1196_rst = rst;
  // Bindings to f1196

  // f1198
  logic [0:0] f1198_wen;
  logic [31:0] f1198_wdata;
  logic [0:0] f1198_clk;
  logic [0:0] f1198_rst;
  logic [31:0] f1198_rdata;
  sr_buffer_32_1 f1198(.wen(f1198_wen), .wdata(f1198_wdata), .clk(f1198_clk), .rst(f1198_rst), .rdata(f1198_rdata));
  assign f1198_clk = clk;
  assign f1198_rst = rst;
  // Bindings to f1198

  // f1200
  logic [0:0] f1200_wen;
  logic [31:0] f1200_wdata;
  logic [0:0] f1200_clk;
  logic [0:0] f1200_rst;
  logic [31:0] f1200_rdata;
  sr_buffer_32_1 f1200(.wen(f1200_wen), .wdata(f1200_wdata), .clk(f1200_clk), .rst(f1200_rst), .rdata(f1200_rdata));
  assign f1200_clk = clk;
  assign f1200_rst = rst;
  // Bindings to f1200

  // f1202
  logic [0:0] f1202_wen;
  logic [31:0] f1202_wdata;
  logic [0:0] f1202_clk;
  logic [0:0] f1202_rst;
  logic [31:0] f1202_rdata;
  sr_buffer_32_1 f1202(.wen(f1202_wen), .wdata(f1202_wdata), .clk(f1202_clk), .rst(f1202_rst), .rdata(f1202_rdata));
  assign f1202_clk = clk;
  assign f1202_rst = rst;
  // Bindings to f1202

  // f1204
  logic [0:0] f1204_wen;
  logic [31:0] f1204_wdata;
  logic [0:0] f1204_clk;
  logic [0:0] f1204_rst;
  logic [31:0] f1204_rdata;
  sr_buffer_32_1 f1204(.wen(f1204_wen), .wdata(f1204_wdata), .clk(f1204_clk), .rst(f1204_rst), .rdata(f1204_rdata));
  assign f1204_clk = clk;
  assign f1204_rst = rst;
  // Bindings to f1204

  // f1206
  logic [0:0] f1206_wen;
  logic [31:0] f1206_wdata;
  logic [0:0] f1206_clk;
  logic [0:0] f1206_rst;
  logic [31:0] f1206_rdata;
  sr_buffer_32_1 f1206(.wen(f1206_wen), .wdata(f1206_wdata), .clk(f1206_clk), .rst(f1206_rst), .rdata(f1206_rdata));
  assign f1206_clk = clk;
  assign f1206_rst = rst;
  // Bindings to f1206

  // f1208
  logic [0:0] f1208_wen;
  logic [31:0] f1208_wdata;
  logic [0:0] f1208_clk;
  logic [0:0] f1208_rst;
  logic [31:0] f1208_rdata;
  sr_buffer_32_1 f1208(.wen(f1208_wen), .wdata(f1208_wdata), .clk(f1208_clk), .rst(f1208_rst), .rdata(f1208_rdata));
  assign f1208_clk = clk;
  assign f1208_rst = rst;
  // Bindings to f1208

  // f1210
  logic [0:0] f1210_wen;
  logic [31:0] f1210_wdata;
  logic [0:0] f1210_clk;
  logic [0:0] f1210_rst;
  logic [31:0] f1210_rdata;
  sr_buffer_32_1 f1210(.wen(f1210_wen), .wdata(f1210_wdata), .clk(f1210_clk), .rst(f1210_rst), .rdata(f1210_rdata));
  assign f1210_clk = clk;
  assign f1210_rst = rst;
  // Bindings to f1210

  // f1212
  logic [0:0] f1212_wen;
  logic [31:0] f1212_wdata;
  logic [0:0] f1212_clk;
  logic [0:0] f1212_rst;
  logic [31:0] f1212_rdata;
  sr_buffer_32_1 f1212(.wen(f1212_wen), .wdata(f1212_wdata), .clk(f1212_clk), .rst(f1212_rst), .rdata(f1212_rdata));
  assign f1212_clk = clk;
  assign f1212_rst = rst;
  // Bindings to f1212

  // f1214
  logic [0:0] f1214_wen;
  logic [31:0] f1214_wdata;
  logic [0:0] f1214_clk;
  logic [0:0] f1214_rst;
  logic [31:0] f1214_rdata;
  sr_buffer_32_1 f1214(.wen(f1214_wen), .wdata(f1214_wdata), .clk(f1214_clk), .rst(f1214_rst), .rdata(f1214_rdata));
  assign f1214_clk = clk;
  assign f1214_rst = rst;
  // Bindings to f1214

  // f1216
  logic [0:0] f1216_wen;
  logic [31:0] f1216_wdata;
  logic [0:0] f1216_clk;
  logic [0:0] f1216_rst;
  logic [31:0] f1216_rdata;
  sr_buffer_32_1 f1216(.wen(f1216_wen), .wdata(f1216_wdata), .clk(f1216_clk), .rst(f1216_rst), .rdata(f1216_rdata));
  assign f1216_clk = clk;
  assign f1216_rst = rst;
  // Bindings to f1216

  // f1218
  logic [0:0] f1218_wen;
  logic [31:0] f1218_wdata;
  logic [0:0] f1218_clk;
  logic [0:0] f1218_rst;
  logic [31:0] f1218_rdata;
  sr_buffer_32_1 f1218(.wen(f1218_wen), .wdata(f1218_wdata), .clk(f1218_clk), .rst(f1218_rst), .rdata(f1218_rdata));
  assign f1218_clk = clk;
  assign f1218_rst = rst;
  // Bindings to f1218

  // f1220
  logic [0:0] f1220_wen;
  logic [31:0] f1220_wdata;
  logic [0:0] f1220_clk;
  logic [0:0] f1220_rst;
  logic [31:0] f1220_rdata;
  sr_buffer_32_1 f1220(.wen(f1220_wen), .wdata(f1220_wdata), .clk(f1220_clk), .rst(f1220_rst), .rdata(f1220_rdata));
  assign f1220_clk = clk;
  assign f1220_rst = rst;
  // Bindings to f1220

  // f1222
  logic [0:0] f1222_wen;
  logic [31:0] f1222_wdata;
  logic [0:0] f1222_clk;
  logic [0:0] f1222_rst;
  logic [31:0] f1222_rdata;
  sr_buffer_32_1 f1222(.wen(f1222_wen), .wdata(f1222_wdata), .clk(f1222_clk), .rst(f1222_rst), .rdata(f1222_rdata));
  assign f1222_clk = clk;
  assign f1222_rst = rst;
  // Bindings to f1222

  // f1224
  logic [0:0] f1224_wen;
  logic [31:0] f1224_wdata;
  logic [0:0] f1224_clk;
  logic [0:0] f1224_rst;
  logic [31:0] f1224_rdata;
  sr_buffer_32_1 f1224(.wen(f1224_wen), .wdata(f1224_wdata), .clk(f1224_clk), .rst(f1224_rst), .rdata(f1224_rdata));
  assign f1224_clk = clk;
  assign f1224_rst = rst;
  // Bindings to f1224

  // f1226
  logic [0:0] f1226_wen;
  logic [31:0] f1226_wdata;
  logic [0:0] f1226_clk;
  logic [0:0] f1226_rst;
  logic [31:0] f1226_rdata;
  sr_buffer_32_1 f1226(.wen(f1226_wen), .wdata(f1226_wdata), .clk(f1226_clk), .rst(f1226_rst), .rdata(f1226_rdata));
  assign f1226_clk = clk;
  assign f1226_rst = rst;
  // Bindings to f1226

  // f1228
  logic [0:0] f1228_wen;
  logic [31:0] f1228_wdata;
  logic [0:0] f1228_clk;
  logic [0:0] f1228_rst;
  logic [31:0] f1228_rdata;
  sr_buffer_32_1 f1228(.wen(f1228_wen), .wdata(f1228_wdata), .clk(f1228_clk), .rst(f1228_rst), .rdata(f1228_rdata));
  assign f1228_clk = clk;
  assign f1228_rst = rst;
  // Bindings to f1228

  // f1230
  logic [0:0] f1230_wen;
  logic [31:0] f1230_wdata;
  logic [0:0] f1230_clk;
  logic [0:0] f1230_rst;
  logic [31:0] f1230_rdata;
  sr_buffer_32_1 f1230(.wen(f1230_wen), .wdata(f1230_wdata), .clk(f1230_clk), .rst(f1230_rst), .rdata(f1230_rdata));
  assign f1230_clk = clk;
  assign f1230_rst = rst;
  // Bindings to f1230

  // f1232
  logic [0:0] f1232_wen;
  logic [31:0] f1232_wdata;
  logic [0:0] f1232_clk;
  logic [0:0] f1232_rst;
  logic [31:0] f1232_rdata;
  sr_buffer_32_1 f1232(.wen(f1232_wen), .wdata(f1232_wdata), .clk(f1232_clk), .rst(f1232_rst), .rdata(f1232_rdata));
  assign f1232_clk = clk;
  assign f1232_rst = rst;
  // Bindings to f1232

  // f1234
  logic [0:0] f1234_wen;
  logic [31:0] f1234_wdata;
  logic [0:0] f1234_clk;
  logic [0:0] f1234_rst;
  logic [31:0] f1234_rdata;
  sr_buffer_32_1 f1234(.wen(f1234_wen), .wdata(f1234_wdata), .clk(f1234_clk), .rst(f1234_rst), .rdata(f1234_rdata));
  assign f1234_clk = clk;
  assign f1234_rst = rst;
  // Bindings to f1234

  // f1236
  logic [0:0] f1236_wen;
  logic [31:0] f1236_wdata;
  logic [0:0] f1236_clk;
  logic [0:0] f1236_rst;
  logic [31:0] f1236_rdata;
  sr_buffer_32_1 f1236(.wen(f1236_wen), .wdata(f1236_wdata), .clk(f1236_clk), .rst(f1236_rst), .rdata(f1236_rdata));
  assign f1236_clk = clk;
  assign f1236_rst = rst;
  // Bindings to f1236

  // f1238
  logic [0:0] f1238_wen;
  logic [31:0] f1238_wdata;
  logic [0:0] f1238_clk;
  logic [0:0] f1238_rst;
  logic [31:0] f1238_rdata;
  sr_buffer_32_1 f1238(.wen(f1238_wen), .wdata(f1238_wdata), .clk(f1238_clk), .rst(f1238_rst), .rdata(f1238_rdata));
  assign f1238_clk = clk;
  assign f1238_rst = rst;
  // Bindings to f1238

  // f1240
  logic [0:0] f1240_wen;
  logic [31:0] f1240_wdata;
  logic [0:0] f1240_clk;
  logic [0:0] f1240_rst;
  logic [31:0] f1240_rdata;
  sr_buffer_32_1 f1240(.wen(f1240_wen), .wdata(f1240_wdata), .clk(f1240_clk), .rst(f1240_rst), .rdata(f1240_rdata));
  assign f1240_clk = clk;
  assign f1240_rst = rst;
  // Bindings to f1240

  // f1242
  logic [0:0] f1242_wen;
  logic [31:0] f1242_wdata;
  logic [0:0] f1242_clk;
  logic [0:0] f1242_rst;
  logic [31:0] f1242_rdata;
  sr_buffer_32_1 f1242(.wen(f1242_wen), .wdata(f1242_wdata), .clk(f1242_clk), .rst(f1242_rst), .rdata(f1242_rdata));
  assign f1242_clk = clk;
  assign f1242_rst = rst;
  // Bindings to f1242

  // f1244
  logic [0:0] f1244_wen;
  logic [31:0] f1244_wdata;
  logic [0:0] f1244_clk;
  logic [0:0] f1244_rst;
  logic [31:0] f1244_rdata;
  sr_buffer_32_1 f1244(.wen(f1244_wen), .wdata(f1244_wdata), .clk(f1244_clk), .rst(f1244_rst), .rdata(f1244_rdata));
  assign f1244_clk = clk;
  assign f1244_rst = rst;
  // Bindings to f1244

  // f1246
  logic [0:0] f1246_wen;
  logic [31:0] f1246_wdata;
  logic [0:0] f1246_clk;
  logic [0:0] f1246_rst;
  logic [31:0] f1246_rdata;
  sr_buffer_32_1 f1246(.wen(f1246_wen), .wdata(f1246_wdata), .clk(f1246_clk), .rst(f1246_rst), .rdata(f1246_rdata));
  assign f1246_clk = clk;
  assign f1246_rst = rst;
  // Bindings to f1246

  // f1248
  logic [0:0] f1248_wen;
  logic [31:0] f1248_wdata;
  logic [0:0] f1248_clk;
  logic [0:0] f1248_rst;
  logic [31:0] f1248_rdata;
  sr_buffer_32_1 f1248(.wen(f1248_wen), .wdata(f1248_wdata), .clk(f1248_clk), .rst(f1248_rst), .rdata(f1248_rdata));
  assign f1248_clk = clk;
  assign f1248_rst = rst;
  // Bindings to f1248

  // f1250
  logic [0:0] f1250_wen;
  logic [31:0] f1250_wdata;
  logic [0:0] f1250_clk;
  logic [0:0] f1250_rst;
  logic [31:0] f1250_rdata;
  sr_buffer_32_1 f1250(.wen(f1250_wen), .wdata(f1250_wdata), .clk(f1250_clk), .rst(f1250_rst), .rdata(f1250_rdata));
  assign f1250_clk = clk;
  assign f1250_rst = rst;
  // Bindings to f1250

  // f1252
  logic [0:0] f1252_wen;
  logic [31:0] f1252_wdata;
  logic [0:0] f1252_clk;
  logic [0:0] f1252_rst;
  logic [31:0] f1252_rdata;
  sr_buffer_32_1 f1252(.wen(f1252_wen), .wdata(f1252_wdata), .clk(f1252_clk), .rst(f1252_rst), .rdata(f1252_rdata));
  assign f1252_clk = clk;
  assign f1252_rst = rst;
  // Bindings to f1252

  // f1254
  logic [0:0] f1254_wen;
  logic [31:0] f1254_wdata;
  logic [0:0] f1254_clk;
  logic [0:0] f1254_rst;
  logic [31:0] f1254_rdata;
  sr_buffer_32_1 f1254(.wen(f1254_wen), .wdata(f1254_wdata), .clk(f1254_clk), .rst(f1254_rst), .rdata(f1254_rdata));
  assign f1254_clk = clk;
  assign f1254_rst = rst;
  // Bindings to f1254

  // f1256
  logic [0:0] f1256_wen;
  logic [31:0] f1256_wdata;
  logic [0:0] f1256_clk;
  logic [0:0] f1256_rst;
  logic [31:0] f1256_rdata;
  sr_buffer_32_1 f1256(.wen(f1256_wen), .wdata(f1256_wdata), .clk(f1256_clk), .rst(f1256_rst), .rdata(f1256_rdata));
  assign f1256_clk = clk;
  assign f1256_rst = rst;
  // Bindings to f1256

  // f1258
  logic [0:0] f1258_wen;
  logic [31:0] f1258_wdata;
  logic [0:0] f1258_clk;
  logic [0:0] f1258_rst;
  logic [31:0] f1258_rdata;
  sr_buffer_32_1 f1258(.wen(f1258_wen), .wdata(f1258_wdata), .clk(f1258_clk), .rst(f1258_rst), .rdata(f1258_rdata));
  assign f1258_clk = clk;
  assign f1258_rst = rst;
  // Bindings to f1258

  // f1260
  logic [0:0] f1260_wen;
  logic [31:0] f1260_wdata;
  logic [0:0] f1260_clk;
  logic [0:0] f1260_rst;
  logic [31:0] f1260_rdata;
  sr_buffer_32_1 f1260(.wen(f1260_wen), .wdata(f1260_wdata), .clk(f1260_clk), .rst(f1260_rst), .rdata(f1260_rdata));
  assign f1260_clk = clk;
  assign f1260_rst = rst;
  // Bindings to f1260

  // f1262
  logic [0:0] f1262_wen;
  logic [31:0] f1262_wdata;
  logic [0:0] f1262_clk;
  logic [0:0] f1262_rst;
  logic [31:0] f1262_rdata;
  sr_buffer_32_1 f1262(.wen(f1262_wen), .wdata(f1262_wdata), .clk(f1262_clk), .rst(f1262_rst), .rdata(f1262_rdata));
  assign f1262_clk = clk;
  assign f1262_rst = rst;
  // Bindings to f1262

  // f1264
  logic [0:0] f1264_wen;
  logic [31:0] f1264_wdata;
  logic [0:0] f1264_clk;
  logic [0:0] f1264_rst;
  logic [31:0] f1264_rdata;
  sr_buffer_32_1 f1264(.wen(f1264_wen), .wdata(f1264_wdata), .clk(f1264_clk), .rst(f1264_rst), .rdata(f1264_rdata));
  assign f1264_clk = clk;
  assign f1264_rst = rst;
  // Bindings to f1264

  // f1266
  logic [0:0] f1266_wen;
  logic [31:0] f1266_wdata;
  logic [0:0] f1266_clk;
  logic [0:0] f1266_rst;
  logic [31:0] f1266_rdata;
  sr_buffer_32_1 f1266(.wen(f1266_wen), .wdata(f1266_wdata), .clk(f1266_clk), .rst(f1266_rst), .rdata(f1266_rdata));
  assign f1266_clk = clk;
  assign f1266_rst = rst;
  // Bindings to f1266

  // f1268
  logic [0:0] f1268_wen;
  logic [31:0] f1268_wdata;
  logic [0:0] f1268_clk;
  logic [0:0] f1268_rst;
  logic [31:0] f1268_rdata;
  sr_buffer_32_1 f1268(.wen(f1268_wen), .wdata(f1268_wdata), .clk(f1268_clk), .rst(f1268_rst), .rdata(f1268_rdata));
  assign f1268_clk = clk;
  assign f1268_rst = rst;
  // Bindings to f1268

  // f1270
  logic [0:0] f1270_wen;
  logic [31:0] f1270_wdata;
  logic [0:0] f1270_clk;
  logic [0:0] f1270_rst;
  logic [31:0] f1270_rdata;
  sr_buffer_32_1 f1270(.wen(f1270_wen), .wdata(f1270_wdata), .clk(f1270_clk), .rst(f1270_rst), .rdata(f1270_rdata));
  assign f1270_clk = clk;
  assign f1270_rst = rst;
  // Bindings to f1270

  // f1272
  logic [0:0] f1272_wen;
  logic [31:0] f1272_wdata;
  logic [0:0] f1272_clk;
  logic [0:0] f1272_rst;
  logic [31:0] f1272_rdata;
  sr_buffer_32_1 f1272(.wen(f1272_wen), .wdata(f1272_wdata), .clk(f1272_clk), .rst(f1272_rst), .rdata(f1272_rdata));
  assign f1272_clk = clk;
  assign f1272_rst = rst;
  // Bindings to f1272

  // f1274
  logic [0:0] f1274_wen;
  logic [31:0] f1274_wdata;
  logic [0:0] f1274_clk;
  logic [0:0] f1274_rst;
  logic [31:0] f1274_rdata;
  sr_buffer_32_1 f1274(.wen(f1274_wen), .wdata(f1274_wdata), .clk(f1274_clk), .rst(f1274_rst), .rdata(f1274_rdata));
  assign f1274_clk = clk;
  assign f1274_rst = rst;
  // Bindings to f1274

  // f1276
  logic [0:0] f1276_wen;
  logic [31:0] f1276_wdata;
  logic [0:0] f1276_clk;
  logic [0:0] f1276_rst;
  logic [31:0] f1276_rdata;
  sr_buffer_32_1 f1276(.wen(f1276_wen), .wdata(f1276_wdata), .clk(f1276_clk), .rst(f1276_rst), .rdata(f1276_rdata));
  assign f1276_clk = clk;
  assign f1276_rst = rst;
  // Bindings to f1276

  // f1278
  logic [0:0] f1278_wen;
  logic [31:0] f1278_wdata;
  logic [0:0] f1278_clk;
  logic [0:0] f1278_rst;
  logic [31:0] f1278_rdata;
  sr_buffer_32_1 f1278(.wen(f1278_wen), .wdata(f1278_wdata), .clk(f1278_clk), .rst(f1278_rst), .rdata(f1278_rdata));
  assign f1278_clk = clk;
  assign f1278_rst = rst;
  // Bindings to f1278

  // f1280
  logic [0:0] f1280_wen;
  logic [31:0] f1280_wdata;
  logic [0:0] f1280_clk;
  logic [0:0] f1280_rst;
  logic [31:0] f1280_rdata;
  sr_buffer_32_1 f1280(.wen(f1280_wen), .wdata(f1280_wdata), .clk(f1280_clk), .rst(f1280_rst), .rdata(f1280_rdata));
  assign f1280_clk = clk;
  assign f1280_rst = rst;
  // Bindings to f1280

  // f1282
  logic [0:0] f1282_wen;
  logic [31:0] f1282_wdata;
  logic [0:0] f1282_clk;
  logic [0:0] f1282_rst;
  logic [31:0] f1282_rdata;
  sr_buffer_32_1 f1282(.wen(f1282_wen), .wdata(f1282_wdata), .clk(f1282_clk), .rst(f1282_rst), .rdata(f1282_rdata));
  assign f1282_clk = clk;
  assign f1282_rst = rst;
  // Bindings to f1282

  // f1284
  logic [0:0] f1284_wen;
  logic [31:0] f1284_wdata;
  logic [0:0] f1284_clk;
  logic [0:0] f1284_rst;
  logic [31:0] f1284_rdata;
  sr_buffer_32_1 f1284(.wen(f1284_wen), .wdata(f1284_wdata), .clk(f1284_clk), .rst(f1284_rst), .rdata(f1284_rdata));
  assign f1284_clk = clk;
  assign f1284_rst = rst;
  // Bindings to f1284

  // f1286
  logic [0:0] f1286_wen;
  logic [31:0] f1286_wdata;
  logic [0:0] f1286_clk;
  logic [0:0] f1286_rst;
  logic [31:0] f1286_rdata;
  sr_buffer_32_1 f1286(.wen(f1286_wen), .wdata(f1286_wdata), .clk(f1286_clk), .rst(f1286_rst), .rdata(f1286_rdata));
  assign f1286_clk = clk;
  assign f1286_rst = rst;
  // Bindings to f1286

  // f1288
  logic [0:0] f1288_wen;
  logic [31:0] f1288_wdata;
  logic [0:0] f1288_clk;
  logic [0:0] f1288_rst;
  logic [31:0] f1288_rdata;
  sr_buffer_32_1 f1288(.wen(f1288_wen), .wdata(f1288_wdata), .clk(f1288_clk), .rst(f1288_rst), .rdata(f1288_rdata));
  assign f1288_clk = clk;
  assign f1288_rst = rst;
  // Bindings to f1288

  // f1290
  logic [0:0] f1290_wen;
  logic [31:0] f1290_wdata;
  logic [0:0] f1290_clk;
  logic [0:0] f1290_rst;
  logic [31:0] f1290_rdata;
  sr_buffer_32_1 f1290(.wen(f1290_wen), .wdata(f1290_wdata), .clk(f1290_clk), .rst(f1290_rst), .rdata(f1290_rdata));
  assign f1290_clk = clk;
  assign f1290_rst = rst;
  // Bindings to f1290

  // f1292
  logic [0:0] f1292_wen;
  logic [31:0] f1292_wdata;
  logic [0:0] f1292_clk;
  logic [0:0] f1292_rst;
  logic [31:0] f1292_rdata;
  sr_buffer_32_1 f1292(.wen(f1292_wen), .wdata(f1292_wdata), .clk(f1292_clk), .rst(f1292_rst), .rdata(f1292_rdata));
  assign f1292_clk = clk;
  assign f1292_rst = rst;
  // Bindings to f1292

  // f1294
  logic [0:0] f1294_wen;
  logic [31:0] f1294_wdata;
  logic [0:0] f1294_clk;
  logic [0:0] f1294_rst;
  logic [31:0] f1294_rdata;
  sr_buffer_32_1 f1294(.wen(f1294_wen), .wdata(f1294_wdata), .clk(f1294_clk), .rst(f1294_rst), .rdata(f1294_rdata));
  assign f1294_clk = clk;
  assign f1294_rst = rst;
  // Bindings to f1294

  // f1296
  logic [0:0] f1296_wen;
  logic [31:0] f1296_wdata;
  logic [0:0] f1296_clk;
  logic [0:0] f1296_rst;
  logic [31:0] f1296_rdata;
  sr_buffer_32_1 f1296(.wen(f1296_wen), .wdata(f1296_wdata), .clk(f1296_clk), .rst(f1296_rst), .rdata(f1296_rdata));
  assign f1296_clk = clk;
  assign f1296_rst = rst;
  // Bindings to f1296

  // f1298
  logic [0:0] f1298_wen;
  logic [31:0] f1298_wdata;
  logic [0:0] f1298_clk;
  logic [0:0] f1298_rst;
  logic [31:0] f1298_rdata;
  sr_buffer_32_1 f1298(.wen(f1298_wen), .wdata(f1298_wdata), .clk(f1298_clk), .rst(f1298_rst), .rdata(f1298_rdata));
  assign f1298_clk = clk;
  assign f1298_rst = rst;
  // Bindings to f1298

  // f1300
  logic [0:0] f1300_wen;
  logic [31:0] f1300_wdata;
  logic [0:0] f1300_clk;
  logic [0:0] f1300_rst;
  logic [31:0] f1300_rdata;
  sr_buffer_32_1 f1300(.wen(f1300_wen), .wdata(f1300_wdata), .clk(f1300_clk), .rst(f1300_rst), .rdata(f1300_rdata));
  assign f1300_clk = clk;
  assign f1300_rst = rst;
  // Bindings to f1300

  // f1302
  logic [0:0] f1302_wen;
  logic [31:0] f1302_wdata;
  logic [0:0] f1302_clk;
  logic [0:0] f1302_rst;
  logic [31:0] f1302_rdata;
  sr_buffer_32_1 f1302(.wen(f1302_wen), .wdata(f1302_wdata), .clk(f1302_clk), .rst(f1302_rst), .rdata(f1302_rdata));
  assign f1302_clk = clk;
  assign f1302_rst = rst;
  // Bindings to f1302

  // f1304
  logic [0:0] f1304_wen;
  logic [31:0] f1304_wdata;
  logic [0:0] f1304_clk;
  logic [0:0] f1304_rst;
  logic [31:0] f1304_rdata;
  sr_buffer_32_1 f1304(.wen(f1304_wen), .wdata(f1304_wdata), .clk(f1304_clk), .rst(f1304_rst), .rdata(f1304_rdata));
  assign f1304_clk = clk;
  assign f1304_rst = rst;
  // Bindings to f1304

  // f1306
  logic [0:0] f1306_wen;
  logic [31:0] f1306_wdata;
  logic [0:0] f1306_clk;
  logic [0:0] f1306_rst;
  logic [31:0] f1306_rdata;
  sr_buffer_32_1 f1306(.wen(f1306_wen), .wdata(f1306_wdata), .clk(f1306_clk), .rst(f1306_rst), .rdata(f1306_rdata));
  assign f1306_clk = clk;
  assign f1306_rst = rst;
  // Bindings to f1306

  // f1308
  logic [0:0] f1308_wen;
  logic [31:0] f1308_wdata;
  logic [0:0] f1308_clk;
  logic [0:0] f1308_rst;
  logic [31:0] f1308_rdata;
  sr_buffer_32_1 f1308(.wen(f1308_wen), .wdata(f1308_wdata), .clk(f1308_clk), .rst(f1308_rst), .rdata(f1308_rdata));
  assign f1308_clk = clk;
  assign f1308_rst = rst;
  // Bindings to f1308

  // f1310
  logic [0:0] f1310_wen;
  logic [31:0] f1310_wdata;
  logic [0:0] f1310_clk;
  logic [0:0] f1310_rst;
  logic [31:0] f1310_rdata;
  sr_buffer_32_1 f1310(.wen(f1310_wen), .wdata(f1310_wdata), .clk(f1310_clk), .rst(f1310_rst), .rdata(f1310_rdata));
  assign f1310_clk = clk;
  assign f1310_rst = rst;
  // Bindings to f1310

  // f1312
  logic [0:0] f1312_wen;
  logic [31:0] f1312_wdata;
  logic [0:0] f1312_clk;
  logic [0:0] f1312_rst;
  logic [31:0] f1312_rdata;
  sr_buffer_32_1 f1312(.wen(f1312_wen), .wdata(f1312_wdata), .clk(f1312_clk), .rst(f1312_rst), .rdata(f1312_rdata));
  assign f1312_clk = clk;
  assign f1312_rst = rst;
  // Bindings to f1312

  // f1314
  logic [0:0] f1314_wen;
  logic [31:0] f1314_wdata;
  logic [0:0] f1314_clk;
  logic [0:0] f1314_rst;
  logic [31:0] f1314_rdata;
  sr_buffer_32_1 f1314(.wen(f1314_wen), .wdata(f1314_wdata), .clk(f1314_clk), .rst(f1314_rst), .rdata(f1314_rdata));
  assign f1314_clk = clk;
  assign f1314_rst = rst;
  // Bindings to f1314

  // f1316
  logic [0:0] f1316_wen;
  logic [31:0] f1316_wdata;
  logic [0:0] f1316_clk;
  logic [0:0] f1316_rst;
  logic [31:0] f1316_rdata;
  sr_buffer_32_1 f1316(.wen(f1316_wen), .wdata(f1316_wdata), .clk(f1316_clk), .rst(f1316_rst), .rdata(f1316_rdata));
  assign f1316_clk = clk;
  assign f1316_rst = rst;
  // Bindings to f1316

  // f1318
  logic [0:0] f1318_wen;
  logic [31:0] f1318_wdata;
  logic [0:0] f1318_clk;
  logic [0:0] f1318_rst;
  logic [31:0] f1318_rdata;
  sr_buffer_32_1 f1318(.wen(f1318_wen), .wdata(f1318_wdata), .clk(f1318_clk), .rst(f1318_rst), .rdata(f1318_rdata));
  assign f1318_clk = clk;
  assign f1318_rst = rst;
  // Bindings to f1318

  // f1320
  logic [0:0] f1320_wen;
  logic [31:0] f1320_wdata;
  logic [0:0] f1320_clk;
  logic [0:0] f1320_rst;
  logic [31:0] f1320_rdata;
  sr_buffer_32_1 f1320(.wen(f1320_wen), .wdata(f1320_wdata), .clk(f1320_clk), .rst(f1320_rst), .rdata(f1320_rdata));
  assign f1320_clk = clk;
  assign f1320_rst = rst;
  // Bindings to f1320

  // f1322
  logic [0:0] f1322_wen;
  logic [31:0] f1322_wdata;
  logic [0:0] f1322_clk;
  logic [0:0] f1322_rst;
  logic [31:0] f1322_rdata;
  sr_buffer_32_1 f1322(.wen(f1322_wen), .wdata(f1322_wdata), .clk(f1322_clk), .rst(f1322_rst), .rdata(f1322_rdata));
  assign f1322_clk = clk;
  assign f1322_rst = rst;
  // Bindings to f1322

  // f1324
  logic [0:0] f1324_wen;
  logic [31:0] f1324_wdata;
  logic [0:0] f1324_clk;
  logic [0:0] f1324_rst;
  logic [31:0] f1324_rdata;
  sr_buffer_32_1 f1324(.wen(f1324_wen), .wdata(f1324_wdata), .clk(f1324_clk), .rst(f1324_rst), .rdata(f1324_rdata));
  assign f1324_clk = clk;
  assign f1324_rst = rst;
  // Bindings to f1324

  // f1326
  logic [0:0] f1326_wen;
  logic [31:0] f1326_wdata;
  logic [0:0] f1326_clk;
  logic [0:0] f1326_rst;
  logic [31:0] f1326_rdata;
  sr_buffer_32_1 f1326(.wen(f1326_wen), .wdata(f1326_wdata), .clk(f1326_clk), .rst(f1326_rst), .rdata(f1326_rdata));
  assign f1326_clk = clk;
  assign f1326_rst = rst;
  // Bindings to f1326

  // f1328
  logic [0:0] f1328_wen;
  logic [31:0] f1328_wdata;
  logic [0:0] f1328_clk;
  logic [0:0] f1328_rst;
  logic [31:0] f1328_rdata;
  sr_buffer_32_1 f1328(.wen(f1328_wen), .wdata(f1328_wdata), .clk(f1328_clk), .rst(f1328_rst), .rdata(f1328_rdata));
  assign f1328_clk = clk;
  assign f1328_rst = rst;
  // Bindings to f1328

  // f1330
  logic [0:0] f1330_wen;
  logic [31:0] f1330_wdata;
  logic [0:0] f1330_clk;
  logic [0:0] f1330_rst;
  logic [31:0] f1330_rdata;
  sr_buffer_32_1 f1330(.wen(f1330_wen), .wdata(f1330_wdata), .clk(f1330_clk), .rst(f1330_rst), .rdata(f1330_rdata));
  assign f1330_clk = clk;
  assign f1330_rst = rst;
  // Bindings to f1330

  // f1332
  logic [0:0] f1332_wen;
  logic [31:0] f1332_wdata;
  logic [0:0] f1332_clk;
  logic [0:0] f1332_rst;
  logic [31:0] f1332_rdata;
  sr_buffer_32_1 f1332(.wen(f1332_wen), .wdata(f1332_wdata), .clk(f1332_clk), .rst(f1332_rst), .rdata(f1332_rdata));
  assign f1332_clk = clk;
  assign f1332_rst = rst;
  // Bindings to f1332

  // f1334
  logic [0:0] f1334_wen;
  logic [31:0] f1334_wdata;
  logic [0:0] f1334_clk;
  logic [0:0] f1334_rst;
  logic [31:0] f1334_rdata;
  sr_buffer_32_1 f1334(.wen(f1334_wen), .wdata(f1334_wdata), .clk(f1334_clk), .rst(f1334_rst), .rdata(f1334_rdata));
  assign f1334_clk = clk;
  assign f1334_rst = rst;
  // Bindings to f1334

  // f1336
  logic [0:0] f1336_wen;
  logic [31:0] f1336_wdata;
  logic [0:0] f1336_clk;
  logic [0:0] f1336_rst;
  logic [31:0] f1336_rdata;
  sr_buffer_32_1 f1336(.wen(f1336_wen), .wdata(f1336_wdata), .clk(f1336_clk), .rst(f1336_rst), .rdata(f1336_rdata));
  assign f1336_clk = clk;
  assign f1336_rst = rst;
  // Bindings to f1336

  // f1338
  logic [0:0] f1338_wen;
  logic [31:0] f1338_wdata;
  logic [0:0] f1338_clk;
  logic [0:0] f1338_rst;
  logic [31:0] f1338_rdata;
  sr_buffer_32_1 f1338(.wen(f1338_wen), .wdata(f1338_wdata), .clk(f1338_clk), .rst(f1338_rst), .rdata(f1338_rdata));
  assign f1338_clk = clk;
  assign f1338_rst = rst;
  // Bindings to f1338

  // f1340
  logic [0:0] f1340_wen;
  logic [31:0] f1340_wdata;
  logic [0:0] f1340_clk;
  logic [0:0] f1340_rst;
  logic [31:0] f1340_rdata;
  sr_buffer_32_1 f1340(.wen(f1340_wen), .wdata(f1340_wdata), .clk(f1340_clk), .rst(f1340_rst), .rdata(f1340_rdata));
  assign f1340_clk = clk;
  assign f1340_rst = rst;
  // Bindings to f1340

  // f1342
  logic [0:0] f1342_wen;
  logic [31:0] f1342_wdata;
  logic [0:0] f1342_clk;
  logic [0:0] f1342_rst;
  logic [31:0] f1342_rdata;
  sr_buffer_32_1 f1342(.wen(f1342_wen), .wdata(f1342_wdata), .clk(f1342_clk), .rst(f1342_rst), .rdata(f1342_rdata));
  assign f1342_clk = clk;
  assign f1342_rst = rst;
  // Bindings to f1342

  // f1344
  logic [0:0] f1344_wen;
  logic [31:0] f1344_wdata;
  logic [0:0] f1344_clk;
  logic [0:0] f1344_rst;
  logic [31:0] f1344_rdata;
  sr_buffer_32_1 f1344(.wen(f1344_wen), .wdata(f1344_wdata), .clk(f1344_clk), .rst(f1344_rst), .rdata(f1344_rdata));
  assign f1344_clk = clk;
  assign f1344_rst = rst;
  // Bindings to f1344

  // f1346
  logic [0:0] f1346_wen;
  logic [31:0] f1346_wdata;
  logic [0:0] f1346_clk;
  logic [0:0] f1346_rst;
  logic [31:0] f1346_rdata;
  sr_buffer_32_1 f1346(.wen(f1346_wen), .wdata(f1346_wdata), .clk(f1346_clk), .rst(f1346_rst), .rdata(f1346_rdata));
  assign f1346_clk = clk;
  assign f1346_rst = rst;
  // Bindings to f1346

  // f1348
  logic [0:0] f1348_wen;
  logic [31:0] f1348_wdata;
  logic [0:0] f1348_clk;
  logic [0:0] f1348_rst;
  logic [31:0] f1348_rdata;
  sr_buffer_32_1 f1348(.wen(f1348_wen), .wdata(f1348_wdata), .clk(f1348_clk), .rst(f1348_rst), .rdata(f1348_rdata));
  assign f1348_clk = clk;
  assign f1348_rst = rst;
  // Bindings to f1348

  // f1350
  logic [0:0] f1350_wen;
  logic [31:0] f1350_wdata;
  logic [0:0] f1350_clk;
  logic [0:0] f1350_rst;
  logic [31:0] f1350_rdata;
  sr_buffer_32_1 f1350(.wen(f1350_wen), .wdata(f1350_wdata), .clk(f1350_clk), .rst(f1350_rst), .rdata(f1350_rdata));
  assign f1350_clk = clk;
  assign f1350_rst = rst;
  // Bindings to f1350

  // f1352
  logic [0:0] f1352_wen;
  logic [31:0] f1352_wdata;
  logic [0:0] f1352_clk;
  logic [0:0] f1352_rst;
  logic [31:0] f1352_rdata;
  sr_buffer_32_1 f1352(.wen(f1352_wen), .wdata(f1352_wdata), .clk(f1352_clk), .rst(f1352_rst), .rdata(f1352_rdata));
  assign f1352_clk = clk;
  assign f1352_rst = rst;
  // Bindings to f1352

  // f1354
  logic [0:0] f1354_wen;
  logic [31:0] f1354_wdata;
  logic [0:0] f1354_clk;
  logic [0:0] f1354_rst;
  logic [31:0] f1354_rdata;
  sr_buffer_32_1 f1354(.wen(f1354_wen), .wdata(f1354_wdata), .clk(f1354_clk), .rst(f1354_rst), .rdata(f1354_rdata));
  assign f1354_clk = clk;
  assign f1354_rst = rst;
  // Bindings to f1354

  // f1356
  logic [0:0] f1356_wen;
  logic [31:0] f1356_wdata;
  logic [0:0] f1356_clk;
  logic [0:0] f1356_rst;
  logic [31:0] f1356_rdata;
  sr_buffer_32_1 f1356(.wen(f1356_wen), .wdata(f1356_wdata), .clk(f1356_clk), .rst(f1356_rst), .rdata(f1356_rdata));
  assign f1356_clk = clk;
  assign f1356_rst = rst;
  // Bindings to f1356

  // f1358
  logic [0:0] f1358_wen;
  logic [31:0] f1358_wdata;
  logic [0:0] f1358_clk;
  logic [0:0] f1358_rst;
  logic [31:0] f1358_rdata;
  sr_buffer_32_1 f1358(.wen(f1358_wen), .wdata(f1358_wdata), .clk(f1358_clk), .rst(f1358_rst), .rdata(f1358_rdata));
  assign f1358_clk = clk;
  assign f1358_rst = rst;
  // Bindings to f1358

  // f1360
  logic [0:0] f1360_wen;
  logic [31:0] f1360_wdata;
  logic [0:0] f1360_clk;
  logic [0:0] f1360_rst;
  logic [31:0] f1360_rdata;
  sr_buffer_32_1 f1360(.wen(f1360_wen), .wdata(f1360_wdata), .clk(f1360_clk), .rst(f1360_rst), .rdata(f1360_rdata));
  assign f1360_clk = clk;
  assign f1360_rst = rst;
  // Bindings to f1360

  // f1362
  logic [0:0] f1362_wen;
  logic [31:0] f1362_wdata;
  logic [0:0] f1362_clk;
  logic [0:0] f1362_rst;
  logic [31:0] f1362_rdata;
  sr_buffer_32_1 f1362(.wen(f1362_wen), .wdata(f1362_wdata), .clk(f1362_clk), .rst(f1362_rst), .rdata(f1362_rdata));
  assign f1362_clk = clk;
  assign f1362_rst = rst;
  // Bindings to f1362

  // f1364
  logic [0:0] f1364_wen;
  logic [31:0] f1364_wdata;
  logic [0:0] f1364_clk;
  logic [0:0] f1364_rst;
  logic [31:0] f1364_rdata;
  sr_buffer_32_1 f1364(.wen(f1364_wen), .wdata(f1364_wdata), .clk(f1364_clk), .rst(f1364_rst), .rdata(f1364_rdata));
  assign f1364_clk = clk;
  assign f1364_rst = rst;
  // Bindings to f1364

  // f1366
  logic [0:0] f1366_wen;
  logic [31:0] f1366_wdata;
  logic [0:0] f1366_clk;
  logic [0:0] f1366_rst;
  logic [31:0] f1366_rdata;
  sr_buffer_32_1 f1366(.wen(f1366_wen), .wdata(f1366_wdata), .clk(f1366_clk), .rst(f1366_rst), .rdata(f1366_rdata));
  assign f1366_clk = clk;
  assign f1366_rst = rst;
  // Bindings to f1366

  // f1368
  logic [0:0] f1368_wen;
  logic [31:0] f1368_wdata;
  logic [0:0] f1368_clk;
  logic [0:0] f1368_rst;
  logic [31:0] f1368_rdata;
  sr_buffer_32_1 f1368(.wen(f1368_wen), .wdata(f1368_wdata), .clk(f1368_clk), .rst(f1368_rst), .rdata(f1368_rdata));
  assign f1368_clk = clk;
  assign f1368_rst = rst;
  // Bindings to f1368

  // f1370
  logic [0:0] f1370_wen;
  logic [31:0] f1370_wdata;
  logic [0:0] f1370_clk;
  logic [0:0] f1370_rst;
  logic [31:0] f1370_rdata;
  sr_buffer_32_1 f1370(.wen(f1370_wen), .wdata(f1370_wdata), .clk(f1370_clk), .rst(f1370_rst), .rdata(f1370_rdata));
  assign f1370_clk = clk;
  assign f1370_rst = rst;
  // Bindings to f1370

  // f1372
  logic [0:0] f1372_wen;
  logic [31:0] f1372_wdata;
  logic [0:0] f1372_clk;
  logic [0:0] f1372_rst;
  logic [31:0] f1372_rdata;
  sr_buffer_32_1 f1372(.wen(f1372_wen), .wdata(f1372_wdata), .clk(f1372_clk), .rst(f1372_rst), .rdata(f1372_rdata));
  assign f1372_clk = clk;
  assign f1372_rst = rst;
  // Bindings to f1372

  // f1374
  logic [0:0] f1374_wen;
  logic [31:0] f1374_wdata;
  logic [0:0] f1374_clk;
  logic [0:0] f1374_rst;
  logic [31:0] f1374_rdata;
  sr_buffer_32_1 f1374(.wen(f1374_wen), .wdata(f1374_wdata), .clk(f1374_clk), .rst(f1374_rst), .rdata(f1374_rdata));
  assign f1374_clk = clk;
  assign f1374_rst = rst;
  // Bindings to f1374

  // f1376
  logic [0:0] f1376_wen;
  logic [31:0] f1376_wdata;
  logic [0:0] f1376_clk;
  logic [0:0] f1376_rst;
  logic [31:0] f1376_rdata;
  sr_buffer_32_1 f1376(.wen(f1376_wen), .wdata(f1376_wdata), .clk(f1376_clk), .rst(f1376_rst), .rdata(f1376_rdata));
  assign f1376_clk = clk;
  assign f1376_rst = rst;
  // Bindings to f1376

  // f1378
  logic [0:0] f1378_wen;
  logic [31:0] f1378_wdata;
  logic [0:0] f1378_clk;
  logic [0:0] f1378_rst;
  logic [31:0] f1378_rdata;
  sr_buffer_32_1 f1378(.wen(f1378_wen), .wdata(f1378_wdata), .clk(f1378_clk), .rst(f1378_rst), .rdata(f1378_rdata));
  assign f1378_clk = clk;
  assign f1378_rst = rst;
  // Bindings to f1378

  // f1380
  logic [0:0] f1380_wen;
  logic [31:0] f1380_wdata;
  logic [0:0] f1380_clk;
  logic [0:0] f1380_rst;
  logic [31:0] f1380_rdata;
  sr_buffer_32_1 f1380(.wen(f1380_wen), .wdata(f1380_wdata), .clk(f1380_clk), .rst(f1380_rst), .rdata(f1380_rdata));
  assign f1380_clk = clk;
  assign f1380_rst = rst;
  // Bindings to f1380

  // f1382
  logic [0:0] f1382_wen;
  logic [31:0] f1382_wdata;
  logic [0:0] f1382_clk;
  logic [0:0] f1382_rst;
  logic [31:0] f1382_rdata;
  sr_buffer_32_1 f1382(.wen(f1382_wen), .wdata(f1382_wdata), .clk(f1382_clk), .rst(f1382_rst), .rdata(f1382_rdata));
  assign f1382_clk = clk;
  assign f1382_rst = rst;
  // Bindings to f1382

  // f1384
  logic [0:0] f1384_wen;
  logic [31:0] f1384_wdata;
  logic [0:0] f1384_clk;
  logic [0:0] f1384_rst;
  logic [31:0] f1384_rdata;
  sr_buffer_32_1 f1384(.wen(f1384_wen), .wdata(f1384_wdata), .clk(f1384_clk), .rst(f1384_rst), .rdata(f1384_rdata));
  assign f1384_clk = clk;
  assign f1384_rst = rst;
  // Bindings to f1384

  // f1386
  logic [0:0] f1386_wen;
  logic [31:0] f1386_wdata;
  logic [0:0] f1386_clk;
  logic [0:0] f1386_rst;
  logic [31:0] f1386_rdata;
  sr_buffer_32_1 f1386(.wen(f1386_wen), .wdata(f1386_wdata), .clk(f1386_clk), .rst(f1386_rst), .rdata(f1386_rdata));
  assign f1386_clk = clk;
  assign f1386_rst = rst;
  // Bindings to f1386

  // f1388
  logic [0:0] f1388_wen;
  logic [31:0] f1388_wdata;
  logic [0:0] f1388_clk;
  logic [0:0] f1388_rst;
  logic [31:0] f1388_rdata;
  sr_buffer_32_1 f1388(.wen(f1388_wen), .wdata(f1388_wdata), .clk(f1388_clk), .rst(f1388_rst), .rdata(f1388_rdata));
  assign f1388_clk = clk;
  assign f1388_rst = rst;
  // Bindings to f1388

  // f1390
  logic [0:0] f1390_wen;
  logic [31:0] f1390_wdata;
  logic [0:0] f1390_clk;
  logic [0:0] f1390_rst;
  logic [31:0] f1390_rdata;
  sr_buffer_32_1 f1390(.wen(f1390_wen), .wdata(f1390_wdata), .clk(f1390_clk), .rst(f1390_rst), .rdata(f1390_rdata));
  assign f1390_clk = clk;
  assign f1390_rst = rst;
  // Bindings to f1390

  // f1392
  logic [0:0] f1392_wen;
  logic [31:0] f1392_wdata;
  logic [0:0] f1392_clk;
  logic [0:0] f1392_rst;
  logic [31:0] f1392_rdata;
  sr_buffer_32_1 f1392(.wen(f1392_wen), .wdata(f1392_wdata), .clk(f1392_clk), .rst(f1392_rst), .rdata(f1392_rdata));
  assign f1392_clk = clk;
  assign f1392_rst = rst;
  // Bindings to f1392

  // f1394
  logic [0:0] f1394_wen;
  logic [31:0] f1394_wdata;
  logic [0:0] f1394_clk;
  logic [0:0] f1394_rst;
  logic [31:0] f1394_rdata;
  sr_buffer_32_1 f1394(.wen(f1394_wen), .wdata(f1394_wdata), .clk(f1394_clk), .rst(f1394_rst), .rdata(f1394_rdata));
  assign f1394_clk = clk;
  assign f1394_rst = rst;
  // Bindings to f1394

  // f1396
  logic [0:0] f1396_wen;
  logic [31:0] f1396_wdata;
  logic [0:0] f1396_clk;
  logic [0:0] f1396_rst;
  logic [31:0] f1396_rdata;
  sr_buffer_32_1 f1396(.wen(f1396_wen), .wdata(f1396_wdata), .clk(f1396_clk), .rst(f1396_rst), .rdata(f1396_rdata));
  assign f1396_clk = clk;
  assign f1396_rst = rst;
  // Bindings to f1396

  // f1398
  logic [0:0] f1398_wen;
  logic [31:0] f1398_wdata;
  logic [0:0] f1398_clk;
  logic [0:0] f1398_rst;
  logic [31:0] f1398_rdata;
  sr_buffer_32_1 f1398(.wen(f1398_wen), .wdata(f1398_wdata), .clk(f1398_clk), .rst(f1398_rst), .rdata(f1398_rdata));
  assign f1398_clk = clk;
  assign f1398_rst = rst;
  // Bindings to f1398

  // f1400
  logic [0:0] f1400_wen;
  logic [31:0] f1400_wdata;
  logic [0:0] f1400_clk;
  logic [0:0] f1400_rst;
  logic [31:0] f1400_rdata;
  sr_buffer_32_1 f1400(.wen(f1400_wen), .wdata(f1400_wdata), .clk(f1400_clk), .rst(f1400_rst), .rdata(f1400_rdata));
  assign f1400_clk = clk;
  assign f1400_rst = rst;
  // Bindings to f1400

  // f1402
  logic [0:0] f1402_wen;
  logic [31:0] f1402_wdata;
  logic [0:0] f1402_clk;
  logic [0:0] f1402_rst;
  logic [31:0] f1402_rdata;
  sr_buffer_32_1 f1402(.wen(f1402_wen), .wdata(f1402_wdata), .clk(f1402_clk), .rst(f1402_rst), .rdata(f1402_rdata));
  assign f1402_clk = clk;
  assign f1402_rst = rst;
  // Bindings to f1402

  // f1404
  logic [0:0] f1404_wen;
  logic [31:0] f1404_wdata;
  logic [0:0] f1404_clk;
  logic [0:0] f1404_rst;
  logic [31:0] f1404_rdata;
  sr_buffer_32_1 f1404(.wen(f1404_wen), .wdata(f1404_wdata), .clk(f1404_clk), .rst(f1404_rst), .rdata(f1404_rdata));
  assign f1404_clk = clk;
  assign f1404_rst = rst;
  // Bindings to f1404

  // f1406
  logic [0:0] f1406_wen;
  logic [31:0] f1406_wdata;
  logic [0:0] f1406_clk;
  logic [0:0] f1406_rst;
  logic [31:0] f1406_rdata;
  sr_buffer_32_1 f1406(.wen(f1406_wen), .wdata(f1406_wdata), .clk(f1406_clk), .rst(f1406_rst), .rdata(f1406_rdata));
  assign f1406_clk = clk;
  assign f1406_rst = rst;
  // Bindings to f1406

  // f1408
  logic [0:0] f1408_wen;
  logic [31:0] f1408_wdata;
  logic [0:0] f1408_clk;
  logic [0:0] f1408_rst;
  logic [31:0] f1408_rdata;
  sr_buffer_32_1 f1408(.wen(f1408_wen), .wdata(f1408_wdata), .clk(f1408_clk), .rst(f1408_rst), .rdata(f1408_rdata));
  assign f1408_clk = clk;
  assign f1408_rst = rst;
  // Bindings to f1408

  // f1410
  logic [0:0] f1410_wen;
  logic [31:0] f1410_wdata;
  logic [0:0] f1410_clk;
  logic [0:0] f1410_rst;
  logic [31:0] f1410_rdata;
  sr_buffer_32_1 f1410(.wen(f1410_wen), .wdata(f1410_wdata), .clk(f1410_clk), .rst(f1410_rst), .rdata(f1410_rdata));
  assign f1410_clk = clk;
  assign f1410_rst = rst;
  // Bindings to f1410

  // f1412
  logic [0:0] f1412_wen;
  logic [31:0] f1412_wdata;
  logic [0:0] f1412_clk;
  logic [0:0] f1412_rst;
  logic [31:0] f1412_rdata;
  sr_buffer_32_1 f1412(.wen(f1412_wen), .wdata(f1412_wdata), .clk(f1412_clk), .rst(f1412_rst), .rdata(f1412_rdata));
  assign f1412_clk = clk;
  assign f1412_rst = rst;
  // Bindings to f1412

  // f1414
  logic [0:0] f1414_wen;
  logic [31:0] f1414_wdata;
  logic [0:0] f1414_clk;
  logic [0:0] f1414_rst;
  logic [31:0] f1414_rdata;
  sr_buffer_32_1 f1414(.wen(f1414_wen), .wdata(f1414_wdata), .clk(f1414_clk), .rst(f1414_rst), .rdata(f1414_rdata));
  assign f1414_clk = clk;
  assign f1414_rst = rst;
  // Bindings to f1414

  // f1416
  logic [0:0] f1416_wen;
  logic [31:0] f1416_wdata;
  logic [0:0] f1416_clk;
  logic [0:0] f1416_rst;
  logic [31:0] f1416_rdata;
  sr_buffer_32_1 f1416(.wen(f1416_wen), .wdata(f1416_wdata), .clk(f1416_clk), .rst(f1416_rst), .rdata(f1416_rdata));
  assign f1416_clk = clk;
  assign f1416_rst = rst;
  // Bindings to f1416

  // f1418
  logic [0:0] f1418_wen;
  logic [31:0] f1418_wdata;
  logic [0:0] f1418_clk;
  logic [0:0] f1418_rst;
  logic [31:0] f1418_rdata;
  sr_buffer_32_1 f1418(.wen(f1418_wen), .wdata(f1418_wdata), .clk(f1418_clk), .rst(f1418_rst), .rdata(f1418_rdata));
  assign f1418_clk = clk;
  assign f1418_rst = rst;
  // Bindings to f1418

  // f1420
  logic [0:0] f1420_wen;
  logic [31:0] f1420_wdata;
  logic [0:0] f1420_clk;
  logic [0:0] f1420_rst;
  logic [31:0] f1420_rdata;
  sr_buffer_32_1 f1420(.wen(f1420_wen), .wdata(f1420_wdata), .clk(f1420_clk), .rst(f1420_rst), .rdata(f1420_rdata));
  assign f1420_clk = clk;
  assign f1420_rst = rst;
  // Bindings to f1420

  // f1422
  logic [0:0] f1422_wen;
  logic [31:0] f1422_wdata;
  logic [0:0] f1422_clk;
  logic [0:0] f1422_rst;
  logic [31:0] f1422_rdata;
  sr_buffer_32_1 f1422(.wen(f1422_wen), .wdata(f1422_wdata), .clk(f1422_clk), .rst(f1422_rst), .rdata(f1422_rdata));
  assign f1422_clk = clk;
  assign f1422_rst = rst;
  // Bindings to f1422

  // f1424
  logic [0:0] f1424_wen;
  logic [31:0] f1424_wdata;
  logic [0:0] f1424_clk;
  logic [0:0] f1424_rst;
  logic [31:0] f1424_rdata;
  sr_buffer_32_1 f1424(.wen(f1424_wen), .wdata(f1424_wdata), .clk(f1424_clk), .rst(f1424_rst), .rdata(f1424_rdata));
  assign f1424_clk = clk;
  assign f1424_rst = rst;
  // Bindings to f1424

  // f1426
  logic [0:0] f1426_wen;
  logic [31:0] f1426_wdata;
  logic [0:0] f1426_clk;
  logic [0:0] f1426_rst;
  logic [31:0] f1426_rdata;
  sr_buffer_32_1 f1426(.wen(f1426_wen), .wdata(f1426_wdata), .clk(f1426_clk), .rst(f1426_rst), .rdata(f1426_rdata));
  assign f1426_clk = clk;
  assign f1426_rst = rst;
  // Bindings to f1426

  // f1428
  logic [0:0] f1428_wen;
  logic [31:0] f1428_wdata;
  logic [0:0] f1428_clk;
  logic [0:0] f1428_rst;
  logic [31:0] f1428_rdata;
  sr_buffer_32_1 f1428(.wen(f1428_wen), .wdata(f1428_wdata), .clk(f1428_clk), .rst(f1428_rst), .rdata(f1428_rdata));
  assign f1428_clk = clk;
  assign f1428_rst = rst;
  // Bindings to f1428

  // f1430
  logic [0:0] f1430_wen;
  logic [31:0] f1430_wdata;
  logic [0:0] f1430_clk;
  logic [0:0] f1430_rst;
  logic [31:0] f1430_rdata;
  sr_buffer_32_1 f1430(.wen(f1430_wen), .wdata(f1430_wdata), .clk(f1430_clk), .rst(f1430_rst), .rdata(f1430_rdata));
  assign f1430_clk = clk;
  assign f1430_rst = rst;
  // Bindings to f1430

  // f1432
  logic [0:0] f1432_wen;
  logic [31:0] f1432_wdata;
  logic [0:0] f1432_clk;
  logic [0:0] f1432_rst;
  logic [31:0] f1432_rdata;
  sr_buffer_32_1 f1432(.wen(f1432_wen), .wdata(f1432_wdata), .clk(f1432_clk), .rst(f1432_rst), .rdata(f1432_rdata));
  assign f1432_clk = clk;
  assign f1432_rst = rst;
  // Bindings to f1432

  // f1434
  logic [0:0] f1434_wen;
  logic [31:0] f1434_wdata;
  logic [0:0] f1434_clk;
  logic [0:0] f1434_rst;
  logic [31:0] f1434_rdata;
  sr_buffer_32_1 f1434(.wen(f1434_wen), .wdata(f1434_wdata), .clk(f1434_clk), .rst(f1434_rst), .rdata(f1434_rdata));
  assign f1434_clk = clk;
  assign f1434_rst = rst;
  // Bindings to f1434

  // f1436
  logic [0:0] f1436_wen;
  logic [31:0] f1436_wdata;
  logic [0:0] f1436_clk;
  logic [0:0] f1436_rst;
  logic [31:0] f1436_rdata;
  sr_buffer_32_1 f1436(.wen(f1436_wen), .wdata(f1436_wdata), .clk(f1436_clk), .rst(f1436_rst), .rdata(f1436_rdata));
  assign f1436_clk = clk;
  assign f1436_rst = rst;
  // Bindings to f1436

  // f1438
  logic [0:0] f1438_wen;
  logic [31:0] f1438_wdata;
  logic [0:0] f1438_clk;
  logic [0:0] f1438_rst;
  logic [31:0] f1438_rdata;
  sr_buffer_32_1 f1438(.wen(f1438_wen), .wdata(f1438_wdata), .clk(f1438_clk), .rst(f1438_rst), .rdata(f1438_rdata));
  assign f1438_clk = clk;
  assign f1438_rst = rst;
  // Bindings to f1438

  // f1440
  logic [0:0] f1440_wen;
  logic [31:0] f1440_wdata;
  logic [0:0] f1440_clk;
  logic [0:0] f1440_rst;
  logic [31:0] f1440_rdata;
  sr_buffer_32_1 f1440(.wen(f1440_wen), .wdata(f1440_wdata), .clk(f1440_clk), .rst(f1440_rst), .rdata(f1440_rdata));
  assign f1440_clk = clk;
  assign f1440_rst = rst;
  // Bindings to f1440

  // f1442
  logic [0:0] f1442_wen;
  logic [31:0] f1442_wdata;
  logic [0:0] f1442_clk;
  logic [0:0] f1442_rst;
  logic [31:0] f1442_rdata;
  sr_buffer_32_1 f1442(.wen(f1442_wen), .wdata(f1442_wdata), .clk(f1442_clk), .rst(f1442_rst), .rdata(f1442_rdata));
  assign f1442_clk = clk;
  assign f1442_rst = rst;
  // Bindings to f1442

  // f1444
  logic [0:0] f1444_wen;
  logic [31:0] f1444_wdata;
  logic [0:0] f1444_clk;
  logic [0:0] f1444_rst;
  logic [31:0] f1444_rdata;
  sr_buffer_32_1 f1444(.wen(f1444_wen), .wdata(f1444_wdata), .clk(f1444_clk), .rst(f1444_rst), .rdata(f1444_rdata));
  assign f1444_clk = clk;
  assign f1444_rst = rst;
  // Bindings to f1444

  // f1446
  logic [0:0] f1446_wen;
  logic [31:0] f1446_wdata;
  logic [0:0] f1446_clk;
  logic [0:0] f1446_rst;
  logic [31:0] f1446_rdata;
  sr_buffer_32_1 f1446(.wen(f1446_wen), .wdata(f1446_wdata), .clk(f1446_clk), .rst(f1446_rst), .rdata(f1446_rdata));
  assign f1446_clk = clk;
  assign f1446_rst = rst;
  // Bindings to f1446

  // f1448
  logic [0:0] f1448_wen;
  logic [31:0] f1448_wdata;
  logic [0:0] f1448_clk;
  logic [0:0] f1448_rst;
  logic [31:0] f1448_rdata;
  sr_buffer_32_1 f1448(.wen(f1448_wen), .wdata(f1448_wdata), .clk(f1448_clk), .rst(f1448_rst), .rdata(f1448_rdata));
  assign f1448_clk = clk;
  assign f1448_rst = rst;
  // Bindings to f1448

  // f1450
  logic [0:0] f1450_wen;
  logic [31:0] f1450_wdata;
  logic [0:0] f1450_clk;
  logic [0:0] f1450_rst;
  logic [31:0] f1450_rdata;
  sr_buffer_32_1 f1450(.wen(f1450_wen), .wdata(f1450_wdata), .clk(f1450_clk), .rst(f1450_rst), .rdata(f1450_rdata));
  assign f1450_clk = clk;
  assign f1450_rst = rst;
  // Bindings to f1450

  // f1452
  logic [0:0] f1452_wen;
  logic [31:0] f1452_wdata;
  logic [0:0] f1452_clk;
  logic [0:0] f1452_rst;
  logic [31:0] f1452_rdata;
  sr_buffer_32_1 f1452(.wen(f1452_wen), .wdata(f1452_wdata), .clk(f1452_clk), .rst(f1452_rst), .rdata(f1452_rdata));
  assign f1452_clk = clk;
  assign f1452_rst = rst;
  // Bindings to f1452

  // f1454
  logic [0:0] f1454_wen;
  logic [31:0] f1454_wdata;
  logic [0:0] f1454_clk;
  logic [0:0] f1454_rst;
  logic [31:0] f1454_rdata;
  sr_buffer_32_1 f1454(.wen(f1454_wen), .wdata(f1454_wdata), .clk(f1454_clk), .rst(f1454_rst), .rdata(f1454_rdata));
  assign f1454_clk = clk;
  assign f1454_rst = rst;
  // Bindings to f1454

  // f1456
  logic [0:0] f1456_wen;
  logic [31:0] f1456_wdata;
  logic [0:0] f1456_clk;
  logic [0:0] f1456_rst;
  logic [31:0] f1456_rdata;
  sr_buffer_32_1 f1456(.wen(f1456_wen), .wdata(f1456_wdata), .clk(f1456_clk), .rst(f1456_rst), .rdata(f1456_rdata));
  assign f1456_clk = clk;
  assign f1456_rst = rst;
  // Bindings to f1456

  // f1458
  logic [0:0] f1458_wen;
  logic [31:0] f1458_wdata;
  logic [0:0] f1458_clk;
  logic [0:0] f1458_rst;
  logic [31:0] f1458_rdata;
  sr_buffer_32_1 f1458(.wen(f1458_wen), .wdata(f1458_wdata), .clk(f1458_clk), .rst(f1458_rst), .rdata(f1458_rdata));
  assign f1458_clk = clk;
  assign f1458_rst = rst;
  // Bindings to f1458

  // f1460
  logic [0:0] f1460_wen;
  logic [31:0] f1460_wdata;
  logic [0:0] f1460_clk;
  logic [0:0] f1460_rst;
  logic [31:0] f1460_rdata;
  sr_buffer_32_1 f1460(.wen(f1460_wen), .wdata(f1460_wdata), .clk(f1460_clk), .rst(f1460_rst), .rdata(f1460_rdata));
  assign f1460_clk = clk;
  assign f1460_rst = rst;
  // Bindings to f1460

  // f1462
  logic [0:0] f1462_wen;
  logic [31:0] f1462_wdata;
  logic [0:0] f1462_clk;
  logic [0:0] f1462_rst;
  logic [31:0] f1462_rdata;
  sr_buffer_32_1 f1462(.wen(f1462_wen), .wdata(f1462_wdata), .clk(f1462_clk), .rst(f1462_rst), .rdata(f1462_rdata));
  assign f1462_clk = clk;
  assign f1462_rst = rst;
  // Bindings to f1462

  // f1464
  logic [0:0] f1464_wen;
  logic [31:0] f1464_wdata;
  logic [0:0] f1464_clk;
  logic [0:0] f1464_rst;
  logic [31:0] f1464_rdata;
  sr_buffer_32_1 f1464(.wen(f1464_wen), .wdata(f1464_wdata), .clk(f1464_clk), .rst(f1464_rst), .rdata(f1464_rdata));
  assign f1464_clk = clk;
  assign f1464_rst = rst;
  // Bindings to f1464

  // f1466
  logic [0:0] f1466_wen;
  logic [31:0] f1466_wdata;
  logic [0:0] f1466_clk;
  logic [0:0] f1466_rst;
  logic [31:0] f1466_rdata;
  sr_buffer_32_1 f1466(.wen(f1466_wen), .wdata(f1466_wdata), .clk(f1466_clk), .rst(f1466_rst), .rdata(f1466_rdata));
  assign f1466_clk = clk;
  assign f1466_rst = rst;
  // Bindings to f1466

  // f1468
  logic [0:0] f1468_wen;
  logic [31:0] f1468_wdata;
  logic [0:0] f1468_clk;
  logic [0:0] f1468_rst;
  logic [31:0] f1468_rdata;
  sr_buffer_32_1 f1468(.wen(f1468_wen), .wdata(f1468_wdata), .clk(f1468_clk), .rst(f1468_rst), .rdata(f1468_rdata));
  assign f1468_clk = clk;
  assign f1468_rst = rst;
  // Bindings to f1468

  // f1470
  logic [0:0] f1470_wen;
  logic [31:0] f1470_wdata;
  logic [0:0] f1470_clk;
  logic [0:0] f1470_rst;
  logic [31:0] f1470_rdata;
  sr_buffer_32_1 f1470(.wen(f1470_wen), .wdata(f1470_wdata), .clk(f1470_clk), .rst(f1470_rst), .rdata(f1470_rdata));
  assign f1470_clk = clk;
  assign f1470_rst = rst;
  // Bindings to f1470

  // f1472
  logic [0:0] f1472_wen;
  logic [31:0] f1472_wdata;
  logic [0:0] f1472_clk;
  logic [0:0] f1472_rst;
  logic [31:0] f1472_rdata;
  sr_buffer_32_1 f1472(.wen(f1472_wen), .wdata(f1472_wdata), .clk(f1472_clk), .rst(f1472_rst), .rdata(f1472_rdata));
  assign f1472_clk = clk;
  assign f1472_rst = rst;
  // Bindings to f1472

  // f1474
  logic [0:0] f1474_wen;
  logic [31:0] f1474_wdata;
  logic [0:0] f1474_clk;
  logic [0:0] f1474_rst;
  logic [31:0] f1474_rdata;
  sr_buffer_32_1 f1474(.wen(f1474_wen), .wdata(f1474_wdata), .clk(f1474_clk), .rst(f1474_rst), .rdata(f1474_rdata));
  assign f1474_clk = clk;
  assign f1474_rst = rst;
  // Bindings to f1474

  // f1476
  logic [0:0] f1476_wen;
  logic [31:0] f1476_wdata;
  logic [0:0] f1476_clk;
  logic [0:0] f1476_rst;
  logic [31:0] f1476_rdata;
  sr_buffer_32_1 f1476(.wen(f1476_wen), .wdata(f1476_wdata), .clk(f1476_clk), .rst(f1476_rst), .rdata(f1476_rdata));
  assign f1476_clk = clk;
  assign f1476_rst = rst;
  // Bindings to f1476

  // f1478
  logic [0:0] f1478_wen;
  logic [31:0] f1478_wdata;
  logic [0:0] f1478_clk;
  logic [0:0] f1478_rst;
  logic [31:0] f1478_rdata;
  sr_buffer_32_1 f1478(.wen(f1478_wen), .wdata(f1478_wdata), .clk(f1478_clk), .rst(f1478_rst), .rdata(f1478_rdata));
  assign f1478_clk = clk;
  assign f1478_rst = rst;
  // Bindings to f1478

  // f1480
  logic [0:0] f1480_wen;
  logic [31:0] f1480_wdata;
  logic [0:0] f1480_clk;
  logic [0:0] f1480_rst;
  logic [31:0] f1480_rdata;
  sr_buffer_32_1 f1480(.wen(f1480_wen), .wdata(f1480_wdata), .clk(f1480_clk), .rst(f1480_rst), .rdata(f1480_rdata));
  assign f1480_clk = clk;
  assign f1480_rst = rst;
  // Bindings to f1480

  // f1482
  logic [0:0] f1482_wen;
  logic [31:0] f1482_wdata;
  logic [0:0] f1482_clk;
  logic [0:0] f1482_rst;
  logic [31:0] f1482_rdata;
  sr_buffer_32_1 f1482(.wen(f1482_wen), .wdata(f1482_wdata), .clk(f1482_clk), .rst(f1482_rst), .rdata(f1482_rdata));
  assign f1482_clk = clk;
  assign f1482_rst = rst;
  // Bindings to f1482

  // f1484
  logic [0:0] f1484_wen;
  logic [31:0] f1484_wdata;
  logic [0:0] f1484_clk;
  logic [0:0] f1484_rst;
  logic [31:0] f1484_rdata;
  sr_buffer_32_1 f1484(.wen(f1484_wen), .wdata(f1484_wdata), .clk(f1484_clk), .rst(f1484_rst), .rdata(f1484_rdata));
  assign f1484_clk = clk;
  assign f1484_rst = rst;
  // Bindings to f1484

  // f1486
  logic [0:0] f1486_wen;
  logic [31:0] f1486_wdata;
  logic [0:0] f1486_clk;
  logic [0:0] f1486_rst;
  logic [31:0] f1486_rdata;
  sr_buffer_32_1 f1486(.wen(f1486_wen), .wdata(f1486_wdata), .clk(f1486_clk), .rst(f1486_rst), .rdata(f1486_rdata));
  assign f1486_clk = clk;
  assign f1486_rst = rst;
  // Bindings to f1486

  // f1488
  logic [0:0] f1488_wen;
  logic [31:0] f1488_wdata;
  logic [0:0] f1488_clk;
  logic [0:0] f1488_rst;
  logic [31:0] f1488_rdata;
  sr_buffer_32_1 f1488(.wen(f1488_wen), .wdata(f1488_wdata), .clk(f1488_clk), .rst(f1488_rst), .rdata(f1488_rdata));
  assign f1488_clk = clk;
  assign f1488_rst = rst;
  // Bindings to f1488

  // f1490
  logic [0:0] f1490_wen;
  logic [31:0] f1490_wdata;
  logic [0:0] f1490_clk;
  logic [0:0] f1490_rst;
  logic [31:0] f1490_rdata;
  sr_buffer_32_1 f1490(.wen(f1490_wen), .wdata(f1490_wdata), .clk(f1490_clk), .rst(f1490_rst), .rdata(f1490_rdata));
  assign f1490_clk = clk;
  assign f1490_rst = rst;
  // Bindings to f1490

  // f1492
  logic [0:0] f1492_wen;
  logic [31:0] f1492_wdata;
  logic [0:0] f1492_clk;
  logic [0:0] f1492_rst;
  logic [31:0] f1492_rdata;
  sr_buffer_32_1 f1492(.wen(f1492_wen), .wdata(f1492_wdata), .clk(f1492_clk), .rst(f1492_rst), .rdata(f1492_rdata));
  assign f1492_clk = clk;
  assign f1492_rst = rst;
  // Bindings to f1492

  // f1494
  logic [0:0] f1494_wen;
  logic [31:0] f1494_wdata;
  logic [0:0] f1494_clk;
  logic [0:0] f1494_rst;
  logic [31:0] f1494_rdata;
  sr_buffer_32_1 f1494(.wen(f1494_wen), .wdata(f1494_wdata), .clk(f1494_clk), .rst(f1494_rst), .rdata(f1494_rdata));
  assign f1494_clk = clk;
  assign f1494_rst = rst;
  // Bindings to f1494

  // f1496
  logic [0:0] f1496_wen;
  logic [31:0] f1496_wdata;
  logic [0:0] f1496_clk;
  logic [0:0] f1496_rst;
  logic [31:0] f1496_rdata;
  sr_buffer_32_1 f1496(.wen(f1496_wen), .wdata(f1496_wdata), .clk(f1496_clk), .rst(f1496_rst), .rdata(f1496_rdata));
  assign f1496_clk = clk;
  assign f1496_rst = rst;
  // Bindings to f1496

  // f1498
  logic [0:0] f1498_wen;
  logic [31:0] f1498_wdata;
  logic [0:0] f1498_clk;
  logic [0:0] f1498_rst;
  logic [31:0] f1498_rdata;
  sr_buffer_32_1 f1498(.wen(f1498_wen), .wdata(f1498_wdata), .clk(f1498_clk), .rst(f1498_rst), .rdata(f1498_rdata));
  assign f1498_clk = clk;
  assign f1498_rst = rst;
  // Bindings to f1498

  // f1500
  logic [0:0] f1500_wen;
  logic [31:0] f1500_wdata;
  logic [0:0] f1500_clk;
  logic [0:0] f1500_rst;
  logic [31:0] f1500_rdata;
  sr_buffer_32_1 f1500(.wen(f1500_wen), .wdata(f1500_wdata), .clk(f1500_clk), .rst(f1500_rst), .rdata(f1500_rdata));
  assign f1500_clk = clk;
  assign f1500_rst = rst;
  // Bindings to f1500

  // f1502
  logic [0:0] f1502_wen;
  logic [31:0] f1502_wdata;
  logic [0:0] f1502_clk;
  logic [0:0] f1502_rst;
  logic [31:0] f1502_rdata;
  sr_buffer_32_1 f1502(.wen(f1502_wen), .wdata(f1502_wdata), .clk(f1502_clk), .rst(f1502_rst), .rdata(f1502_rdata));
  assign f1502_clk = clk;
  assign f1502_rst = rst;
  // Bindings to f1502

  // f1504
  logic [0:0] f1504_wen;
  logic [31:0] f1504_wdata;
  logic [0:0] f1504_clk;
  logic [0:0] f1504_rst;
  logic [31:0] f1504_rdata;
  sr_buffer_32_1 f1504(.wen(f1504_wen), .wdata(f1504_wdata), .clk(f1504_clk), .rst(f1504_rst), .rdata(f1504_rdata));
  assign f1504_clk = clk;
  assign f1504_rst = rst;
  // Bindings to f1504

  // f1506
  logic [0:0] f1506_wen;
  logic [31:0] f1506_wdata;
  logic [0:0] f1506_clk;
  logic [0:0] f1506_rst;
  logic [31:0] f1506_rdata;
  sr_buffer_32_1 f1506(.wen(f1506_wen), .wdata(f1506_wdata), .clk(f1506_clk), .rst(f1506_rst), .rdata(f1506_rdata));
  assign f1506_clk = clk;
  assign f1506_rst = rst;
  // Bindings to f1506

  // f1508
  logic [0:0] f1508_wen;
  logic [31:0] f1508_wdata;
  logic [0:0] f1508_clk;
  logic [0:0] f1508_rst;
  logic [31:0] f1508_rdata;
  sr_buffer_32_1 f1508(.wen(f1508_wen), .wdata(f1508_wdata), .clk(f1508_clk), .rst(f1508_rst), .rdata(f1508_rdata));
  assign f1508_clk = clk;
  assign f1508_rst = rst;
  // Bindings to f1508

  // f1510
  logic [0:0] f1510_wen;
  logic [31:0] f1510_wdata;
  logic [0:0] f1510_clk;
  logic [0:0] f1510_rst;
  logic [31:0] f1510_rdata;
  sr_buffer_32_1 f1510(.wen(f1510_wen), .wdata(f1510_wdata), .clk(f1510_clk), .rst(f1510_rst), .rdata(f1510_rdata));
  assign f1510_clk = clk;
  assign f1510_rst = rst;
  // Bindings to f1510

  // f1512
  logic [0:0] f1512_wen;
  logic [31:0] f1512_wdata;
  logic [0:0] f1512_clk;
  logic [0:0] f1512_rst;
  logic [31:0] f1512_rdata;
  sr_buffer_32_1 f1512(.wen(f1512_wen), .wdata(f1512_wdata), .clk(f1512_clk), .rst(f1512_rst), .rdata(f1512_rdata));
  assign f1512_clk = clk;
  assign f1512_rst = rst;
  // Bindings to f1512

  // f1514
  logic [0:0] f1514_wen;
  logic [31:0] f1514_wdata;
  logic [0:0] f1514_clk;
  logic [0:0] f1514_rst;
  logic [31:0] f1514_rdata;
  sr_buffer_32_1 f1514(.wen(f1514_wen), .wdata(f1514_wdata), .clk(f1514_clk), .rst(f1514_rst), .rdata(f1514_rdata));
  assign f1514_clk = clk;
  assign f1514_rst = rst;
  // Bindings to f1514

  // f1516
  logic [0:0] f1516_wen;
  logic [31:0] f1516_wdata;
  logic [0:0] f1516_clk;
  logic [0:0] f1516_rst;
  logic [31:0] f1516_rdata;
  sr_buffer_32_1 f1516(.wen(f1516_wen), .wdata(f1516_wdata), .clk(f1516_clk), .rst(f1516_rst), .rdata(f1516_rdata));
  assign f1516_clk = clk;
  assign f1516_rst = rst;
  // Bindings to f1516

  // f1518
  logic [0:0] f1518_wen;
  logic [31:0] f1518_wdata;
  logic [0:0] f1518_clk;
  logic [0:0] f1518_rst;
  logic [31:0] f1518_rdata;
  sr_buffer_32_1 f1518(.wen(f1518_wen), .wdata(f1518_wdata), .clk(f1518_clk), .rst(f1518_rst), .rdata(f1518_rdata));
  assign f1518_clk = clk;
  assign f1518_rst = rst;
  // Bindings to f1518

  // f1520
  logic [0:0] f1520_wen;
  logic [31:0] f1520_wdata;
  logic [0:0] f1520_clk;
  logic [0:0] f1520_rst;
  logic [31:0] f1520_rdata;
  sr_buffer_32_1 f1520(.wen(f1520_wen), .wdata(f1520_wdata), .clk(f1520_clk), .rst(f1520_rst), .rdata(f1520_rdata));
  assign f1520_clk = clk;
  assign f1520_rst = rst;
  // Bindings to f1520

  // f1522
  logic [0:0] f1522_wen;
  logic [31:0] f1522_wdata;
  logic [0:0] f1522_clk;
  logic [0:0] f1522_rst;
  logic [31:0] f1522_rdata;
  sr_buffer_32_1 f1522(.wen(f1522_wen), .wdata(f1522_wdata), .clk(f1522_clk), .rst(f1522_rst), .rdata(f1522_rdata));
  assign f1522_clk = clk;
  assign f1522_rst = rst;
  // Bindings to f1522

  // f1524
  logic [0:0] f1524_wen;
  logic [31:0] f1524_wdata;
  logic [0:0] f1524_clk;
  logic [0:0] f1524_rst;
  logic [31:0] f1524_rdata;
  sr_buffer_32_1 f1524(.wen(f1524_wen), .wdata(f1524_wdata), .clk(f1524_clk), .rst(f1524_rst), .rdata(f1524_rdata));
  assign f1524_clk = clk;
  assign f1524_rst = rst;
  // Bindings to f1524

  // f1526
  logic [0:0] f1526_wen;
  logic [31:0] f1526_wdata;
  logic [0:0] f1526_clk;
  logic [0:0] f1526_rst;
  logic [31:0] f1526_rdata;
  sr_buffer_32_1 f1526(.wen(f1526_wen), .wdata(f1526_wdata), .clk(f1526_clk), .rst(f1526_rst), .rdata(f1526_rdata));
  assign f1526_clk = clk;
  assign f1526_rst = rst;
  // Bindings to f1526

  // f1528
  logic [0:0] f1528_wen;
  logic [31:0] f1528_wdata;
  logic [0:0] f1528_clk;
  logic [0:0] f1528_rst;
  logic [31:0] f1528_rdata;
  sr_buffer_32_1 f1528(.wen(f1528_wen), .wdata(f1528_wdata), .clk(f1528_clk), .rst(f1528_rst), .rdata(f1528_rdata));
  assign f1528_clk = clk;
  assign f1528_rst = rst;
  // Bindings to f1528

  // f1530
  logic [0:0] f1530_wen;
  logic [31:0] f1530_wdata;
  logic [0:0] f1530_clk;
  logic [0:0] f1530_rst;
  logic [31:0] f1530_rdata;
  sr_buffer_32_1 f1530(.wen(f1530_wen), .wdata(f1530_wdata), .clk(f1530_clk), .rst(f1530_rst), .rdata(f1530_rdata));
  assign f1530_clk = clk;
  assign f1530_rst = rst;
  // Bindings to f1530

  // f1532
  logic [0:0] f1532_wen;
  logic [31:0] f1532_wdata;
  logic [0:0] f1532_clk;
  logic [0:0] f1532_rst;
  logic [31:0] f1532_rdata;
  sr_buffer_32_1 f1532(.wen(f1532_wen), .wdata(f1532_wdata), .clk(f1532_clk), .rst(f1532_rst), .rdata(f1532_rdata));
  assign f1532_clk = clk;
  assign f1532_rst = rst;
  // Bindings to f1532

  // f1534
  logic [0:0] f1534_wen;
  logic [31:0] f1534_wdata;
  logic [0:0] f1534_clk;
  logic [0:0] f1534_rst;
  logic [31:0] f1534_rdata;
  sr_buffer_32_1 f1534(.wen(f1534_wen), .wdata(f1534_wdata), .clk(f1534_clk), .rst(f1534_rst), .rdata(f1534_rdata));
  assign f1534_clk = clk;
  assign f1534_rst = rst;
  // Bindings to f1534

  // f1536
  logic [0:0] f1536_wen;
  logic [31:0] f1536_wdata;
  logic [0:0] f1536_clk;
  logic [0:0] f1536_rst;
  logic [31:0] f1536_rdata;
  sr_buffer_32_1 f1536(.wen(f1536_wen), .wdata(f1536_wdata), .clk(f1536_clk), .rst(f1536_rst), .rdata(f1536_rdata));
  assign f1536_clk = clk;
  assign f1536_rst = rst;
  // Bindings to f1536

  // f1538
  logic [0:0] f1538_wen;
  logic [31:0] f1538_wdata;
  logic [0:0] f1538_clk;
  logic [0:0] f1538_rst;
  logic [31:0] f1538_rdata;
  sr_buffer_32_1 f1538(.wen(f1538_wen), .wdata(f1538_wdata), .clk(f1538_clk), .rst(f1538_rst), .rdata(f1538_rdata));
  assign f1538_clk = clk;
  assign f1538_rst = rst;
  // Bindings to f1538

  // f1540
  logic [0:0] f1540_wen;
  logic [31:0] f1540_wdata;
  logic [0:0] f1540_clk;
  logic [0:0] f1540_rst;
  logic [31:0] f1540_rdata;
  sr_buffer_32_1 f1540(.wen(f1540_wen), .wdata(f1540_wdata), .clk(f1540_clk), .rst(f1540_rst), .rdata(f1540_rdata));
  assign f1540_clk = clk;
  assign f1540_rst = rst;
  // Bindings to f1540

  // f1542
  logic [0:0] f1542_wen;
  logic [31:0] f1542_wdata;
  logic [0:0] f1542_clk;
  logic [0:0] f1542_rst;
  logic [31:0] f1542_rdata;
  sr_buffer_32_1 f1542(.wen(f1542_wen), .wdata(f1542_wdata), .clk(f1542_clk), .rst(f1542_rst), .rdata(f1542_rdata));
  assign f1542_clk = clk;
  assign f1542_rst = rst;
  // Bindings to f1542

  // f1544
  logic [0:0] f1544_wen;
  logic [31:0] f1544_wdata;
  logic [0:0] f1544_clk;
  logic [0:0] f1544_rst;
  logic [31:0] f1544_rdata;
  sr_buffer_32_1 f1544(.wen(f1544_wen), .wdata(f1544_wdata), .clk(f1544_clk), .rst(f1544_rst), .rdata(f1544_rdata));
  assign f1544_clk = clk;
  assign f1544_rst = rst;
  // Bindings to f1544

  // f1546
  logic [0:0] f1546_wen;
  logic [31:0] f1546_wdata;
  logic [0:0] f1546_clk;
  logic [0:0] f1546_rst;
  logic [31:0] f1546_rdata;
  sr_buffer_32_1 f1546(.wen(f1546_wen), .wdata(f1546_wdata), .clk(f1546_clk), .rst(f1546_rst), .rdata(f1546_rdata));
  assign f1546_clk = clk;
  assign f1546_rst = rst;
  // Bindings to f1546

  // f1548
  logic [0:0] f1548_wen;
  logic [31:0] f1548_wdata;
  logic [0:0] f1548_clk;
  logic [0:0] f1548_rst;
  logic [31:0] f1548_rdata;
  sr_buffer_32_1 f1548(.wen(f1548_wen), .wdata(f1548_wdata), .clk(f1548_clk), .rst(f1548_rst), .rdata(f1548_rdata));
  assign f1548_clk = clk;
  assign f1548_rst = rst;
  // Bindings to f1548

  // f1550
  logic [0:0] f1550_wen;
  logic [31:0] f1550_wdata;
  logic [0:0] f1550_clk;
  logic [0:0] f1550_rst;
  logic [31:0] f1550_rdata;
  sr_buffer_32_1 f1550(.wen(f1550_wen), .wdata(f1550_wdata), .clk(f1550_clk), .rst(f1550_rst), .rdata(f1550_rdata));
  assign f1550_clk = clk;
  assign f1550_rst = rst;
  // Bindings to f1550

  // f1552
  logic [0:0] f1552_wen;
  logic [31:0] f1552_wdata;
  logic [0:0] f1552_clk;
  logic [0:0] f1552_rst;
  logic [31:0] f1552_rdata;
  sr_buffer_32_1 f1552(.wen(f1552_wen), .wdata(f1552_wdata), .clk(f1552_clk), .rst(f1552_rst), .rdata(f1552_rdata));
  assign f1552_clk = clk;
  assign f1552_rst = rst;
  // Bindings to f1552

  // f1554
  logic [0:0] f1554_wen;
  logic [31:0] f1554_wdata;
  logic [0:0] f1554_clk;
  logic [0:0] f1554_rst;
  logic [31:0] f1554_rdata;
  sr_buffer_32_1 f1554(.wen(f1554_wen), .wdata(f1554_wdata), .clk(f1554_clk), .rst(f1554_rst), .rdata(f1554_rdata));
  assign f1554_clk = clk;
  assign f1554_rst = rst;
  // Bindings to f1554

  // f1556
  logic [0:0] f1556_wen;
  logic [31:0] f1556_wdata;
  logic [0:0] f1556_clk;
  logic [0:0] f1556_rst;
  logic [31:0] f1556_rdata;
  sr_buffer_32_1 f1556(.wen(f1556_wen), .wdata(f1556_wdata), .clk(f1556_clk), .rst(f1556_rst), .rdata(f1556_rdata));
  assign f1556_clk = clk;
  assign f1556_rst = rst;
  // Bindings to f1556

  // f1558
  logic [0:0] f1558_wen;
  logic [31:0] f1558_wdata;
  logic [0:0] f1558_clk;
  logic [0:0] f1558_rst;
  logic [31:0] f1558_rdata;
  sr_buffer_32_1 f1558(.wen(f1558_wen), .wdata(f1558_wdata), .clk(f1558_clk), .rst(f1558_rst), .rdata(f1558_rdata));
  assign f1558_clk = clk;
  assign f1558_rst = rst;
  // Bindings to f1558

  // f1560
  logic [0:0] f1560_wen;
  logic [31:0] f1560_wdata;
  logic [0:0] f1560_clk;
  logic [0:0] f1560_rst;
  logic [31:0] f1560_rdata;
  sr_buffer_32_1 f1560(.wen(f1560_wen), .wdata(f1560_wdata), .clk(f1560_clk), .rst(f1560_rst), .rdata(f1560_rdata));
  assign f1560_clk = clk;
  assign f1560_rst = rst;
  // Bindings to f1560

  // f1562
  logic [0:0] f1562_wen;
  logic [31:0] f1562_wdata;
  logic [0:0] f1562_clk;
  logic [0:0] f1562_rst;
  logic [31:0] f1562_rdata;
  sr_buffer_32_1 f1562(.wen(f1562_wen), .wdata(f1562_wdata), .clk(f1562_clk), .rst(f1562_rst), .rdata(f1562_rdata));
  assign f1562_clk = clk;
  assign f1562_rst = rst;
  // Bindings to f1562

  // f1564
  logic [0:0] f1564_wen;
  logic [31:0] f1564_wdata;
  logic [0:0] f1564_clk;
  logic [0:0] f1564_rst;
  logic [31:0] f1564_rdata;
  sr_buffer_32_1 f1564(.wen(f1564_wen), .wdata(f1564_wdata), .clk(f1564_clk), .rst(f1564_rst), .rdata(f1564_rdata));
  assign f1564_clk = clk;
  assign f1564_rst = rst;
  // Bindings to f1564

  // f1566
  logic [0:0] f1566_wen;
  logic [31:0] f1566_wdata;
  logic [0:0] f1566_clk;
  logic [0:0] f1566_rst;
  logic [31:0] f1566_rdata;
  sr_buffer_32_1 f1566(.wen(f1566_wen), .wdata(f1566_wdata), .clk(f1566_clk), .rst(f1566_rst), .rdata(f1566_rdata));
  assign f1566_clk = clk;
  assign f1566_rst = rst;
  // Bindings to f1566

  // f1568
  logic [0:0] f1568_wen;
  logic [31:0] f1568_wdata;
  logic [0:0] f1568_clk;
  logic [0:0] f1568_rst;
  logic [31:0] f1568_rdata;
  sr_buffer_32_1 f1568(.wen(f1568_wen), .wdata(f1568_wdata), .clk(f1568_clk), .rst(f1568_rst), .rdata(f1568_rdata));
  assign f1568_clk = clk;
  assign f1568_rst = rst;
  // Bindings to f1568

  // f1570
  logic [0:0] f1570_wen;
  logic [31:0] f1570_wdata;
  logic [0:0] f1570_clk;
  logic [0:0] f1570_rst;
  logic [31:0] f1570_rdata;
  sr_buffer_32_1 f1570(.wen(f1570_wen), .wdata(f1570_wdata), .clk(f1570_clk), .rst(f1570_rst), .rdata(f1570_rdata));
  assign f1570_clk = clk;
  assign f1570_rst = rst;
  // Bindings to f1570

  // f1572
  logic [0:0] f1572_wen;
  logic [31:0] f1572_wdata;
  logic [0:0] f1572_clk;
  logic [0:0] f1572_rst;
  logic [31:0] f1572_rdata;
  sr_buffer_32_1 f1572(.wen(f1572_wen), .wdata(f1572_wdata), .clk(f1572_clk), .rst(f1572_rst), .rdata(f1572_rdata));
  assign f1572_clk = clk;
  assign f1572_rst = rst;
  // Bindings to f1572

  // f1574
  logic [0:0] f1574_wen;
  logic [31:0] f1574_wdata;
  logic [0:0] f1574_clk;
  logic [0:0] f1574_rst;
  logic [31:0] f1574_rdata;
  sr_buffer_32_1 f1574(.wen(f1574_wen), .wdata(f1574_wdata), .clk(f1574_clk), .rst(f1574_rst), .rdata(f1574_rdata));
  assign f1574_clk = clk;
  assign f1574_rst = rst;
  // Bindings to f1574

  // f1576
  logic [0:0] f1576_wen;
  logic [31:0] f1576_wdata;
  logic [0:0] f1576_clk;
  logic [0:0] f1576_rst;
  logic [31:0] f1576_rdata;
  sr_buffer_32_1 f1576(.wen(f1576_wen), .wdata(f1576_wdata), .clk(f1576_clk), .rst(f1576_rst), .rdata(f1576_rdata));
  assign f1576_clk = clk;
  assign f1576_rst = rst;
  // Bindings to f1576

  // f1578
  logic [0:0] f1578_wen;
  logic [31:0] f1578_wdata;
  logic [0:0] f1578_clk;
  logic [0:0] f1578_rst;
  logic [31:0] f1578_rdata;
  sr_buffer_32_1 f1578(.wen(f1578_wen), .wdata(f1578_wdata), .clk(f1578_clk), .rst(f1578_rst), .rdata(f1578_rdata));
  assign f1578_clk = clk;
  assign f1578_rst = rst;
  // Bindings to f1578

  // f1580
  logic [0:0] f1580_wen;
  logic [31:0] f1580_wdata;
  logic [0:0] f1580_clk;
  logic [0:0] f1580_rst;
  logic [31:0] f1580_rdata;
  sr_buffer_32_1 f1580(.wen(f1580_wen), .wdata(f1580_wdata), .clk(f1580_clk), .rst(f1580_rst), .rdata(f1580_rdata));
  assign f1580_clk = clk;
  assign f1580_rst = rst;
  // Bindings to f1580

  // f1582
  logic [0:0] f1582_wen;
  logic [31:0] f1582_wdata;
  logic [0:0] f1582_clk;
  logic [0:0] f1582_rst;
  logic [31:0] f1582_rdata;
  sr_buffer_32_1 f1582(.wen(f1582_wen), .wdata(f1582_wdata), .clk(f1582_clk), .rst(f1582_rst), .rdata(f1582_rdata));
  assign f1582_clk = clk;
  assign f1582_rst = rst;
  // Bindings to f1582

  // f1584
  logic [0:0] f1584_wen;
  logic [31:0] f1584_wdata;
  logic [0:0] f1584_clk;
  logic [0:0] f1584_rst;
  logic [31:0] f1584_rdata;
  sr_buffer_32_1 f1584(.wen(f1584_wen), .wdata(f1584_wdata), .clk(f1584_clk), .rst(f1584_rst), .rdata(f1584_rdata));
  assign f1584_clk = clk;
  assign f1584_rst = rst;
  // Bindings to f1584

  // f1586
  logic [0:0] f1586_wen;
  logic [31:0] f1586_wdata;
  logic [0:0] f1586_clk;
  logic [0:0] f1586_rst;
  logic [31:0] f1586_rdata;
  sr_buffer_32_1 f1586(.wen(f1586_wen), .wdata(f1586_wdata), .clk(f1586_clk), .rst(f1586_rst), .rdata(f1586_rdata));
  assign f1586_clk = clk;
  assign f1586_rst = rst;
  // Bindings to f1586

  // f1588
  logic [0:0] f1588_wen;
  logic [31:0] f1588_wdata;
  logic [0:0] f1588_clk;
  logic [0:0] f1588_rst;
  logic [31:0] f1588_rdata;
  sr_buffer_32_1 f1588(.wen(f1588_wen), .wdata(f1588_wdata), .clk(f1588_clk), .rst(f1588_rst), .rdata(f1588_rdata));
  assign f1588_clk = clk;
  assign f1588_rst = rst;
  // Bindings to f1588

  // f1590
  logic [0:0] f1590_wen;
  logic [31:0] f1590_wdata;
  logic [0:0] f1590_clk;
  logic [0:0] f1590_rst;
  logic [31:0] f1590_rdata;
  sr_buffer_32_1 f1590(.wen(f1590_wen), .wdata(f1590_wdata), .clk(f1590_clk), .rst(f1590_rst), .rdata(f1590_rdata));
  assign f1590_clk = clk;
  assign f1590_rst = rst;
  // Bindings to f1590

  // f1592
  logic [0:0] f1592_wen;
  logic [31:0] f1592_wdata;
  logic [0:0] f1592_clk;
  logic [0:0] f1592_rst;
  logic [31:0] f1592_rdata;
  sr_buffer_32_1 f1592(.wen(f1592_wen), .wdata(f1592_wdata), .clk(f1592_clk), .rst(f1592_rst), .rdata(f1592_rdata));
  assign f1592_clk = clk;
  assign f1592_rst = rst;
  // Bindings to f1592

  // f1594
  logic [0:0] f1594_wen;
  logic [31:0] f1594_wdata;
  logic [0:0] f1594_clk;
  logic [0:0] f1594_rst;
  logic [31:0] f1594_rdata;
  sr_buffer_32_1 f1594(.wen(f1594_wen), .wdata(f1594_wdata), .clk(f1594_clk), .rst(f1594_rst), .rdata(f1594_rdata));
  assign f1594_clk = clk;
  assign f1594_rst = rst;
  // Bindings to f1594

  // f1596
  logic [0:0] f1596_wen;
  logic [31:0] f1596_wdata;
  logic [0:0] f1596_clk;
  logic [0:0] f1596_rst;
  logic [31:0] f1596_rdata;
  sr_buffer_32_1 f1596(.wen(f1596_wen), .wdata(f1596_wdata), .clk(f1596_clk), .rst(f1596_rst), .rdata(f1596_rdata));
  assign f1596_clk = clk;
  assign f1596_rst = rst;
  // Bindings to f1596

  // f1598
  logic [0:0] f1598_wen;
  logic [31:0] f1598_wdata;
  logic [0:0] f1598_clk;
  logic [0:0] f1598_rst;
  logic [31:0] f1598_rdata;
  sr_buffer_32_1 f1598(.wen(f1598_wen), .wdata(f1598_wdata), .clk(f1598_clk), .rst(f1598_rst), .rdata(f1598_rdata));
  assign f1598_clk = clk;
  assign f1598_rst = rst;
  // Bindings to f1598

  // f1600
  logic [0:0] f1600_wen;
  logic [31:0] f1600_wdata;
  logic [0:0] f1600_clk;
  logic [0:0] f1600_rst;
  logic [31:0] f1600_rdata;
  sr_buffer_32_1 f1600(.wen(f1600_wen), .wdata(f1600_wdata), .clk(f1600_clk), .rst(f1600_rst), .rdata(f1600_rdata));
  assign f1600_clk = clk;
  assign f1600_rst = rst;
  // Bindings to f1600

  // f1602
  logic [0:0] f1602_wen;
  logic [31:0] f1602_wdata;
  logic [0:0] f1602_clk;
  logic [0:0] f1602_rst;
  logic [31:0] f1602_rdata;
  sr_buffer_32_1 f1602(.wen(f1602_wen), .wdata(f1602_wdata), .clk(f1602_clk), .rst(f1602_rst), .rdata(f1602_rdata));
  assign f1602_clk = clk;
  assign f1602_rst = rst;
  // Bindings to f1602

  // f1604
  logic [0:0] f1604_wen;
  logic [31:0] f1604_wdata;
  logic [0:0] f1604_clk;
  logic [0:0] f1604_rst;
  logic [31:0] f1604_rdata;
  sr_buffer_32_1 f1604(.wen(f1604_wen), .wdata(f1604_wdata), .clk(f1604_clk), .rst(f1604_rst), .rdata(f1604_rdata));
  assign f1604_clk = clk;
  assign f1604_rst = rst;
  // Bindings to f1604

  // f1606
  logic [0:0] f1606_wen;
  logic [31:0] f1606_wdata;
  logic [0:0] f1606_clk;
  logic [0:0] f1606_rst;
  logic [31:0] f1606_rdata;
  sr_buffer_32_1 f1606(.wen(f1606_wen), .wdata(f1606_wdata), .clk(f1606_clk), .rst(f1606_rst), .rdata(f1606_rdata));
  assign f1606_clk = clk;
  assign f1606_rst = rst;
  // Bindings to f1606

  // f1608
  logic [0:0] f1608_wen;
  logic [31:0] f1608_wdata;
  logic [0:0] f1608_clk;
  logic [0:0] f1608_rst;
  logic [31:0] f1608_rdata;
  sr_buffer_32_1 f1608(.wen(f1608_wen), .wdata(f1608_wdata), .clk(f1608_clk), .rst(f1608_rst), .rdata(f1608_rdata));
  assign f1608_clk = clk;
  assign f1608_rst = rst;
  // Bindings to f1608

  // f1610
  logic [0:0] f1610_wen;
  logic [31:0] f1610_wdata;
  logic [0:0] f1610_clk;
  logic [0:0] f1610_rst;
  logic [31:0] f1610_rdata;
  sr_buffer_32_1 f1610(.wen(f1610_wen), .wdata(f1610_wdata), .clk(f1610_clk), .rst(f1610_rst), .rdata(f1610_rdata));
  assign f1610_clk = clk;
  assign f1610_rst = rst;
  // Bindings to f1610

  // f1612
  logic [0:0] f1612_wen;
  logic [31:0] f1612_wdata;
  logic [0:0] f1612_clk;
  logic [0:0] f1612_rst;
  logic [31:0] f1612_rdata;
  sr_buffer_32_1 f1612(.wen(f1612_wen), .wdata(f1612_wdata), .clk(f1612_clk), .rst(f1612_rst), .rdata(f1612_rdata));
  assign f1612_clk = clk;
  assign f1612_rst = rst;
  // Bindings to f1612

  // f1614
  logic [0:0] f1614_wen;
  logic [31:0] f1614_wdata;
  logic [0:0] f1614_clk;
  logic [0:0] f1614_rst;
  logic [31:0] f1614_rdata;
  sr_buffer_32_1 f1614(.wen(f1614_wen), .wdata(f1614_wdata), .clk(f1614_clk), .rst(f1614_rst), .rdata(f1614_rdata));
  assign f1614_clk = clk;
  assign f1614_rst = rst;
  // Bindings to f1614

  // f1616
  logic [0:0] f1616_wen;
  logic [31:0] f1616_wdata;
  logic [0:0] f1616_clk;
  logic [0:0] f1616_rst;
  logic [31:0] f1616_rdata;
  sr_buffer_32_1 f1616(.wen(f1616_wen), .wdata(f1616_wdata), .clk(f1616_clk), .rst(f1616_rst), .rdata(f1616_rdata));
  assign f1616_clk = clk;
  assign f1616_rst = rst;
  // Bindings to f1616

  // f1618
  logic [0:0] f1618_wen;
  logic [31:0] f1618_wdata;
  logic [0:0] f1618_clk;
  logic [0:0] f1618_rst;
  logic [31:0] f1618_rdata;
  sr_buffer_32_1 f1618(.wen(f1618_wen), .wdata(f1618_wdata), .clk(f1618_clk), .rst(f1618_rst), .rdata(f1618_rdata));
  assign f1618_clk = clk;
  assign f1618_rst = rst;
  // Bindings to f1618

  // f1620
  logic [0:0] f1620_wen;
  logic [31:0] f1620_wdata;
  logic [0:0] f1620_clk;
  logic [0:0] f1620_rst;
  logic [31:0] f1620_rdata;
  sr_buffer_32_1 f1620(.wen(f1620_wen), .wdata(f1620_wdata), .clk(f1620_clk), .rst(f1620_rst), .rdata(f1620_rdata));
  assign f1620_clk = clk;
  assign f1620_rst = rst;
  // Bindings to f1620

  // f1622
  logic [0:0] f1622_wen;
  logic [31:0] f1622_wdata;
  logic [0:0] f1622_clk;
  logic [0:0] f1622_rst;
  logic [31:0] f1622_rdata;
  sr_buffer_32_1 f1622(.wen(f1622_wen), .wdata(f1622_wdata), .clk(f1622_clk), .rst(f1622_rst), .rdata(f1622_rdata));
  assign f1622_clk = clk;
  assign f1622_rst = rst;
  // Bindings to f1622

  // f1624
  logic [0:0] f1624_wen;
  logic [31:0] f1624_wdata;
  logic [0:0] f1624_clk;
  logic [0:0] f1624_rst;
  logic [31:0] f1624_rdata;
  sr_buffer_32_1 f1624(.wen(f1624_wen), .wdata(f1624_wdata), .clk(f1624_clk), .rst(f1624_rst), .rdata(f1624_rdata));
  assign f1624_clk = clk;
  assign f1624_rst = rst;
  // Bindings to f1624

  // f1626
  logic [0:0] f1626_wen;
  logic [31:0] f1626_wdata;
  logic [0:0] f1626_clk;
  logic [0:0] f1626_rst;
  logic [31:0] f1626_rdata;
  sr_buffer_32_1 f1626(.wen(f1626_wen), .wdata(f1626_wdata), .clk(f1626_clk), .rst(f1626_rst), .rdata(f1626_rdata));
  assign f1626_clk = clk;
  assign f1626_rst = rst;
  // Bindings to f1626

  // f1628
  logic [0:0] f1628_wen;
  logic [31:0] f1628_wdata;
  logic [0:0] f1628_clk;
  logic [0:0] f1628_rst;
  logic [31:0] f1628_rdata;
  sr_buffer_32_1 f1628(.wen(f1628_wen), .wdata(f1628_wdata), .clk(f1628_clk), .rst(f1628_rst), .rdata(f1628_rdata));
  assign f1628_clk = clk;
  assign f1628_rst = rst;
  // Bindings to f1628

  // f1630
  logic [0:0] f1630_wen;
  logic [31:0] f1630_wdata;
  logic [0:0] f1630_clk;
  logic [0:0] f1630_rst;
  logic [31:0] f1630_rdata;
  sr_buffer_32_1 f1630(.wen(f1630_wen), .wdata(f1630_wdata), .clk(f1630_clk), .rst(f1630_rst), .rdata(f1630_rdata));
  assign f1630_clk = clk;
  assign f1630_rst = rst;
  // Bindings to f1630

  // f1632
  logic [0:0] f1632_wen;
  logic [31:0] f1632_wdata;
  logic [0:0] f1632_clk;
  logic [0:0] f1632_rst;
  logic [31:0] f1632_rdata;
  sr_buffer_32_1 f1632(.wen(f1632_wen), .wdata(f1632_wdata), .clk(f1632_clk), .rst(f1632_rst), .rdata(f1632_rdata));
  assign f1632_clk = clk;
  assign f1632_rst = rst;
  // Bindings to f1632

  // f1634
  logic [0:0] f1634_wen;
  logic [31:0] f1634_wdata;
  logic [0:0] f1634_clk;
  logic [0:0] f1634_rst;
  logic [31:0] f1634_rdata;
  sr_buffer_32_1 f1634(.wen(f1634_wen), .wdata(f1634_wdata), .clk(f1634_clk), .rst(f1634_rst), .rdata(f1634_rdata));
  assign f1634_clk = clk;
  assign f1634_rst = rst;
  // Bindings to f1634

  // f1636
  logic [0:0] f1636_wen;
  logic [31:0] f1636_wdata;
  logic [0:0] f1636_clk;
  logic [0:0] f1636_rst;
  logic [31:0] f1636_rdata;
  sr_buffer_32_1 f1636(.wen(f1636_wen), .wdata(f1636_wdata), .clk(f1636_clk), .rst(f1636_rst), .rdata(f1636_rdata));
  assign f1636_clk = clk;
  assign f1636_rst = rst;
  // Bindings to f1636

  // f1638
  logic [0:0] f1638_wen;
  logic [31:0] f1638_wdata;
  logic [0:0] f1638_clk;
  logic [0:0] f1638_rst;
  logic [31:0] f1638_rdata;
  sr_buffer_32_1 f1638(.wen(f1638_wen), .wdata(f1638_wdata), .clk(f1638_clk), .rst(f1638_rst), .rdata(f1638_rdata));
  assign f1638_clk = clk;
  assign f1638_rst = rst;
  // Bindings to f1638

  // f1640
  logic [0:0] f1640_wen;
  logic [31:0] f1640_wdata;
  logic [0:0] f1640_clk;
  logic [0:0] f1640_rst;
  logic [31:0] f1640_rdata;
  sr_buffer_32_1 f1640(.wen(f1640_wen), .wdata(f1640_wdata), .clk(f1640_clk), .rst(f1640_rst), .rdata(f1640_rdata));
  assign f1640_clk = clk;
  assign f1640_rst = rst;
  // Bindings to f1640

  // f1642
  logic [0:0] f1642_wen;
  logic [31:0] f1642_wdata;
  logic [0:0] f1642_clk;
  logic [0:0] f1642_rst;
  logic [31:0] f1642_rdata;
  sr_buffer_32_1 f1642(.wen(f1642_wen), .wdata(f1642_wdata), .clk(f1642_clk), .rst(f1642_rst), .rdata(f1642_rdata));
  assign f1642_clk = clk;
  assign f1642_rst = rst;
  // Bindings to f1642

  // f1644
  logic [0:0] f1644_wen;
  logic [31:0] f1644_wdata;
  logic [0:0] f1644_clk;
  logic [0:0] f1644_rst;
  logic [31:0] f1644_rdata;
  sr_buffer_32_1 f1644(.wen(f1644_wen), .wdata(f1644_wdata), .clk(f1644_clk), .rst(f1644_rst), .rdata(f1644_rdata));
  assign f1644_clk = clk;
  assign f1644_rst = rst;
  // Bindings to f1644

  // f1646
  logic [0:0] f1646_wen;
  logic [31:0] f1646_wdata;
  logic [0:0] f1646_clk;
  logic [0:0] f1646_rst;
  logic [31:0] f1646_rdata;
  sr_buffer_32_1 f1646(.wen(f1646_wen), .wdata(f1646_wdata), .clk(f1646_clk), .rst(f1646_rst), .rdata(f1646_rdata));
  assign f1646_clk = clk;
  assign f1646_rst = rst;
  // Bindings to f1646

  // f1648
  logic [0:0] f1648_wen;
  logic [31:0] f1648_wdata;
  logic [0:0] f1648_clk;
  logic [0:0] f1648_rst;
  logic [31:0] f1648_rdata;
  sr_buffer_32_1 f1648(.wen(f1648_wen), .wdata(f1648_wdata), .clk(f1648_clk), .rst(f1648_rst), .rdata(f1648_rdata));
  assign f1648_clk = clk;
  assign f1648_rst = rst;
  // Bindings to f1648

  // f1650
  logic [0:0] f1650_wen;
  logic [31:0] f1650_wdata;
  logic [0:0] f1650_clk;
  logic [0:0] f1650_rst;
  logic [31:0] f1650_rdata;
  sr_buffer_32_1 f1650(.wen(f1650_wen), .wdata(f1650_wdata), .clk(f1650_clk), .rst(f1650_rst), .rdata(f1650_rdata));
  assign f1650_clk = clk;
  assign f1650_rst = rst;
  // Bindings to f1650

  // f1652
  logic [0:0] f1652_wen;
  logic [31:0] f1652_wdata;
  logic [0:0] f1652_clk;
  logic [0:0] f1652_rst;
  logic [31:0] f1652_rdata;
  sr_buffer_32_1 f1652(.wen(f1652_wen), .wdata(f1652_wdata), .clk(f1652_clk), .rst(f1652_rst), .rdata(f1652_rdata));
  assign f1652_clk = clk;
  assign f1652_rst = rst;
  // Bindings to f1652

  // f1654
  logic [0:0] f1654_wen;
  logic [31:0] f1654_wdata;
  logic [0:0] f1654_clk;
  logic [0:0] f1654_rst;
  logic [31:0] f1654_rdata;
  sr_buffer_32_1 f1654(.wen(f1654_wen), .wdata(f1654_wdata), .clk(f1654_clk), .rst(f1654_rst), .rdata(f1654_rdata));
  assign f1654_clk = clk;
  assign f1654_rst = rst;
  // Bindings to f1654

  // f1656
  logic [0:0] f1656_wen;
  logic [31:0] f1656_wdata;
  logic [0:0] f1656_clk;
  logic [0:0] f1656_rst;
  logic [31:0] f1656_rdata;
  sr_buffer_32_1 f1656(.wen(f1656_wen), .wdata(f1656_wdata), .clk(f1656_clk), .rst(f1656_rst), .rdata(f1656_rdata));
  assign f1656_clk = clk;
  assign f1656_rst = rst;
  // Bindings to f1656

  // f1658
  logic [0:0] f1658_wen;
  logic [31:0] f1658_wdata;
  logic [0:0] f1658_clk;
  logic [0:0] f1658_rst;
  logic [31:0] f1658_rdata;
  sr_buffer_32_1 f1658(.wen(f1658_wen), .wdata(f1658_wdata), .clk(f1658_clk), .rst(f1658_rst), .rdata(f1658_rdata));
  assign f1658_clk = clk;
  assign f1658_rst = rst;
  // Bindings to f1658

  // f1660
  logic [0:0] f1660_wen;
  logic [31:0] f1660_wdata;
  logic [0:0] f1660_clk;
  logic [0:0] f1660_rst;
  logic [31:0] f1660_rdata;
  sr_buffer_32_1 f1660(.wen(f1660_wen), .wdata(f1660_wdata), .clk(f1660_clk), .rst(f1660_rst), .rdata(f1660_rdata));
  assign f1660_clk = clk;
  assign f1660_rst = rst;
  // Bindings to f1660

  // f1662
  logic [0:0] f1662_wen;
  logic [31:0] f1662_wdata;
  logic [0:0] f1662_clk;
  logic [0:0] f1662_rst;
  logic [31:0] f1662_rdata;
  sr_buffer_32_1 f1662(.wen(f1662_wen), .wdata(f1662_wdata), .clk(f1662_clk), .rst(f1662_rst), .rdata(f1662_rdata));
  assign f1662_clk = clk;
  assign f1662_rst = rst;
  // Bindings to f1662

  // f1664
  logic [0:0] f1664_wen;
  logic [31:0] f1664_wdata;
  logic [0:0] f1664_clk;
  logic [0:0] f1664_rst;
  logic [31:0] f1664_rdata;
  sr_buffer_32_1 f1664(.wen(f1664_wen), .wdata(f1664_wdata), .clk(f1664_clk), .rst(f1664_rst), .rdata(f1664_rdata));
  assign f1664_clk = clk;
  assign f1664_rst = rst;
  // Bindings to f1664

  // f1666
  logic [0:0] f1666_wen;
  logic [31:0] f1666_wdata;
  logic [0:0] f1666_clk;
  logic [0:0] f1666_rst;
  logic [31:0] f1666_rdata;
  sr_buffer_32_1 f1666(.wen(f1666_wen), .wdata(f1666_wdata), .clk(f1666_clk), .rst(f1666_rst), .rdata(f1666_rdata));
  assign f1666_clk = clk;
  assign f1666_rst = rst;
  // Bindings to f1666

  // f1668
  logic [0:0] f1668_wen;
  logic [31:0] f1668_wdata;
  logic [0:0] f1668_clk;
  logic [0:0] f1668_rst;
  logic [31:0] f1668_rdata;
  sr_buffer_32_1 f1668(.wen(f1668_wen), .wdata(f1668_wdata), .clk(f1668_clk), .rst(f1668_rst), .rdata(f1668_rdata));
  assign f1668_clk = clk;
  assign f1668_rst = rst;
  // Bindings to f1668

  // f1670
  logic [0:0] f1670_wen;
  logic [31:0] f1670_wdata;
  logic [0:0] f1670_clk;
  logic [0:0] f1670_rst;
  logic [31:0] f1670_rdata;
  sr_buffer_32_1 f1670(.wen(f1670_wen), .wdata(f1670_wdata), .clk(f1670_clk), .rst(f1670_rst), .rdata(f1670_rdata));
  assign f1670_clk = clk;
  assign f1670_rst = rst;
  // Bindings to f1670

  // f1672
  logic [0:0] f1672_wen;
  logic [31:0] f1672_wdata;
  logic [0:0] f1672_clk;
  logic [0:0] f1672_rst;
  logic [31:0] f1672_rdata;
  sr_buffer_32_1 f1672(.wen(f1672_wen), .wdata(f1672_wdata), .clk(f1672_clk), .rst(f1672_rst), .rdata(f1672_rdata));
  assign f1672_clk = clk;
  assign f1672_rst = rst;
  // Bindings to f1672

  // f1674
  logic [0:0] f1674_wen;
  logic [31:0] f1674_wdata;
  logic [0:0] f1674_clk;
  logic [0:0] f1674_rst;
  logic [31:0] f1674_rdata;
  sr_buffer_32_1 f1674(.wen(f1674_wen), .wdata(f1674_wdata), .clk(f1674_clk), .rst(f1674_rst), .rdata(f1674_rdata));
  assign f1674_clk = clk;
  assign f1674_rst = rst;
  // Bindings to f1674

  // f1676
  logic [0:0] f1676_wen;
  logic [31:0] f1676_wdata;
  logic [0:0] f1676_clk;
  logic [0:0] f1676_rst;
  logic [31:0] f1676_rdata;
  sr_buffer_32_1 f1676(.wen(f1676_wen), .wdata(f1676_wdata), .clk(f1676_clk), .rst(f1676_rst), .rdata(f1676_rdata));
  assign f1676_clk = clk;
  assign f1676_rst = rst;
  // Bindings to f1676

  // f1678
  logic [0:0] f1678_wen;
  logic [31:0] f1678_wdata;
  logic [0:0] f1678_clk;
  logic [0:0] f1678_rst;
  logic [31:0] f1678_rdata;
  sr_buffer_32_1 f1678(.wen(f1678_wen), .wdata(f1678_wdata), .clk(f1678_clk), .rst(f1678_rst), .rdata(f1678_rdata));
  assign f1678_clk = clk;
  assign f1678_rst = rst;
  // Bindings to f1678

  // f1680
  logic [0:0] f1680_wen;
  logic [31:0] f1680_wdata;
  logic [0:0] f1680_clk;
  logic [0:0] f1680_rst;
  logic [31:0] f1680_rdata;
  sr_buffer_32_1 f1680(.wen(f1680_wen), .wdata(f1680_wdata), .clk(f1680_clk), .rst(f1680_rst), .rdata(f1680_rdata));
  assign f1680_clk = clk;
  assign f1680_rst = rst;
  // Bindings to f1680

  // f1682
  logic [0:0] f1682_wen;
  logic [31:0] f1682_wdata;
  logic [0:0] f1682_clk;
  logic [0:0] f1682_rst;
  logic [31:0] f1682_rdata;
  sr_buffer_32_1 f1682(.wen(f1682_wen), .wdata(f1682_wdata), .clk(f1682_clk), .rst(f1682_rst), .rdata(f1682_rdata));
  assign f1682_clk = clk;
  assign f1682_rst = rst;
  // Bindings to f1682

  // f1684
  logic [0:0] f1684_wen;
  logic [31:0] f1684_wdata;
  logic [0:0] f1684_clk;
  logic [0:0] f1684_rst;
  logic [31:0] f1684_rdata;
  sr_buffer_32_1 f1684(.wen(f1684_wen), .wdata(f1684_wdata), .clk(f1684_clk), .rst(f1684_rst), .rdata(f1684_rdata));
  assign f1684_clk = clk;
  assign f1684_rst = rst;
  // Bindings to f1684

  // f1686
  logic [0:0] f1686_wen;
  logic [31:0] f1686_wdata;
  logic [0:0] f1686_clk;
  logic [0:0] f1686_rst;
  logic [31:0] f1686_rdata;
  sr_buffer_32_1 f1686(.wen(f1686_wen), .wdata(f1686_wdata), .clk(f1686_clk), .rst(f1686_rst), .rdata(f1686_rdata));
  assign f1686_clk = clk;
  assign f1686_rst = rst;
  // Bindings to f1686

  // f1688
  logic [0:0] f1688_wen;
  logic [31:0] f1688_wdata;
  logic [0:0] f1688_clk;
  logic [0:0] f1688_rst;
  logic [31:0] f1688_rdata;
  sr_buffer_32_1 f1688(.wen(f1688_wen), .wdata(f1688_wdata), .clk(f1688_clk), .rst(f1688_rst), .rdata(f1688_rdata));
  assign f1688_clk = clk;
  assign f1688_rst = rst;
  // Bindings to f1688

  // f1690
  logic [0:0] f1690_wen;
  logic [31:0] f1690_wdata;
  logic [0:0] f1690_clk;
  logic [0:0] f1690_rst;
  logic [31:0] f1690_rdata;
  sr_buffer_32_1 f1690(.wen(f1690_wen), .wdata(f1690_wdata), .clk(f1690_clk), .rst(f1690_rst), .rdata(f1690_rdata));
  assign f1690_clk = clk;
  assign f1690_rst = rst;
  // Bindings to f1690

  // f1692
  logic [0:0] f1692_wen;
  logic [31:0] f1692_wdata;
  logic [0:0] f1692_clk;
  logic [0:0] f1692_rst;
  logic [31:0] f1692_rdata;
  sr_buffer_32_1 f1692(.wen(f1692_wen), .wdata(f1692_wdata), .clk(f1692_clk), .rst(f1692_rst), .rdata(f1692_rdata));
  assign f1692_clk = clk;
  assign f1692_rst = rst;
  // Bindings to f1692

  // f1694
  logic [0:0] f1694_wen;
  logic [31:0] f1694_wdata;
  logic [0:0] f1694_clk;
  logic [0:0] f1694_rst;
  logic [31:0] f1694_rdata;
  sr_buffer_32_1 f1694(.wen(f1694_wen), .wdata(f1694_wdata), .clk(f1694_clk), .rst(f1694_rst), .rdata(f1694_rdata));
  assign f1694_clk = clk;
  assign f1694_rst = rst;
  // Bindings to f1694

  // f1696
  logic [0:0] f1696_wen;
  logic [31:0] f1696_wdata;
  logic [0:0] f1696_clk;
  logic [0:0] f1696_rst;
  logic [31:0] f1696_rdata;
  sr_buffer_32_1 f1696(.wen(f1696_wen), .wdata(f1696_wdata), .clk(f1696_clk), .rst(f1696_rst), .rdata(f1696_rdata));
  assign f1696_clk = clk;
  assign f1696_rst = rst;
  // Bindings to f1696

  // f1698
  logic [0:0] f1698_wen;
  logic [31:0] f1698_wdata;
  logic [0:0] f1698_clk;
  logic [0:0] f1698_rst;
  logic [31:0] f1698_rdata;
  sr_buffer_32_1 f1698(.wen(f1698_wen), .wdata(f1698_wdata), .clk(f1698_clk), .rst(f1698_rst), .rdata(f1698_rdata));
  assign f1698_clk = clk;
  assign f1698_rst = rst;
  // Bindings to f1698

  // f1700
  logic [0:0] f1700_wen;
  logic [31:0] f1700_wdata;
  logic [0:0] f1700_clk;
  logic [0:0] f1700_rst;
  logic [31:0] f1700_rdata;
  sr_buffer_32_1 f1700(.wen(f1700_wen), .wdata(f1700_wdata), .clk(f1700_clk), .rst(f1700_rst), .rdata(f1700_rdata));
  assign f1700_clk = clk;
  assign f1700_rst = rst;
  // Bindings to f1700

  // f1702
  logic [0:0] f1702_wen;
  logic [31:0] f1702_wdata;
  logic [0:0] f1702_clk;
  logic [0:0] f1702_rst;
  logic [31:0] f1702_rdata;
  sr_buffer_32_1 f1702(.wen(f1702_wen), .wdata(f1702_wdata), .clk(f1702_clk), .rst(f1702_rst), .rdata(f1702_rdata));
  assign f1702_clk = clk;
  assign f1702_rst = rst;
  // Bindings to f1702

  // f1704
  logic [0:0] f1704_wen;
  logic [31:0] f1704_wdata;
  logic [0:0] f1704_clk;
  logic [0:0] f1704_rst;
  logic [31:0] f1704_rdata;
  sr_buffer_32_1 f1704(.wen(f1704_wen), .wdata(f1704_wdata), .clk(f1704_clk), .rst(f1704_rst), .rdata(f1704_rdata));
  assign f1704_clk = clk;
  assign f1704_rst = rst;
  // Bindings to f1704

  // f1706
  logic [0:0] f1706_wen;
  logic [31:0] f1706_wdata;
  logic [0:0] f1706_clk;
  logic [0:0] f1706_rst;
  logic [31:0] f1706_rdata;
  sr_buffer_32_1 f1706(.wen(f1706_wen), .wdata(f1706_wdata), .clk(f1706_clk), .rst(f1706_rst), .rdata(f1706_rdata));
  assign f1706_clk = clk;
  assign f1706_rst = rst;
  // Bindings to f1706

  // f1708
  logic [0:0] f1708_wen;
  logic [31:0] f1708_wdata;
  logic [0:0] f1708_clk;
  logic [0:0] f1708_rst;
  logic [31:0] f1708_rdata;
  sr_buffer_32_1 f1708(.wen(f1708_wen), .wdata(f1708_wdata), .clk(f1708_clk), .rst(f1708_rst), .rdata(f1708_rdata));
  assign f1708_clk = clk;
  assign f1708_rst = rst;
  // Bindings to f1708

  // f1710
  logic [0:0] f1710_wen;
  logic [31:0] f1710_wdata;
  logic [0:0] f1710_clk;
  logic [0:0] f1710_rst;
  logic [31:0] f1710_rdata;
  sr_buffer_32_1 f1710(.wen(f1710_wen), .wdata(f1710_wdata), .clk(f1710_clk), .rst(f1710_rst), .rdata(f1710_rdata));
  assign f1710_clk = clk;
  assign f1710_rst = rst;
  // Bindings to f1710

  // f1712
  logic [0:0] f1712_wen;
  logic [31:0] f1712_wdata;
  logic [0:0] f1712_clk;
  logic [0:0] f1712_rst;
  logic [31:0] f1712_rdata;
  sr_buffer_32_1 f1712(.wen(f1712_wen), .wdata(f1712_wdata), .clk(f1712_clk), .rst(f1712_rst), .rdata(f1712_rdata));
  assign f1712_clk = clk;
  assign f1712_rst = rst;
  // Bindings to f1712

  // f1714
  logic [0:0] f1714_wen;
  logic [31:0] f1714_wdata;
  logic [0:0] f1714_clk;
  logic [0:0] f1714_rst;
  logic [31:0] f1714_rdata;
  sr_buffer_32_1 f1714(.wen(f1714_wen), .wdata(f1714_wdata), .clk(f1714_clk), .rst(f1714_rst), .rdata(f1714_rdata));
  assign f1714_clk = clk;
  assign f1714_rst = rst;
  // Bindings to f1714

  // f1716
  logic [0:0] f1716_wen;
  logic [31:0] f1716_wdata;
  logic [0:0] f1716_clk;
  logic [0:0] f1716_rst;
  logic [31:0] f1716_rdata;
  sr_buffer_32_1 f1716(.wen(f1716_wen), .wdata(f1716_wdata), .clk(f1716_clk), .rst(f1716_rst), .rdata(f1716_rdata));
  assign f1716_clk = clk;
  assign f1716_rst = rst;
  // Bindings to f1716

  // f1718
  logic [0:0] f1718_wen;
  logic [31:0] f1718_wdata;
  logic [0:0] f1718_clk;
  logic [0:0] f1718_rst;
  logic [31:0] f1718_rdata;
  sr_buffer_32_1 f1718(.wen(f1718_wen), .wdata(f1718_wdata), .clk(f1718_clk), .rst(f1718_rst), .rdata(f1718_rdata));
  assign f1718_clk = clk;
  assign f1718_rst = rst;
  // Bindings to f1718

  // f1720
  logic [0:0] f1720_wen;
  logic [31:0] f1720_wdata;
  logic [0:0] f1720_clk;
  logic [0:0] f1720_rst;
  logic [31:0] f1720_rdata;
  sr_buffer_32_1 f1720(.wen(f1720_wen), .wdata(f1720_wdata), .clk(f1720_clk), .rst(f1720_rst), .rdata(f1720_rdata));
  assign f1720_clk = clk;
  assign f1720_rst = rst;
  // Bindings to f1720

  // f1722
  logic [0:0] f1722_wen;
  logic [31:0] f1722_wdata;
  logic [0:0] f1722_clk;
  logic [0:0] f1722_rst;
  logic [31:0] f1722_rdata;
  sr_buffer_32_1 f1722(.wen(f1722_wen), .wdata(f1722_wdata), .clk(f1722_clk), .rst(f1722_rst), .rdata(f1722_rdata));
  assign f1722_clk = clk;
  assign f1722_rst = rst;
  // Bindings to f1722

  // f1724
  logic [0:0] f1724_wen;
  logic [31:0] f1724_wdata;
  logic [0:0] f1724_clk;
  logic [0:0] f1724_rst;
  logic [31:0] f1724_rdata;
  sr_buffer_32_1 f1724(.wen(f1724_wen), .wdata(f1724_wdata), .clk(f1724_clk), .rst(f1724_rst), .rdata(f1724_rdata));
  assign f1724_clk = clk;
  assign f1724_rst = rst;
  // Bindings to f1724

  // f1726
  logic [0:0] f1726_wen;
  logic [31:0] f1726_wdata;
  logic [0:0] f1726_clk;
  logic [0:0] f1726_rst;
  logic [31:0] f1726_rdata;
  sr_buffer_32_1 f1726(.wen(f1726_wen), .wdata(f1726_wdata), .clk(f1726_clk), .rst(f1726_rst), .rdata(f1726_rdata));
  assign f1726_clk = clk;
  assign f1726_rst = rst;
  // Bindings to f1726

  // f1728
  logic [0:0] f1728_wen;
  logic [31:0] f1728_wdata;
  logic [0:0] f1728_clk;
  logic [0:0] f1728_rst;
  logic [31:0] f1728_rdata;
  sr_buffer_32_1 f1728(.wen(f1728_wen), .wdata(f1728_wdata), .clk(f1728_clk), .rst(f1728_rst), .rdata(f1728_rdata));
  assign f1728_clk = clk;
  assign f1728_rst = rst;
  // Bindings to f1728

  // f1730
  logic [0:0] f1730_wen;
  logic [31:0] f1730_wdata;
  logic [0:0] f1730_clk;
  logic [0:0] f1730_rst;
  logic [31:0] f1730_rdata;
  sr_buffer_32_1 f1730(.wen(f1730_wen), .wdata(f1730_wdata), .clk(f1730_clk), .rst(f1730_rst), .rdata(f1730_rdata));
  assign f1730_clk = clk;
  assign f1730_rst = rst;
  // Bindings to f1730

  // f1732
  logic [0:0] f1732_wen;
  logic [31:0] f1732_wdata;
  logic [0:0] f1732_clk;
  logic [0:0] f1732_rst;
  logic [31:0] f1732_rdata;
  sr_buffer_32_1 f1732(.wen(f1732_wen), .wdata(f1732_wdata), .clk(f1732_clk), .rst(f1732_rst), .rdata(f1732_rdata));
  assign f1732_clk = clk;
  assign f1732_rst = rst;
  // Bindings to f1732

  // f1734
  logic [0:0] f1734_wen;
  logic [31:0] f1734_wdata;
  logic [0:0] f1734_clk;
  logic [0:0] f1734_rst;
  logic [31:0] f1734_rdata;
  sr_buffer_32_1 f1734(.wen(f1734_wen), .wdata(f1734_wdata), .clk(f1734_clk), .rst(f1734_rst), .rdata(f1734_rdata));
  assign f1734_clk = clk;
  assign f1734_rst = rst;
  // Bindings to f1734

  // f1736
  logic [0:0] f1736_wen;
  logic [31:0] f1736_wdata;
  logic [0:0] f1736_clk;
  logic [0:0] f1736_rst;
  logic [31:0] f1736_rdata;
  sr_buffer_32_1 f1736(.wen(f1736_wen), .wdata(f1736_wdata), .clk(f1736_clk), .rst(f1736_rst), .rdata(f1736_rdata));
  assign f1736_clk = clk;
  assign f1736_rst = rst;
  // Bindings to f1736

  // f1738
  logic [0:0] f1738_wen;
  logic [31:0] f1738_wdata;
  logic [0:0] f1738_clk;
  logic [0:0] f1738_rst;
  logic [31:0] f1738_rdata;
  sr_buffer_32_1 f1738(.wen(f1738_wen), .wdata(f1738_wdata), .clk(f1738_clk), .rst(f1738_rst), .rdata(f1738_rdata));
  assign f1738_clk = clk;
  assign f1738_rst = rst;
  // Bindings to f1738

  // f1740
  logic [0:0] f1740_wen;
  logic [31:0] f1740_wdata;
  logic [0:0] f1740_clk;
  logic [0:0] f1740_rst;
  logic [31:0] f1740_rdata;
  sr_buffer_32_1 f1740(.wen(f1740_wen), .wdata(f1740_wdata), .clk(f1740_clk), .rst(f1740_rst), .rdata(f1740_rdata));
  assign f1740_clk = clk;
  assign f1740_rst = rst;
  // Bindings to f1740

  // f1742
  logic [0:0] f1742_wen;
  logic [31:0] f1742_wdata;
  logic [0:0] f1742_clk;
  logic [0:0] f1742_rst;
  logic [31:0] f1742_rdata;
  sr_buffer_32_1 f1742(.wen(f1742_wen), .wdata(f1742_wdata), .clk(f1742_clk), .rst(f1742_rst), .rdata(f1742_rdata));
  assign f1742_clk = clk;
  assign f1742_rst = rst;
  // Bindings to f1742

  // f1744
  logic [0:0] f1744_wen;
  logic [31:0] f1744_wdata;
  logic [0:0] f1744_clk;
  logic [0:0] f1744_rst;
  logic [31:0] f1744_rdata;
  sr_buffer_32_1 f1744(.wen(f1744_wen), .wdata(f1744_wdata), .clk(f1744_clk), .rst(f1744_rst), .rdata(f1744_rdata));
  assign f1744_clk = clk;
  assign f1744_rst = rst;
  // Bindings to f1744

  // f1746
  logic [0:0] f1746_wen;
  logic [31:0] f1746_wdata;
  logic [0:0] f1746_clk;
  logic [0:0] f1746_rst;
  logic [31:0] f1746_rdata;
  sr_buffer_32_1 f1746(.wen(f1746_wen), .wdata(f1746_wdata), .clk(f1746_clk), .rst(f1746_rst), .rdata(f1746_rdata));
  assign f1746_clk = clk;
  assign f1746_rst = rst;
  // Bindings to f1746

  // f1748
  logic [0:0] f1748_wen;
  logic [31:0] f1748_wdata;
  logic [0:0] f1748_clk;
  logic [0:0] f1748_rst;
  logic [31:0] f1748_rdata;
  sr_buffer_32_1 f1748(.wen(f1748_wen), .wdata(f1748_wdata), .clk(f1748_clk), .rst(f1748_rst), .rdata(f1748_rdata));
  assign f1748_clk = clk;
  assign f1748_rst = rst;
  // Bindings to f1748

  // f1750
  logic [0:0] f1750_wen;
  logic [31:0] f1750_wdata;
  logic [0:0] f1750_clk;
  logic [0:0] f1750_rst;
  logic [31:0] f1750_rdata;
  sr_buffer_32_1 f1750(.wen(f1750_wen), .wdata(f1750_wdata), .clk(f1750_clk), .rst(f1750_rst), .rdata(f1750_rdata));
  assign f1750_clk = clk;
  assign f1750_rst = rst;
  // Bindings to f1750

  // f1752
  logic [0:0] f1752_wen;
  logic [31:0] f1752_wdata;
  logic [0:0] f1752_clk;
  logic [0:0] f1752_rst;
  logic [31:0] f1752_rdata;
  sr_buffer_32_1 f1752(.wen(f1752_wen), .wdata(f1752_wdata), .clk(f1752_clk), .rst(f1752_rst), .rdata(f1752_rdata));
  assign f1752_clk = clk;
  assign f1752_rst = rst;
  // Bindings to f1752

  // f1754
  logic [0:0] f1754_wen;
  logic [31:0] f1754_wdata;
  logic [0:0] f1754_clk;
  logic [0:0] f1754_rst;
  logic [31:0] f1754_rdata;
  sr_buffer_32_1 f1754(.wen(f1754_wen), .wdata(f1754_wdata), .clk(f1754_clk), .rst(f1754_rst), .rdata(f1754_rdata));
  assign f1754_clk = clk;
  assign f1754_rst = rst;
  // Bindings to f1754

  // f1756
  logic [0:0] f1756_wen;
  logic [31:0] f1756_wdata;
  logic [0:0] f1756_clk;
  logic [0:0] f1756_rst;
  logic [31:0] f1756_rdata;
  sr_buffer_32_1 f1756(.wen(f1756_wen), .wdata(f1756_wdata), .clk(f1756_clk), .rst(f1756_rst), .rdata(f1756_rdata));
  assign f1756_clk = clk;
  assign f1756_rst = rst;
  // Bindings to f1756

  // f1758
  logic [0:0] f1758_wen;
  logic [31:0] f1758_wdata;
  logic [0:0] f1758_clk;
  logic [0:0] f1758_rst;
  logic [31:0] f1758_rdata;
  sr_buffer_32_1 f1758(.wen(f1758_wen), .wdata(f1758_wdata), .clk(f1758_clk), .rst(f1758_rst), .rdata(f1758_rdata));
  assign f1758_clk = clk;
  assign f1758_rst = rst;
  // Bindings to f1758

  // f1760
  logic [0:0] f1760_wen;
  logic [31:0] f1760_wdata;
  logic [0:0] f1760_clk;
  logic [0:0] f1760_rst;
  logic [31:0] f1760_rdata;
  sr_buffer_32_1 f1760(.wen(f1760_wen), .wdata(f1760_wdata), .clk(f1760_clk), .rst(f1760_rst), .rdata(f1760_rdata));
  assign f1760_clk = clk;
  assign f1760_rst = rst;
  // Bindings to f1760

  // f1762
  logic [0:0] f1762_wen;
  logic [31:0] f1762_wdata;
  logic [0:0] f1762_clk;
  logic [0:0] f1762_rst;
  logic [31:0] f1762_rdata;
  sr_buffer_32_1 f1762(.wen(f1762_wen), .wdata(f1762_wdata), .clk(f1762_clk), .rst(f1762_rst), .rdata(f1762_rdata));
  assign f1762_clk = clk;
  assign f1762_rst = rst;
  // Bindings to f1762

  // f1764
  logic [0:0] f1764_wen;
  logic [31:0] f1764_wdata;
  logic [0:0] f1764_clk;
  logic [0:0] f1764_rst;
  logic [31:0] f1764_rdata;
  sr_buffer_32_1 f1764(.wen(f1764_wen), .wdata(f1764_wdata), .clk(f1764_clk), .rst(f1764_rst), .rdata(f1764_rdata));
  assign f1764_clk = clk;
  assign f1764_rst = rst;
  // Bindings to f1764

  // f1766
  logic [0:0] f1766_wen;
  logic [31:0] f1766_wdata;
  logic [0:0] f1766_clk;
  logic [0:0] f1766_rst;
  logic [31:0] f1766_rdata;
  sr_buffer_32_1 f1766(.wen(f1766_wen), .wdata(f1766_wdata), .clk(f1766_clk), .rst(f1766_rst), .rdata(f1766_rdata));
  assign f1766_clk = clk;
  assign f1766_rst = rst;
  // Bindings to f1766

  // f1768
  logic [0:0] f1768_wen;
  logic [31:0] f1768_wdata;
  logic [0:0] f1768_clk;
  logic [0:0] f1768_rst;
  logic [31:0] f1768_rdata;
  sr_buffer_32_1 f1768(.wen(f1768_wen), .wdata(f1768_wdata), .clk(f1768_clk), .rst(f1768_rst), .rdata(f1768_rdata));
  assign f1768_clk = clk;
  assign f1768_rst = rst;
  // Bindings to f1768

  // f1770
  logic [0:0] f1770_wen;
  logic [31:0] f1770_wdata;
  logic [0:0] f1770_clk;
  logic [0:0] f1770_rst;
  logic [31:0] f1770_rdata;
  sr_buffer_32_1 f1770(.wen(f1770_wen), .wdata(f1770_wdata), .clk(f1770_clk), .rst(f1770_rst), .rdata(f1770_rdata));
  assign f1770_clk = clk;
  assign f1770_rst = rst;
  // Bindings to f1770

  // f1772
  logic [0:0] f1772_wen;
  logic [31:0] f1772_wdata;
  logic [0:0] f1772_clk;
  logic [0:0] f1772_rst;
  logic [31:0] f1772_rdata;
  sr_buffer_32_1 f1772(.wen(f1772_wen), .wdata(f1772_wdata), .clk(f1772_clk), .rst(f1772_rst), .rdata(f1772_rdata));
  assign f1772_clk = clk;
  assign f1772_rst = rst;
  // Bindings to f1772

  // f1774
  logic [0:0] f1774_wen;
  logic [31:0] f1774_wdata;
  logic [0:0] f1774_clk;
  logic [0:0] f1774_rst;
  logic [31:0] f1774_rdata;
  sr_buffer_32_1 f1774(.wen(f1774_wen), .wdata(f1774_wdata), .clk(f1774_clk), .rst(f1774_rst), .rdata(f1774_rdata));
  assign f1774_clk = clk;
  assign f1774_rst = rst;
  // Bindings to f1774

  // f1776
  logic [0:0] f1776_wen;
  logic [31:0] f1776_wdata;
  logic [0:0] f1776_clk;
  logic [0:0] f1776_rst;
  logic [31:0] f1776_rdata;
  sr_buffer_32_1 f1776(.wen(f1776_wen), .wdata(f1776_wdata), .clk(f1776_clk), .rst(f1776_rst), .rdata(f1776_rdata));
  assign f1776_clk = clk;
  assign f1776_rst = rst;
  // Bindings to f1776

  // f1778
  logic [0:0] f1778_wen;
  logic [31:0] f1778_wdata;
  logic [0:0] f1778_clk;
  logic [0:0] f1778_rst;
  logic [31:0] f1778_rdata;
  sr_buffer_32_1 f1778(.wen(f1778_wen), .wdata(f1778_wdata), .clk(f1778_clk), .rst(f1778_rst), .rdata(f1778_rdata));
  assign f1778_clk = clk;
  assign f1778_rst = rst;
  // Bindings to f1778

  // f1780
  logic [0:0] f1780_wen;
  logic [31:0] f1780_wdata;
  logic [0:0] f1780_clk;
  logic [0:0] f1780_rst;
  logic [31:0] f1780_rdata;
  sr_buffer_32_1 f1780(.wen(f1780_wen), .wdata(f1780_wdata), .clk(f1780_clk), .rst(f1780_rst), .rdata(f1780_rdata));
  assign f1780_clk = clk;
  assign f1780_rst = rst;
  // Bindings to f1780

  // f1782
  logic [0:0] f1782_wen;
  logic [31:0] f1782_wdata;
  logic [0:0] f1782_clk;
  logic [0:0] f1782_rst;
  logic [31:0] f1782_rdata;
  sr_buffer_32_1 f1782(.wen(f1782_wen), .wdata(f1782_wdata), .clk(f1782_clk), .rst(f1782_rst), .rdata(f1782_rdata));
  assign f1782_clk = clk;
  assign f1782_rst = rst;
  // Bindings to f1782

  // f1784
  logic [0:0] f1784_wen;
  logic [31:0] f1784_wdata;
  logic [0:0] f1784_clk;
  logic [0:0] f1784_rst;
  logic [31:0] f1784_rdata;
  sr_buffer_32_1 f1784(.wen(f1784_wen), .wdata(f1784_wdata), .clk(f1784_clk), .rst(f1784_rst), .rdata(f1784_rdata));
  assign f1784_clk = clk;
  assign f1784_rst = rst;
  // Bindings to f1784

  // f1786
  logic [0:0] f1786_wen;
  logic [31:0] f1786_wdata;
  logic [0:0] f1786_clk;
  logic [0:0] f1786_rst;
  logic [31:0] f1786_rdata;
  sr_buffer_32_1 f1786(.wen(f1786_wen), .wdata(f1786_wdata), .clk(f1786_clk), .rst(f1786_rst), .rdata(f1786_rdata));
  assign f1786_clk = clk;
  assign f1786_rst = rst;
  // Bindings to f1786

  // f1788
  logic [0:0] f1788_wen;
  logic [31:0] f1788_wdata;
  logic [0:0] f1788_clk;
  logic [0:0] f1788_rst;
  logic [31:0] f1788_rdata;
  sr_buffer_32_1 f1788(.wen(f1788_wen), .wdata(f1788_wdata), .clk(f1788_clk), .rst(f1788_rst), .rdata(f1788_rdata));
  assign f1788_clk = clk;
  assign f1788_rst = rst;
  // Bindings to f1788

  // f1790
  logic [0:0] f1790_wen;
  logic [31:0] f1790_wdata;
  logic [0:0] f1790_clk;
  logic [0:0] f1790_rst;
  logic [31:0] f1790_rdata;
  sr_buffer_32_1 f1790(.wen(f1790_wen), .wdata(f1790_wdata), .clk(f1790_clk), .rst(f1790_rst), .rdata(f1790_rdata));
  assign f1790_clk = clk;
  assign f1790_rst = rst;
  // Bindings to f1790

  // f1792
  logic [0:0] f1792_wen;
  logic [31:0] f1792_wdata;
  logic [0:0] f1792_clk;
  logic [0:0] f1792_rst;
  logic [31:0] f1792_rdata;
  sr_buffer_32_1 f1792(.wen(f1792_wen), .wdata(f1792_wdata), .clk(f1792_clk), .rst(f1792_rst), .rdata(f1792_rdata));
  assign f1792_clk = clk;
  assign f1792_rst = rst;
  // Bindings to f1792

  // f1794
  logic [0:0] f1794_wen;
  logic [31:0] f1794_wdata;
  logic [0:0] f1794_clk;
  logic [0:0] f1794_rst;
  logic [31:0] f1794_rdata;
  sr_buffer_32_1 f1794(.wen(f1794_wen), .wdata(f1794_wdata), .clk(f1794_clk), .rst(f1794_rst), .rdata(f1794_rdata));
  assign f1794_clk = clk;
  assign f1794_rst = rst;
  // Bindings to f1794

  // f1796
  logic [0:0] f1796_wen;
  logic [31:0] f1796_wdata;
  logic [0:0] f1796_clk;
  logic [0:0] f1796_rst;
  logic [31:0] f1796_rdata;
  sr_buffer_32_1 f1796(.wen(f1796_wen), .wdata(f1796_wdata), .clk(f1796_clk), .rst(f1796_rst), .rdata(f1796_rdata));
  assign f1796_clk = clk;
  assign f1796_rst = rst;
  // Bindings to f1796

  // f1798
  logic [0:0] f1798_wen;
  logic [31:0] f1798_wdata;
  logic [0:0] f1798_clk;
  logic [0:0] f1798_rst;
  logic [31:0] f1798_rdata;
  sr_buffer_32_1 f1798(.wen(f1798_wen), .wdata(f1798_wdata), .clk(f1798_clk), .rst(f1798_rst), .rdata(f1798_rdata));
  assign f1798_clk = clk;
  assign f1798_rst = rst;
  // Bindings to f1798

  // f1800
  logic [0:0] f1800_wen;
  logic [31:0] f1800_wdata;
  logic [0:0] f1800_clk;
  logic [0:0] f1800_rst;
  logic [31:0] f1800_rdata;
  sr_buffer_32_1 f1800(.wen(f1800_wen), .wdata(f1800_wdata), .clk(f1800_clk), .rst(f1800_rst), .rdata(f1800_rdata));
  assign f1800_clk = clk;
  assign f1800_rst = rst;
  // Bindings to f1800

  // f1802
  logic [0:0] f1802_wen;
  logic [31:0] f1802_wdata;
  logic [0:0] f1802_clk;
  logic [0:0] f1802_rst;
  logic [31:0] f1802_rdata;
  sr_buffer_32_1 f1802(.wen(f1802_wen), .wdata(f1802_wdata), .clk(f1802_clk), .rst(f1802_rst), .rdata(f1802_rdata));
  assign f1802_clk = clk;
  assign f1802_rst = rst;
  // Bindings to f1802

  // f1804
  logic [0:0] f1804_wen;
  logic [31:0] f1804_wdata;
  logic [0:0] f1804_clk;
  logic [0:0] f1804_rst;
  logic [31:0] f1804_rdata;
  sr_buffer_32_1 f1804(.wen(f1804_wen), .wdata(f1804_wdata), .clk(f1804_clk), .rst(f1804_rst), .rdata(f1804_rdata));
  assign f1804_clk = clk;
  assign f1804_rst = rst;
  // Bindings to f1804

  // f1806
  logic [0:0] f1806_wen;
  logic [31:0] f1806_wdata;
  logic [0:0] f1806_clk;
  logic [0:0] f1806_rst;
  logic [31:0] f1806_rdata;
  sr_buffer_32_1 f1806(.wen(f1806_wen), .wdata(f1806_wdata), .clk(f1806_clk), .rst(f1806_rst), .rdata(f1806_rdata));
  assign f1806_clk = clk;
  assign f1806_rst = rst;
  // Bindings to f1806

  // f1808
  logic [0:0] f1808_wen;
  logic [31:0] f1808_wdata;
  logic [0:0] f1808_clk;
  logic [0:0] f1808_rst;
  logic [31:0] f1808_rdata;
  sr_buffer_32_1 f1808(.wen(f1808_wen), .wdata(f1808_wdata), .clk(f1808_clk), .rst(f1808_rst), .rdata(f1808_rdata));
  assign f1808_clk = clk;
  assign f1808_rst = rst;
  // Bindings to f1808

  // f1810
  logic [0:0] f1810_wen;
  logic [31:0] f1810_wdata;
  logic [0:0] f1810_clk;
  logic [0:0] f1810_rst;
  logic [31:0] f1810_rdata;
  sr_buffer_32_1 f1810(.wen(f1810_wen), .wdata(f1810_wdata), .clk(f1810_clk), .rst(f1810_rst), .rdata(f1810_rdata));
  assign f1810_clk = clk;
  assign f1810_rst = rst;
  // Bindings to f1810

  // f1812
  logic [0:0] f1812_wen;
  logic [31:0] f1812_wdata;
  logic [0:0] f1812_clk;
  logic [0:0] f1812_rst;
  logic [31:0] f1812_rdata;
  sr_buffer_32_1 f1812(.wen(f1812_wen), .wdata(f1812_wdata), .clk(f1812_clk), .rst(f1812_rst), .rdata(f1812_rdata));
  assign f1812_clk = clk;
  assign f1812_rst = rst;
  // Bindings to f1812

  // f1814
  logic [0:0] f1814_wen;
  logic [31:0] f1814_wdata;
  logic [0:0] f1814_clk;
  logic [0:0] f1814_rst;
  logic [31:0] f1814_rdata;
  sr_buffer_32_1 f1814(.wen(f1814_wen), .wdata(f1814_wdata), .clk(f1814_clk), .rst(f1814_rst), .rdata(f1814_rdata));
  assign f1814_clk = clk;
  assign f1814_rst = rst;
  // Bindings to f1814

  // f1816
  logic [0:0] f1816_wen;
  logic [31:0] f1816_wdata;
  logic [0:0] f1816_clk;
  logic [0:0] f1816_rst;
  logic [31:0] f1816_rdata;
  sr_buffer_32_1 f1816(.wen(f1816_wen), .wdata(f1816_wdata), .clk(f1816_clk), .rst(f1816_rst), .rdata(f1816_rdata));
  assign f1816_clk = clk;
  assign f1816_rst = rst;
  // Bindings to f1816

  // f1818
  logic [0:0] f1818_wen;
  logic [31:0] f1818_wdata;
  logic [0:0] f1818_clk;
  logic [0:0] f1818_rst;
  logic [31:0] f1818_rdata;
  sr_buffer_32_1 f1818(.wen(f1818_wen), .wdata(f1818_wdata), .clk(f1818_clk), .rst(f1818_rst), .rdata(f1818_rdata));
  assign f1818_clk = clk;
  assign f1818_rst = rst;
  // Bindings to f1818

  // f1820
  logic [0:0] f1820_wen;
  logic [31:0] f1820_wdata;
  logic [0:0] f1820_clk;
  logic [0:0] f1820_rst;
  logic [31:0] f1820_rdata;
  sr_buffer_32_1 f1820(.wen(f1820_wen), .wdata(f1820_wdata), .clk(f1820_clk), .rst(f1820_rst), .rdata(f1820_rdata));
  assign f1820_clk = clk;
  assign f1820_rst = rst;
  // Bindings to f1820

  // f1822
  logic [0:0] f1822_wen;
  logic [31:0] f1822_wdata;
  logic [0:0] f1822_clk;
  logic [0:0] f1822_rst;
  logic [31:0] f1822_rdata;
  sr_buffer_32_1 f1822(.wen(f1822_wen), .wdata(f1822_wdata), .clk(f1822_clk), .rst(f1822_rst), .rdata(f1822_rdata));
  assign f1822_clk = clk;
  assign f1822_rst = rst;
  // Bindings to f1822

  // f1824
  logic [0:0] f1824_wen;
  logic [31:0] f1824_wdata;
  logic [0:0] f1824_clk;
  logic [0:0] f1824_rst;
  logic [31:0] f1824_rdata;
  sr_buffer_32_1 f1824(.wen(f1824_wen), .wdata(f1824_wdata), .clk(f1824_clk), .rst(f1824_rst), .rdata(f1824_rdata));
  assign f1824_clk = clk;
  assign f1824_rst = rst;
  // Bindings to f1824

  // f1826
  logic [0:0] f1826_wen;
  logic [31:0] f1826_wdata;
  logic [0:0] f1826_clk;
  logic [0:0] f1826_rst;
  logic [31:0] f1826_rdata;
  sr_buffer_32_1 f1826(.wen(f1826_wen), .wdata(f1826_wdata), .clk(f1826_clk), .rst(f1826_rst), .rdata(f1826_rdata));
  assign f1826_clk = clk;
  assign f1826_rst = rst;
  // Bindings to f1826

  // f1828
  logic [0:0] f1828_wen;
  logic [31:0] f1828_wdata;
  logic [0:0] f1828_clk;
  logic [0:0] f1828_rst;
  logic [31:0] f1828_rdata;
  sr_buffer_32_1 f1828(.wen(f1828_wen), .wdata(f1828_wdata), .clk(f1828_clk), .rst(f1828_rst), .rdata(f1828_rdata));
  assign f1828_clk = clk;
  assign f1828_rst = rst;
  // Bindings to f1828

  // f1830
  logic [0:0] f1830_wen;
  logic [31:0] f1830_wdata;
  logic [0:0] f1830_clk;
  logic [0:0] f1830_rst;
  logic [31:0] f1830_rdata;
  sr_buffer_32_1 f1830(.wen(f1830_wen), .wdata(f1830_wdata), .clk(f1830_clk), .rst(f1830_rst), .rdata(f1830_rdata));
  assign f1830_clk = clk;
  assign f1830_rst = rst;
  // Bindings to f1830

  // f1832
  logic [0:0] f1832_wen;
  logic [31:0] f1832_wdata;
  logic [0:0] f1832_clk;
  logic [0:0] f1832_rst;
  logic [31:0] f1832_rdata;
  sr_buffer_32_1 f1832(.wen(f1832_wen), .wdata(f1832_wdata), .clk(f1832_clk), .rst(f1832_rst), .rdata(f1832_rdata));
  assign f1832_clk = clk;
  assign f1832_rst = rst;
  // Bindings to f1832

  // f1834
  logic [0:0] f1834_wen;
  logic [31:0] f1834_wdata;
  logic [0:0] f1834_clk;
  logic [0:0] f1834_rst;
  logic [31:0] f1834_rdata;
  sr_buffer_32_1 f1834(.wen(f1834_wen), .wdata(f1834_wdata), .clk(f1834_clk), .rst(f1834_rst), .rdata(f1834_rdata));
  assign f1834_clk = clk;
  assign f1834_rst = rst;
  // Bindings to f1834

  // f1836
  logic [0:0] f1836_wen;
  logic [31:0] f1836_wdata;
  logic [0:0] f1836_clk;
  logic [0:0] f1836_rst;
  logic [31:0] f1836_rdata;
  sr_buffer_32_1 f1836(.wen(f1836_wen), .wdata(f1836_wdata), .clk(f1836_clk), .rst(f1836_rst), .rdata(f1836_rdata));
  assign f1836_clk = clk;
  assign f1836_rst = rst;
  // Bindings to f1836

  // f1838
  logic [0:0] f1838_wen;
  logic [31:0] f1838_wdata;
  logic [0:0] f1838_clk;
  logic [0:0] f1838_rst;
  logic [31:0] f1838_rdata;
  sr_buffer_32_1 f1838(.wen(f1838_wen), .wdata(f1838_wdata), .clk(f1838_clk), .rst(f1838_rst), .rdata(f1838_rdata));
  assign f1838_clk = clk;
  assign f1838_rst = rst;
  // Bindings to f1838

  // f1840
  logic [0:0] f1840_wen;
  logic [31:0] f1840_wdata;
  logic [0:0] f1840_clk;
  logic [0:0] f1840_rst;
  logic [31:0] f1840_rdata;
  sr_buffer_32_1 f1840(.wen(f1840_wen), .wdata(f1840_wdata), .clk(f1840_clk), .rst(f1840_rst), .rdata(f1840_rdata));
  assign f1840_clk = clk;
  assign f1840_rst = rst;
  // Bindings to f1840

  // f1842
  logic [0:0] f1842_wen;
  logic [31:0] f1842_wdata;
  logic [0:0] f1842_clk;
  logic [0:0] f1842_rst;
  logic [31:0] f1842_rdata;
  sr_buffer_32_1 f1842(.wen(f1842_wen), .wdata(f1842_wdata), .clk(f1842_clk), .rst(f1842_rst), .rdata(f1842_rdata));
  assign f1842_clk = clk;
  assign f1842_rst = rst;
  // Bindings to f1842

  // f1844
  logic [0:0] f1844_wen;
  logic [31:0] f1844_wdata;
  logic [0:0] f1844_clk;
  logic [0:0] f1844_rst;
  logic [31:0] f1844_rdata;
  sr_buffer_32_1 f1844(.wen(f1844_wen), .wdata(f1844_wdata), .clk(f1844_clk), .rst(f1844_rst), .rdata(f1844_rdata));
  assign f1844_clk = clk;
  assign f1844_rst = rst;
  // Bindings to f1844

  // f1846
  logic [0:0] f1846_wen;
  logic [31:0] f1846_wdata;
  logic [0:0] f1846_clk;
  logic [0:0] f1846_rst;
  logic [31:0] f1846_rdata;
  sr_buffer_32_1 f1846(.wen(f1846_wen), .wdata(f1846_wdata), .clk(f1846_clk), .rst(f1846_rst), .rdata(f1846_rdata));
  assign f1846_clk = clk;
  assign f1846_rst = rst;
  // Bindings to f1846

  // f1848
  logic [0:0] f1848_wen;
  logic [31:0] f1848_wdata;
  logic [0:0] f1848_clk;
  logic [0:0] f1848_rst;
  logic [31:0] f1848_rdata;
  sr_buffer_32_1 f1848(.wen(f1848_wen), .wdata(f1848_wdata), .clk(f1848_clk), .rst(f1848_rst), .rdata(f1848_rdata));
  assign f1848_clk = clk;
  assign f1848_rst = rst;
  // Bindings to f1848

  // f1850
  logic [0:0] f1850_wen;
  logic [31:0] f1850_wdata;
  logic [0:0] f1850_clk;
  logic [0:0] f1850_rst;
  logic [31:0] f1850_rdata;
  sr_buffer_32_1 f1850(.wen(f1850_wen), .wdata(f1850_wdata), .clk(f1850_clk), .rst(f1850_rst), .rdata(f1850_rdata));
  assign f1850_clk = clk;
  assign f1850_rst = rst;
  // Bindings to f1850

  // f1852
  logic [0:0] f1852_wen;
  logic [31:0] f1852_wdata;
  logic [0:0] f1852_clk;
  logic [0:0] f1852_rst;
  logic [31:0] f1852_rdata;
  sr_buffer_32_1 f1852(.wen(f1852_wen), .wdata(f1852_wdata), .clk(f1852_clk), .rst(f1852_rst), .rdata(f1852_rdata));
  assign f1852_clk = clk;
  assign f1852_rst = rst;
  // Bindings to f1852

  // f1854
  logic [0:0] f1854_wen;
  logic [31:0] f1854_wdata;
  logic [0:0] f1854_clk;
  logic [0:0] f1854_rst;
  logic [31:0] f1854_rdata;
  sr_buffer_32_1 f1854(.wen(f1854_wen), .wdata(f1854_wdata), .clk(f1854_clk), .rst(f1854_rst), .rdata(f1854_rdata));
  assign f1854_clk = clk;
  assign f1854_rst = rst;
  // Bindings to f1854

  // f1856
  logic [0:0] f1856_wen;
  logic [31:0] f1856_wdata;
  logic [0:0] f1856_clk;
  logic [0:0] f1856_rst;
  logic [31:0] f1856_rdata;
  sr_buffer_32_1 f1856(.wen(f1856_wen), .wdata(f1856_wdata), .clk(f1856_clk), .rst(f1856_rst), .rdata(f1856_rdata));
  assign f1856_clk = clk;
  assign f1856_rst = rst;
  // Bindings to f1856

  // f1858
  logic [0:0] f1858_wen;
  logic [31:0] f1858_wdata;
  logic [0:0] f1858_clk;
  logic [0:0] f1858_rst;
  logic [31:0] f1858_rdata;
  sr_buffer_32_1 f1858(.wen(f1858_wen), .wdata(f1858_wdata), .clk(f1858_clk), .rst(f1858_rst), .rdata(f1858_rdata));
  assign f1858_clk = clk;
  assign f1858_rst = rst;
  // Bindings to f1858

  // f1860
  logic [0:0] f1860_wen;
  logic [31:0] f1860_wdata;
  logic [0:0] f1860_clk;
  logic [0:0] f1860_rst;
  logic [31:0] f1860_rdata;
  sr_buffer_32_1 f1860(.wen(f1860_wen), .wdata(f1860_wdata), .clk(f1860_clk), .rst(f1860_rst), .rdata(f1860_rdata));
  assign f1860_clk = clk;
  assign f1860_rst = rst;
  // Bindings to f1860

  // f1862
  logic [0:0] f1862_wen;
  logic [31:0] f1862_wdata;
  logic [0:0] f1862_clk;
  logic [0:0] f1862_rst;
  logic [31:0] f1862_rdata;
  sr_buffer_32_1 f1862(.wen(f1862_wen), .wdata(f1862_wdata), .clk(f1862_clk), .rst(f1862_rst), .rdata(f1862_rdata));
  assign f1862_clk = clk;
  assign f1862_rst = rst;
  // Bindings to f1862

  // f1864
  logic [0:0] f1864_wen;
  logic [31:0] f1864_wdata;
  logic [0:0] f1864_clk;
  logic [0:0] f1864_rst;
  logic [31:0] f1864_rdata;
  sr_buffer_32_1 f1864(.wen(f1864_wen), .wdata(f1864_wdata), .clk(f1864_clk), .rst(f1864_rst), .rdata(f1864_rdata));
  assign f1864_clk = clk;
  assign f1864_rst = rst;
  // Bindings to f1864

  // f1866
  logic [0:0] f1866_wen;
  logic [31:0] f1866_wdata;
  logic [0:0] f1866_clk;
  logic [0:0] f1866_rst;
  logic [31:0] f1866_rdata;
  sr_buffer_32_1 f1866(.wen(f1866_wen), .wdata(f1866_wdata), .clk(f1866_clk), .rst(f1866_rst), .rdata(f1866_rdata));
  assign f1866_clk = clk;
  assign f1866_rst = rst;
  // Bindings to f1866

  // f1868
  logic [0:0] f1868_wen;
  logic [31:0] f1868_wdata;
  logic [0:0] f1868_clk;
  logic [0:0] f1868_rst;
  logic [31:0] f1868_rdata;
  sr_buffer_32_1 f1868(.wen(f1868_wen), .wdata(f1868_wdata), .clk(f1868_clk), .rst(f1868_rst), .rdata(f1868_rdata));
  assign f1868_clk = clk;
  assign f1868_rst = rst;
  // Bindings to f1868

  // f1870
  logic [0:0] f1870_wen;
  logic [31:0] f1870_wdata;
  logic [0:0] f1870_clk;
  logic [0:0] f1870_rst;
  logic [31:0] f1870_rdata;
  sr_buffer_32_1 f1870(.wen(f1870_wen), .wdata(f1870_wdata), .clk(f1870_clk), .rst(f1870_rst), .rdata(f1870_rdata));
  assign f1870_clk = clk;
  assign f1870_rst = rst;
  // Bindings to f1870

  // f1872
  logic [0:0] f1872_wen;
  logic [31:0] f1872_wdata;
  logic [0:0] f1872_clk;
  logic [0:0] f1872_rst;
  logic [31:0] f1872_rdata;
  sr_buffer_32_1 f1872(.wen(f1872_wen), .wdata(f1872_wdata), .clk(f1872_clk), .rst(f1872_rst), .rdata(f1872_rdata));
  assign f1872_clk = clk;
  assign f1872_rst = rst;
  // Bindings to f1872

  // f1874
  logic [0:0] f1874_wen;
  logic [31:0] f1874_wdata;
  logic [0:0] f1874_clk;
  logic [0:0] f1874_rst;
  logic [31:0] f1874_rdata;
  sr_buffer_32_1 f1874(.wen(f1874_wen), .wdata(f1874_wdata), .clk(f1874_clk), .rst(f1874_rst), .rdata(f1874_rdata));
  assign f1874_clk = clk;
  assign f1874_rst = rst;
  // Bindings to f1874

  // f1876
  logic [0:0] f1876_wen;
  logic [31:0] f1876_wdata;
  logic [0:0] f1876_clk;
  logic [0:0] f1876_rst;
  logic [31:0] f1876_rdata;
  sr_buffer_32_1 f1876(.wen(f1876_wen), .wdata(f1876_wdata), .clk(f1876_clk), .rst(f1876_rst), .rdata(f1876_rdata));
  assign f1876_clk = clk;
  assign f1876_rst = rst;
  // Bindings to f1876

  // f1878
  logic [0:0] f1878_wen;
  logic [31:0] f1878_wdata;
  logic [0:0] f1878_clk;
  logic [0:0] f1878_rst;
  logic [31:0] f1878_rdata;
  sr_buffer_32_1 f1878(.wen(f1878_wen), .wdata(f1878_wdata), .clk(f1878_clk), .rst(f1878_rst), .rdata(f1878_rdata));
  assign f1878_clk = clk;
  assign f1878_rst = rst;
  // Bindings to f1878

  // f1880
  logic [0:0] f1880_wen;
  logic [31:0] f1880_wdata;
  logic [0:0] f1880_clk;
  logic [0:0] f1880_rst;
  logic [31:0] f1880_rdata;
  sr_buffer_32_1 f1880(.wen(f1880_wen), .wdata(f1880_wdata), .clk(f1880_clk), .rst(f1880_rst), .rdata(f1880_rdata));
  assign f1880_clk = clk;
  assign f1880_rst = rst;
  // Bindings to f1880

  // f1882
  logic [0:0] f1882_wen;
  logic [31:0] f1882_wdata;
  logic [0:0] f1882_clk;
  logic [0:0] f1882_rst;
  logic [31:0] f1882_rdata;
  sr_buffer_32_1 f1882(.wen(f1882_wen), .wdata(f1882_wdata), .clk(f1882_clk), .rst(f1882_rst), .rdata(f1882_rdata));
  assign f1882_clk = clk;
  assign f1882_rst = rst;
  // Bindings to f1882

  // f1884
  logic [0:0] f1884_wen;
  logic [31:0] f1884_wdata;
  logic [0:0] f1884_clk;
  logic [0:0] f1884_rst;
  logic [31:0] f1884_rdata;
  sr_buffer_32_1 f1884(.wen(f1884_wen), .wdata(f1884_wdata), .clk(f1884_clk), .rst(f1884_rst), .rdata(f1884_rdata));
  assign f1884_clk = clk;
  assign f1884_rst = rst;
  // Bindings to f1884

  // f1886
  logic [0:0] f1886_wen;
  logic [31:0] f1886_wdata;
  logic [0:0] f1886_clk;
  logic [0:0] f1886_rst;
  logic [31:0] f1886_rdata;
  sr_buffer_32_1 f1886(.wen(f1886_wen), .wdata(f1886_wdata), .clk(f1886_clk), .rst(f1886_rst), .rdata(f1886_rdata));
  assign f1886_clk = clk;
  assign f1886_rst = rst;
  // Bindings to f1886

  // f1888
  logic [0:0] f1888_wen;
  logic [31:0] f1888_wdata;
  logic [0:0] f1888_clk;
  logic [0:0] f1888_rst;
  logic [31:0] f1888_rdata;
  sr_buffer_32_1 f1888(.wen(f1888_wen), .wdata(f1888_wdata), .clk(f1888_clk), .rst(f1888_rst), .rdata(f1888_rdata));
  assign f1888_clk = clk;
  assign f1888_rst = rst;
  // Bindings to f1888

  // f1890
  logic [0:0] f1890_wen;
  logic [31:0] f1890_wdata;
  logic [0:0] f1890_clk;
  logic [0:0] f1890_rst;
  logic [31:0] f1890_rdata;
  sr_buffer_32_1 f1890(.wen(f1890_wen), .wdata(f1890_wdata), .clk(f1890_clk), .rst(f1890_rst), .rdata(f1890_rdata));
  assign f1890_clk = clk;
  assign f1890_rst = rst;
  // Bindings to f1890

  // f1892
  logic [0:0] f1892_wen;
  logic [31:0] f1892_wdata;
  logic [0:0] f1892_clk;
  logic [0:0] f1892_rst;
  logic [31:0] f1892_rdata;
  sr_buffer_32_1 f1892(.wen(f1892_wen), .wdata(f1892_wdata), .clk(f1892_clk), .rst(f1892_rst), .rdata(f1892_rdata));
  assign f1892_clk = clk;
  assign f1892_rst = rst;
  // Bindings to f1892

  // f1894
  logic [0:0] f1894_wen;
  logic [31:0] f1894_wdata;
  logic [0:0] f1894_clk;
  logic [0:0] f1894_rst;
  logic [31:0] f1894_rdata;
  sr_buffer_32_1 f1894(.wen(f1894_wen), .wdata(f1894_wdata), .clk(f1894_clk), .rst(f1894_rst), .rdata(f1894_rdata));
  assign f1894_clk = clk;
  assign f1894_rst = rst;
  // Bindings to f1894

  // f1896
  logic [0:0] f1896_wen;
  logic [31:0] f1896_wdata;
  logic [0:0] f1896_clk;
  logic [0:0] f1896_rst;
  logic [31:0] f1896_rdata;
  sr_buffer_32_1 f1896(.wen(f1896_wen), .wdata(f1896_wdata), .clk(f1896_clk), .rst(f1896_rst), .rdata(f1896_rdata));
  assign f1896_clk = clk;
  assign f1896_rst = rst;
  // Bindings to f1896

  // f1898
  logic [0:0] f1898_wen;
  logic [31:0] f1898_wdata;
  logic [0:0] f1898_clk;
  logic [0:0] f1898_rst;
  logic [31:0] f1898_rdata;
  sr_buffer_32_1 f1898(.wen(f1898_wen), .wdata(f1898_wdata), .clk(f1898_clk), .rst(f1898_rst), .rdata(f1898_rdata));
  assign f1898_clk = clk;
  assign f1898_rst = rst;
  // Bindings to f1898

  // f1900
  logic [0:0] f1900_wen;
  logic [31:0] f1900_wdata;
  logic [0:0] f1900_clk;
  logic [0:0] f1900_rst;
  logic [31:0] f1900_rdata;
  sr_buffer_32_1 f1900(.wen(f1900_wen), .wdata(f1900_wdata), .clk(f1900_clk), .rst(f1900_rst), .rdata(f1900_rdata));
  assign f1900_clk = clk;
  assign f1900_rst = rst;
  // Bindings to f1900

  // f1902
  logic [0:0] f1902_wen;
  logic [31:0] f1902_wdata;
  logic [0:0] f1902_clk;
  logic [0:0] f1902_rst;
  logic [31:0] f1902_rdata;
  sr_buffer_32_1 f1902(.wen(f1902_wen), .wdata(f1902_wdata), .clk(f1902_clk), .rst(f1902_rst), .rdata(f1902_rdata));
  assign f1902_clk = clk;
  assign f1902_rst = rst;
  // Bindings to f1902

  // f1904
  logic [0:0] f1904_wen;
  logic [31:0] f1904_wdata;
  logic [0:0] f1904_clk;
  logic [0:0] f1904_rst;
  logic [31:0] f1904_rdata;
  sr_buffer_32_1 f1904(.wen(f1904_wen), .wdata(f1904_wdata), .clk(f1904_clk), .rst(f1904_rst), .rdata(f1904_rdata));
  assign f1904_clk = clk;
  assign f1904_rst = rst;
  // Bindings to f1904

  // f1906
  logic [0:0] f1906_wen;
  logic [31:0] f1906_wdata;
  logic [0:0] f1906_clk;
  logic [0:0] f1906_rst;
  logic [31:0] f1906_rdata;
  sr_buffer_32_1 f1906(.wen(f1906_wen), .wdata(f1906_wdata), .clk(f1906_clk), .rst(f1906_rst), .rdata(f1906_rdata));
  assign f1906_clk = clk;
  assign f1906_rst = rst;
  // Bindings to f1906

  // f1908
  logic [0:0] f1908_wen;
  logic [31:0] f1908_wdata;
  logic [0:0] f1908_clk;
  logic [0:0] f1908_rst;
  logic [31:0] f1908_rdata;
  sr_buffer_32_1 f1908(.wen(f1908_wen), .wdata(f1908_wdata), .clk(f1908_clk), .rst(f1908_rst), .rdata(f1908_rdata));
  assign f1908_clk = clk;
  assign f1908_rst = rst;
  // Bindings to f1908

  // f1910
  logic [0:0] f1910_wen;
  logic [31:0] f1910_wdata;
  logic [0:0] f1910_clk;
  logic [0:0] f1910_rst;
  logic [31:0] f1910_rdata;
  sr_buffer_32_1 f1910(.wen(f1910_wen), .wdata(f1910_wdata), .clk(f1910_clk), .rst(f1910_rst), .rdata(f1910_rdata));
  assign f1910_clk = clk;
  assign f1910_rst = rst;
  // Bindings to f1910

  // f1912
  logic [0:0] f1912_wen;
  logic [31:0] f1912_wdata;
  logic [0:0] f1912_clk;
  logic [0:0] f1912_rst;
  logic [31:0] f1912_rdata;
  sr_buffer_32_1 f1912(.wen(f1912_wen), .wdata(f1912_wdata), .clk(f1912_clk), .rst(f1912_rst), .rdata(f1912_rdata));
  assign f1912_clk = clk;
  assign f1912_rst = rst;
  // Bindings to f1912

  // f1914
  logic [0:0] f1914_wen;
  logic [31:0] f1914_wdata;
  logic [0:0] f1914_clk;
  logic [0:0] f1914_rst;
  logic [31:0] f1914_rdata;
  sr_buffer_32_1 f1914(.wen(f1914_wen), .wdata(f1914_wdata), .clk(f1914_clk), .rst(f1914_rst), .rdata(f1914_rdata));
  assign f1914_clk = clk;
  assign f1914_rst = rst;
  // Bindings to f1914

  // f1916
  logic [0:0] f1916_wen;
  logic [31:0] f1916_wdata;
  logic [0:0] f1916_clk;
  logic [0:0] f1916_rst;
  logic [31:0] f1916_rdata;
  sr_buffer_32_1 f1916(.wen(f1916_wen), .wdata(f1916_wdata), .clk(f1916_clk), .rst(f1916_rst), .rdata(f1916_rdata));
  assign f1916_clk = clk;
  assign f1916_rst = rst;
  // Bindings to f1916

  // f1918
  logic [0:0] f1918_wen;
  logic [31:0] f1918_wdata;
  logic [0:0] f1918_clk;
  logic [0:0] f1918_rst;
  logic [31:0] f1918_rdata;
  sr_buffer_32_1 f1918(.wen(f1918_wen), .wdata(f1918_wdata), .clk(f1918_clk), .rst(f1918_rst), .rdata(f1918_rdata));
  assign f1918_clk = clk;
  assign f1918_rst = rst;
  // Bindings to f1918

  // f1920
  logic [0:0] f1920_wen;
  logic [31:0] f1920_wdata;
  logic [0:0] f1920_clk;
  logic [0:0] f1920_rst;
  logic [31:0] f1920_rdata;
  sr_buffer_32_1 f1920(.wen(f1920_wen), .wdata(f1920_wdata), .clk(f1920_clk), .rst(f1920_rst), .rdata(f1920_rdata));
  assign f1920_clk = clk;
  assign f1920_rst = rst;
  // Bindings to f1920

  // f1922
  logic [0:0] f1922_wen;
  logic [31:0] f1922_wdata;
  logic [0:0] f1922_clk;
  logic [0:0] f1922_rst;
  logic [31:0] f1922_rdata;
  sr_buffer_32_1 f1922(.wen(f1922_wen), .wdata(f1922_wdata), .clk(f1922_clk), .rst(f1922_rst), .rdata(f1922_rdata));
  assign f1922_clk = clk;
  assign f1922_rst = rst;
  // Bindings to f1922

  // f1924
  logic [0:0] f1924_wen;
  logic [31:0] f1924_wdata;
  logic [0:0] f1924_clk;
  logic [0:0] f1924_rst;
  logic [31:0] f1924_rdata;
  sr_buffer_32_1 f1924(.wen(f1924_wen), .wdata(f1924_wdata), .clk(f1924_clk), .rst(f1924_rst), .rdata(f1924_rdata));
  assign f1924_clk = clk;
  assign f1924_rst = rst;
  // Bindings to f1924

  // f1926
  logic [0:0] f1926_wen;
  logic [31:0] f1926_wdata;
  logic [0:0] f1926_clk;
  logic [0:0] f1926_rst;
  logic [31:0] f1926_rdata;
  sr_buffer_32_1 f1926(.wen(f1926_wen), .wdata(f1926_wdata), .clk(f1926_clk), .rst(f1926_rst), .rdata(f1926_rdata));
  assign f1926_clk = clk;
  assign f1926_rst = rst;
  // Bindings to f1926

  // f1928
  logic [0:0] f1928_wen;
  logic [31:0] f1928_wdata;
  logic [0:0] f1928_clk;
  logic [0:0] f1928_rst;
  logic [31:0] f1928_rdata;
  sr_buffer_32_1 f1928(.wen(f1928_wen), .wdata(f1928_wdata), .clk(f1928_clk), .rst(f1928_rst), .rdata(f1928_rdata));
  assign f1928_clk = clk;
  assign f1928_rst = rst;
  // Bindings to f1928

  // f1930
  logic [0:0] f1930_wen;
  logic [31:0] f1930_wdata;
  logic [0:0] f1930_clk;
  logic [0:0] f1930_rst;
  logic [31:0] f1930_rdata;
  sr_buffer_32_1 f1930(.wen(f1930_wen), .wdata(f1930_wdata), .clk(f1930_clk), .rst(f1930_rst), .rdata(f1930_rdata));
  assign f1930_clk = clk;
  assign f1930_rst = rst;
  // Bindings to f1930

  // f1932
  logic [0:0] f1932_wen;
  logic [31:0] f1932_wdata;
  logic [0:0] f1932_clk;
  logic [0:0] f1932_rst;
  logic [31:0] f1932_rdata;
  sr_buffer_32_1 f1932(.wen(f1932_wen), .wdata(f1932_wdata), .clk(f1932_clk), .rst(f1932_rst), .rdata(f1932_rdata));
  assign f1932_clk = clk;
  assign f1932_rst = rst;
  // Bindings to f1932

  // f1934
  logic [0:0] f1934_wen;
  logic [31:0] f1934_wdata;
  logic [0:0] f1934_clk;
  logic [0:0] f1934_rst;
  logic [31:0] f1934_rdata;
  sr_buffer_32_1 f1934(.wen(f1934_wen), .wdata(f1934_wdata), .clk(f1934_clk), .rst(f1934_rst), .rdata(f1934_rdata));
  assign f1934_clk = clk;
  assign f1934_rst = rst;
  // Bindings to f1934

  // f1936
  logic [0:0] f1936_wen;
  logic [31:0] f1936_wdata;
  logic [0:0] f1936_clk;
  logic [0:0] f1936_rst;
  logic [31:0] f1936_rdata;
  sr_buffer_32_1 f1936(.wen(f1936_wen), .wdata(f1936_wdata), .clk(f1936_clk), .rst(f1936_rst), .rdata(f1936_rdata));
  assign f1936_clk = clk;
  assign f1936_rst = rst;
  // Bindings to f1936

  // f1938
  logic [0:0] f1938_wen;
  logic [31:0] f1938_wdata;
  logic [0:0] f1938_clk;
  logic [0:0] f1938_rst;
  logic [31:0] f1938_rdata;
  sr_buffer_32_1 f1938(.wen(f1938_wen), .wdata(f1938_wdata), .clk(f1938_clk), .rst(f1938_rst), .rdata(f1938_rdata));
  assign f1938_clk = clk;
  assign f1938_rst = rst;
  // Bindings to f1938

  // f1940
  logic [0:0] f1940_wen;
  logic [31:0] f1940_wdata;
  logic [0:0] f1940_clk;
  logic [0:0] f1940_rst;
  logic [31:0] f1940_rdata;
  sr_buffer_32_1 f1940(.wen(f1940_wen), .wdata(f1940_wdata), .clk(f1940_clk), .rst(f1940_rst), .rdata(f1940_rdata));
  assign f1940_clk = clk;
  assign f1940_rst = rst;
  // Bindings to f1940

  // f1942
  logic [0:0] f1942_wen;
  logic [31:0] f1942_wdata;
  logic [0:0] f1942_clk;
  logic [0:0] f1942_rst;
  logic [31:0] f1942_rdata;
  sr_buffer_32_1 f1942(.wen(f1942_wen), .wdata(f1942_wdata), .clk(f1942_clk), .rst(f1942_rst), .rdata(f1942_rdata));
  assign f1942_clk = clk;
  assign f1942_rst = rst;
  // Bindings to f1942

  // f1944
  logic [0:0] f1944_wen;
  logic [31:0] f1944_wdata;
  logic [0:0] f1944_clk;
  logic [0:0] f1944_rst;
  logic [31:0] f1944_rdata;
  sr_buffer_32_1 f1944(.wen(f1944_wen), .wdata(f1944_wdata), .clk(f1944_clk), .rst(f1944_rst), .rdata(f1944_rdata));
  assign f1944_clk = clk;
  assign f1944_rst = rst;
  // Bindings to f1944

  // f1946
  logic [0:0] f1946_wen;
  logic [31:0] f1946_wdata;
  logic [0:0] f1946_clk;
  logic [0:0] f1946_rst;
  logic [31:0] f1946_rdata;
  sr_buffer_32_1 f1946(.wen(f1946_wen), .wdata(f1946_wdata), .clk(f1946_clk), .rst(f1946_rst), .rdata(f1946_rdata));
  assign f1946_clk = clk;
  assign f1946_rst = rst;
  // Bindings to f1946

  // f1948
  logic [0:0] f1948_wen;
  logic [31:0] f1948_wdata;
  logic [0:0] f1948_clk;
  logic [0:0] f1948_rst;
  logic [31:0] f1948_rdata;
  sr_buffer_32_1 f1948(.wen(f1948_wen), .wdata(f1948_wdata), .clk(f1948_clk), .rst(f1948_rst), .rdata(f1948_rdata));
  assign f1948_clk = clk;
  assign f1948_rst = rst;
  // Bindings to f1948

  // f1950
  logic [0:0] f1950_wen;
  logic [31:0] f1950_wdata;
  logic [0:0] f1950_clk;
  logic [0:0] f1950_rst;
  logic [31:0] f1950_rdata;
  sr_buffer_32_1 f1950(.wen(f1950_wen), .wdata(f1950_wdata), .clk(f1950_clk), .rst(f1950_rst), .rdata(f1950_rdata));
  assign f1950_clk = clk;
  assign f1950_rst = rst;
  // Bindings to f1950

  // f1952
  logic [0:0] f1952_wen;
  logic [31:0] f1952_wdata;
  logic [0:0] f1952_clk;
  logic [0:0] f1952_rst;
  logic [31:0] f1952_rdata;
  sr_buffer_32_1 f1952(.wen(f1952_wen), .wdata(f1952_wdata), .clk(f1952_clk), .rst(f1952_rst), .rdata(f1952_rdata));
  assign f1952_clk = clk;
  assign f1952_rst = rst;
  // Bindings to f1952

  // f1954
  logic [0:0] f1954_wen;
  logic [31:0] f1954_wdata;
  logic [0:0] f1954_clk;
  logic [0:0] f1954_rst;
  logic [31:0] f1954_rdata;
  sr_buffer_32_1 f1954(.wen(f1954_wen), .wdata(f1954_wdata), .clk(f1954_clk), .rst(f1954_rst), .rdata(f1954_rdata));
  assign f1954_clk = clk;
  assign f1954_rst = rst;
  // Bindings to f1954

  // f1956
  logic [0:0] f1956_wen;
  logic [31:0] f1956_wdata;
  logic [0:0] f1956_clk;
  logic [0:0] f1956_rst;
  logic [31:0] f1956_rdata;
  sr_buffer_32_1 f1956(.wen(f1956_wen), .wdata(f1956_wdata), .clk(f1956_clk), .rst(f1956_rst), .rdata(f1956_rdata));
  assign f1956_clk = clk;
  assign f1956_rst = rst;
  // Bindings to f1956

  // f1958
  logic [0:0] f1958_wen;
  logic [31:0] f1958_wdata;
  logic [0:0] f1958_clk;
  logic [0:0] f1958_rst;
  logic [31:0] f1958_rdata;
  sr_buffer_32_1 f1958(.wen(f1958_wen), .wdata(f1958_wdata), .clk(f1958_clk), .rst(f1958_rst), .rdata(f1958_rdata));
  assign f1958_clk = clk;
  assign f1958_rst = rst;
  // Bindings to f1958

  // f1960
  logic [0:0] f1960_wen;
  logic [31:0] f1960_wdata;
  logic [0:0] f1960_clk;
  logic [0:0] f1960_rst;
  logic [31:0] f1960_rdata;
  sr_buffer_32_1 f1960(.wen(f1960_wen), .wdata(f1960_wdata), .clk(f1960_clk), .rst(f1960_rst), .rdata(f1960_rdata));
  assign f1960_clk = clk;
  assign f1960_rst = rst;
  // Bindings to f1960

  // f1962
  logic [0:0] f1962_wen;
  logic [31:0] f1962_wdata;
  logic [0:0] f1962_clk;
  logic [0:0] f1962_rst;
  logic [31:0] f1962_rdata;
  sr_buffer_32_1 f1962(.wen(f1962_wen), .wdata(f1962_wdata), .clk(f1962_clk), .rst(f1962_rst), .rdata(f1962_rdata));
  assign f1962_clk = clk;
  assign f1962_rst = rst;
  // Bindings to f1962

  // f1964
  logic [0:0] f1964_wen;
  logic [31:0] f1964_wdata;
  logic [0:0] f1964_clk;
  logic [0:0] f1964_rst;
  logic [31:0] f1964_rdata;
  sr_buffer_32_1 f1964(.wen(f1964_wen), .wdata(f1964_wdata), .clk(f1964_clk), .rst(f1964_rst), .rdata(f1964_rdata));
  assign f1964_clk = clk;
  assign f1964_rst = rst;
  // Bindings to f1964

  // f1966
  logic [0:0] f1966_wen;
  logic [31:0] f1966_wdata;
  logic [0:0] f1966_clk;
  logic [0:0] f1966_rst;
  logic [31:0] f1966_rdata;
  sr_buffer_32_1 f1966(.wen(f1966_wen), .wdata(f1966_wdata), .clk(f1966_clk), .rst(f1966_rst), .rdata(f1966_rdata));
  assign f1966_clk = clk;
  assign f1966_rst = rst;
  // Bindings to f1966

  // f1968
  logic [0:0] f1968_wen;
  logic [31:0] f1968_wdata;
  logic [0:0] f1968_clk;
  logic [0:0] f1968_rst;
  logic [31:0] f1968_rdata;
  sr_buffer_32_1 f1968(.wen(f1968_wen), .wdata(f1968_wdata), .clk(f1968_clk), .rst(f1968_rst), .rdata(f1968_rdata));
  assign f1968_clk = clk;
  assign f1968_rst = rst;
  // Bindings to f1968

  // f1970
  logic [0:0] f1970_wen;
  logic [31:0] f1970_wdata;
  logic [0:0] f1970_clk;
  logic [0:0] f1970_rst;
  logic [31:0] f1970_rdata;
  sr_buffer_32_1 f1970(.wen(f1970_wen), .wdata(f1970_wdata), .clk(f1970_clk), .rst(f1970_rst), .rdata(f1970_rdata));
  assign f1970_clk = clk;
  assign f1970_rst = rst;
  // Bindings to f1970

  // f1972
  logic [0:0] f1972_wen;
  logic [31:0] f1972_wdata;
  logic [0:0] f1972_clk;
  logic [0:0] f1972_rst;
  logic [31:0] f1972_rdata;
  sr_buffer_32_1 f1972(.wen(f1972_wen), .wdata(f1972_wdata), .clk(f1972_clk), .rst(f1972_rst), .rdata(f1972_rdata));
  assign f1972_clk = clk;
  assign f1972_rst = rst;
  // Bindings to f1972

  // f1974
  logic [0:0] f1974_wen;
  logic [31:0] f1974_wdata;
  logic [0:0] f1974_clk;
  logic [0:0] f1974_rst;
  logic [31:0] f1974_rdata;
  sr_buffer_32_1 f1974(.wen(f1974_wen), .wdata(f1974_wdata), .clk(f1974_clk), .rst(f1974_rst), .rdata(f1974_rdata));
  assign f1974_clk = clk;
  assign f1974_rst = rst;
  // Bindings to f1974

  // f1976
  logic [0:0] f1976_wen;
  logic [31:0] f1976_wdata;
  logic [0:0] f1976_clk;
  logic [0:0] f1976_rst;
  logic [31:0] f1976_rdata;
  sr_buffer_32_1 f1976(.wen(f1976_wen), .wdata(f1976_wdata), .clk(f1976_clk), .rst(f1976_rst), .rdata(f1976_rdata));
  assign f1976_clk = clk;
  assign f1976_rst = rst;
  // Bindings to f1976

  // f1978
  logic [0:0] f1978_wen;
  logic [31:0] f1978_wdata;
  logic [0:0] f1978_clk;
  logic [0:0] f1978_rst;
  logic [31:0] f1978_rdata;
  sr_buffer_32_1 f1978(.wen(f1978_wen), .wdata(f1978_wdata), .clk(f1978_clk), .rst(f1978_rst), .rdata(f1978_rdata));
  assign f1978_clk = clk;
  assign f1978_rst = rst;
  // Bindings to f1978

  // f1980
  logic [0:0] f1980_wen;
  logic [31:0] f1980_wdata;
  logic [0:0] f1980_clk;
  logic [0:0] f1980_rst;
  logic [31:0] f1980_rdata;
  sr_buffer_32_1 f1980(.wen(f1980_wen), .wdata(f1980_wdata), .clk(f1980_clk), .rst(f1980_rst), .rdata(f1980_rdata));
  assign f1980_clk = clk;
  assign f1980_rst = rst;
  // Bindings to f1980

  // f1982
  logic [0:0] f1982_wen;
  logic [31:0] f1982_wdata;
  logic [0:0] f1982_clk;
  logic [0:0] f1982_rst;
  logic [31:0] f1982_rdata;
  sr_buffer_32_1 f1982(.wen(f1982_wen), .wdata(f1982_wdata), .clk(f1982_clk), .rst(f1982_rst), .rdata(f1982_rdata));
  assign f1982_clk = clk;
  assign f1982_rst = rst;
  // Bindings to f1982

  // f1984
  logic [0:0] f1984_wen;
  logic [31:0] f1984_wdata;
  logic [0:0] f1984_clk;
  logic [0:0] f1984_rst;
  logic [31:0] f1984_rdata;
  sr_buffer_32_1 f1984(.wen(f1984_wen), .wdata(f1984_wdata), .clk(f1984_clk), .rst(f1984_rst), .rdata(f1984_rdata));
  assign f1984_clk = clk;
  assign f1984_rst = rst;
  // Bindings to f1984

  // f1986
  logic [0:0] f1986_wen;
  logic [31:0] f1986_wdata;
  logic [0:0] f1986_clk;
  logic [0:0] f1986_rst;
  logic [31:0] f1986_rdata;
  sr_buffer_32_1 f1986(.wen(f1986_wen), .wdata(f1986_wdata), .clk(f1986_clk), .rst(f1986_rst), .rdata(f1986_rdata));
  assign f1986_clk = clk;
  assign f1986_rst = rst;
  // Bindings to f1986

  // f1988
  logic [0:0] f1988_wen;
  logic [31:0] f1988_wdata;
  logic [0:0] f1988_clk;
  logic [0:0] f1988_rst;
  logic [31:0] f1988_rdata;
  sr_buffer_32_1 f1988(.wen(f1988_wen), .wdata(f1988_wdata), .clk(f1988_clk), .rst(f1988_rst), .rdata(f1988_rdata));
  assign f1988_clk = clk;
  assign f1988_rst = rst;
  // Bindings to f1988

  // f1990
  logic [0:0] f1990_wen;
  logic [31:0] f1990_wdata;
  logic [0:0] f1990_clk;
  logic [0:0] f1990_rst;
  logic [31:0] f1990_rdata;
  sr_buffer_32_1 f1990(.wen(f1990_wen), .wdata(f1990_wdata), .clk(f1990_clk), .rst(f1990_rst), .rdata(f1990_rdata));
  assign f1990_clk = clk;
  assign f1990_rst = rst;
  // Bindings to f1990

  // f1992
  logic [0:0] f1992_wen;
  logic [31:0] f1992_wdata;
  logic [0:0] f1992_clk;
  logic [0:0] f1992_rst;
  logic [31:0] f1992_rdata;
  sr_buffer_32_1 f1992(.wen(f1992_wen), .wdata(f1992_wdata), .clk(f1992_clk), .rst(f1992_rst), .rdata(f1992_rdata));
  assign f1992_clk = clk;
  assign f1992_rst = rst;
  // Bindings to f1992

  // f1994
  logic [0:0] f1994_wen;
  logic [31:0] f1994_wdata;
  logic [0:0] f1994_clk;
  logic [0:0] f1994_rst;
  logic [31:0] f1994_rdata;
  sr_buffer_32_1 f1994(.wen(f1994_wen), .wdata(f1994_wdata), .clk(f1994_clk), .rst(f1994_rst), .rdata(f1994_rdata));
  assign f1994_clk = clk;
  assign f1994_rst = rst;
  // Bindings to f1994

  // f1996
  logic [0:0] f1996_wen;
  logic [31:0] f1996_wdata;
  logic [0:0] f1996_clk;
  logic [0:0] f1996_rst;
  logic [31:0] f1996_rdata;
  sr_buffer_32_1 f1996(.wen(f1996_wen), .wdata(f1996_wdata), .clk(f1996_clk), .rst(f1996_rst), .rdata(f1996_rdata));
  assign f1996_clk = clk;
  assign f1996_rst = rst;
  // Bindings to f1996

  // f1998
  logic [0:0] f1998_wen;
  logic [31:0] f1998_wdata;
  logic [0:0] f1998_clk;
  logic [0:0] f1998_rst;
  logic [31:0] f1998_rdata;
  sr_buffer_32_1 f1998(.wen(f1998_wen), .wdata(f1998_wdata), .clk(f1998_clk), .rst(f1998_rst), .rdata(f1998_rdata));
  assign f1998_clk = clk;
  assign f1998_rst = rst;
  // Bindings to f1998

  // f2000
  logic [0:0] f2000_wen;
  logic [31:0] f2000_wdata;
  logic [0:0] f2000_clk;
  logic [0:0] f2000_rst;
  logic [31:0] f2000_rdata;
  sr_buffer_32_1 f2000(.wen(f2000_wen), .wdata(f2000_wdata), .clk(f2000_clk), .rst(f2000_rst), .rdata(f2000_rdata));
  assign f2000_clk = clk;
  assign f2000_rst = rst;
  // Bindings to f2000

  // f2002
  logic [0:0] f2002_wen;
  logic [31:0] f2002_wdata;
  logic [0:0] f2002_clk;
  logic [0:0] f2002_rst;
  logic [31:0] f2002_rdata;
  sr_buffer_32_1 f2002(.wen(f2002_wen), .wdata(f2002_wdata), .clk(f2002_clk), .rst(f2002_rst), .rdata(f2002_rdata));
  assign f2002_clk = clk;
  assign f2002_rst = rst;
  // Bindings to f2002

  // f2004
  logic [0:0] f2004_wen;
  logic [31:0] f2004_wdata;
  logic [0:0] f2004_clk;
  logic [0:0] f2004_rst;
  logic [31:0] f2004_rdata;
  sr_buffer_32_1 f2004(.wen(f2004_wen), .wdata(f2004_wdata), .clk(f2004_clk), .rst(f2004_rst), .rdata(f2004_rdata));
  assign f2004_clk = clk;
  assign f2004_rst = rst;
  // Bindings to f2004

  // f2006
  logic [0:0] f2006_wen;
  logic [31:0] f2006_wdata;
  logic [0:0] f2006_clk;
  logic [0:0] f2006_rst;
  logic [31:0] f2006_rdata;
  sr_buffer_32_1 f2006(.wen(f2006_wen), .wdata(f2006_wdata), .clk(f2006_clk), .rst(f2006_rst), .rdata(f2006_rdata));
  assign f2006_clk = clk;
  assign f2006_rst = rst;
  // Bindings to f2006

  // f2008
  logic [0:0] f2008_wen;
  logic [31:0] f2008_wdata;
  logic [0:0] f2008_clk;
  logic [0:0] f2008_rst;
  logic [31:0] f2008_rdata;
  sr_buffer_32_1 f2008(.wen(f2008_wen), .wdata(f2008_wdata), .clk(f2008_clk), .rst(f2008_rst), .rdata(f2008_rdata));
  assign f2008_clk = clk;
  assign f2008_rst = rst;
  // Bindings to f2008

  // f2010
  logic [0:0] f2010_wen;
  logic [31:0] f2010_wdata;
  logic [0:0] f2010_clk;
  logic [0:0] f2010_rst;
  logic [31:0] f2010_rdata;
  sr_buffer_32_1 f2010(.wen(f2010_wen), .wdata(f2010_wdata), .clk(f2010_clk), .rst(f2010_rst), .rdata(f2010_rdata));
  assign f2010_clk = clk;
  assign f2010_rst = rst;
  // Bindings to f2010

  // f2012
  logic [0:0] f2012_wen;
  logic [31:0] f2012_wdata;
  logic [0:0] f2012_clk;
  logic [0:0] f2012_rst;
  logic [31:0] f2012_rdata;
  sr_buffer_32_1 f2012(.wen(f2012_wen), .wdata(f2012_wdata), .clk(f2012_clk), .rst(f2012_rst), .rdata(f2012_rdata));
  assign f2012_clk = clk;
  assign f2012_rst = rst;
  // Bindings to f2012

  // f2014
  logic [0:0] f2014_wen;
  logic [31:0] f2014_wdata;
  logic [0:0] f2014_clk;
  logic [0:0] f2014_rst;
  logic [31:0] f2014_rdata;
  sr_buffer_32_1 f2014(.wen(f2014_wen), .wdata(f2014_wdata), .clk(f2014_clk), .rst(f2014_rst), .rdata(f2014_rdata));
  assign f2014_clk = clk;
  assign f2014_rst = rst;
  // Bindings to f2014

  // f2016
  logic [0:0] f2016_wen;
  logic [31:0] f2016_wdata;
  logic [0:0] f2016_clk;
  logic [0:0] f2016_rst;
  logic [31:0] f2016_rdata;
  sr_buffer_32_1 f2016(.wen(f2016_wen), .wdata(f2016_wdata), .clk(f2016_clk), .rst(f2016_rst), .rdata(f2016_rdata));
  assign f2016_clk = clk;
  assign f2016_rst = rst;
  // Bindings to f2016

  // f2018
  logic [0:0] f2018_wen;
  logic [31:0] f2018_wdata;
  logic [0:0] f2018_clk;
  logic [0:0] f2018_rst;
  logic [31:0] f2018_rdata;
  sr_buffer_32_1 f2018(.wen(f2018_wen), .wdata(f2018_wdata), .clk(f2018_clk), .rst(f2018_rst), .rdata(f2018_rdata));
  assign f2018_clk = clk;
  assign f2018_rst = rst;
  // Bindings to f2018

  // f2020
  logic [0:0] f2020_wen;
  logic [31:0] f2020_wdata;
  logic [0:0] f2020_clk;
  logic [0:0] f2020_rst;
  logic [31:0] f2020_rdata;
  sr_buffer_32_1 f2020(.wen(f2020_wen), .wdata(f2020_wdata), .clk(f2020_clk), .rst(f2020_rst), .rdata(f2020_rdata));
  assign f2020_clk = clk;
  assign f2020_rst = rst;
  // Bindings to f2020

  // f2022
  logic [0:0] f2022_wen;
  logic [31:0] f2022_wdata;
  logic [0:0] f2022_clk;
  logic [0:0] f2022_rst;
  logic [31:0] f2022_rdata;
  sr_buffer_32_1 f2022(.wen(f2022_wen), .wdata(f2022_wdata), .clk(f2022_clk), .rst(f2022_rst), .rdata(f2022_rdata));
  assign f2022_clk = clk;
  assign f2022_rst = rst;
  // Bindings to f2022

  // f2024
  logic [0:0] f2024_wen;
  logic [31:0] f2024_wdata;
  logic [0:0] f2024_clk;
  logic [0:0] f2024_rst;
  logic [31:0] f2024_rdata;
  sr_buffer_32_1 f2024(.wen(f2024_wen), .wdata(f2024_wdata), .clk(f2024_clk), .rst(f2024_rst), .rdata(f2024_rdata));
  assign f2024_clk = clk;
  assign f2024_rst = rst;
  // Bindings to f2024

  // f2026
  logic [0:0] f2026_wen;
  logic [31:0] f2026_wdata;
  logic [0:0] f2026_clk;
  logic [0:0] f2026_rst;
  logic [31:0] f2026_rdata;
  sr_buffer_32_1 f2026(.wen(f2026_wen), .wdata(f2026_wdata), .clk(f2026_clk), .rst(f2026_rst), .rdata(f2026_rdata));
  assign f2026_clk = clk;
  assign f2026_rst = rst;
  // Bindings to f2026

  // f2028
  logic [0:0] f2028_wen;
  logic [31:0] f2028_wdata;
  logic [0:0] f2028_clk;
  logic [0:0] f2028_rst;
  logic [31:0] f2028_rdata;
  sr_buffer_32_1 f2028(.wen(f2028_wen), .wdata(f2028_wdata), .clk(f2028_clk), .rst(f2028_rst), .rdata(f2028_rdata));
  assign f2028_clk = clk;
  assign f2028_rst = rst;
  // Bindings to f2028

  // f2030
  logic [0:0] f2030_wen;
  logic [31:0] f2030_wdata;
  logic [0:0] f2030_clk;
  logic [0:0] f2030_rst;
  logic [31:0] f2030_rdata;
  sr_buffer_32_1 f2030(.wen(f2030_wen), .wdata(f2030_wdata), .clk(f2030_clk), .rst(f2030_rst), .rdata(f2030_rdata));
  assign f2030_clk = clk;
  assign f2030_rst = rst;
  // Bindings to f2030

  // f2032
  logic [0:0] f2032_wen;
  logic [31:0] f2032_wdata;
  logic [0:0] f2032_clk;
  logic [0:0] f2032_rst;
  logic [31:0] f2032_rdata;
  sr_buffer_32_1 f2032(.wen(f2032_wen), .wdata(f2032_wdata), .clk(f2032_clk), .rst(f2032_rst), .rdata(f2032_rdata));
  assign f2032_clk = clk;
  assign f2032_rst = rst;
  // Bindings to f2032

  // f2034
  logic [0:0] f2034_wen;
  logic [31:0] f2034_wdata;
  logic [0:0] f2034_clk;
  logic [0:0] f2034_rst;
  logic [31:0] f2034_rdata;
  sr_buffer_32_1 f2034(.wen(f2034_wen), .wdata(f2034_wdata), .clk(f2034_clk), .rst(f2034_rst), .rdata(f2034_rdata));
  assign f2034_clk = clk;
  assign f2034_rst = rst;
  // Bindings to f2034

  // f2036
  logic [0:0] f2036_wen;
  logic [31:0] f2036_wdata;
  logic [0:0] f2036_clk;
  logic [0:0] f2036_rst;
  logic [31:0] f2036_rdata;
  sr_buffer_32_1 f2036(.wen(f2036_wen), .wdata(f2036_wdata), .clk(f2036_clk), .rst(f2036_rst), .rdata(f2036_rdata));
  assign f2036_clk = clk;
  assign f2036_rst = rst;
  // Bindings to f2036

  // f2038
  logic [0:0] f2038_wen;
  logic [31:0] f2038_wdata;
  logic [0:0] f2038_clk;
  logic [0:0] f2038_rst;
  logic [31:0] f2038_rdata;
  sr_buffer_32_1 f2038(.wen(f2038_wen), .wdata(f2038_wdata), .clk(f2038_clk), .rst(f2038_rst), .rdata(f2038_rdata));
  assign f2038_clk = clk;
  assign f2038_rst = rst;
  // Bindings to f2038

  // f2040
  logic [0:0] f2040_wen;
  logic [31:0] f2040_wdata;
  logic [0:0] f2040_clk;
  logic [0:0] f2040_rst;
  logic [31:0] f2040_rdata;
  sr_buffer_32_1 f2040(.wen(f2040_wen), .wdata(f2040_wdata), .clk(f2040_clk), .rst(f2040_rst), .rdata(f2040_rdata));
  assign f2040_clk = clk;
  assign f2040_rst = rst;
  // Bindings to f2040

  // f2042
  logic [0:0] f2042_wen;
  logic [31:0] f2042_wdata;
  logic [0:0] f2042_clk;
  logic [0:0] f2042_rst;
  logic [31:0] f2042_rdata;
  sr_buffer_32_1 f2042(.wen(f2042_wen), .wdata(f2042_wdata), .clk(f2042_clk), .rst(f2042_rst), .rdata(f2042_rdata));
  assign f2042_clk = clk;
  assign f2042_rst = rst;
  // Bindings to f2042

  // f2044
  logic [0:0] f2044_wen;
  logic [31:0] f2044_wdata;
  logic [0:0] f2044_clk;
  logic [0:0] f2044_rst;
  logic [31:0] f2044_rdata;
  sr_buffer_32_1 f2044(.wen(f2044_wen), .wdata(f2044_wdata), .clk(f2044_clk), .rst(f2044_rst), .rdata(f2044_rdata));
  assign f2044_clk = clk;
  assign f2044_rst = rst;
  // Bindings to f2044

  // f2046
  logic [0:0] f2046_wen;
  logic [31:0] f2046_wdata;
  logic [0:0] f2046_clk;
  logic [0:0] f2046_rst;
  logic [31:0] f2046_rdata;
  sr_buffer_32_1 f2046(.wen(f2046_wen), .wdata(f2046_wdata), .clk(f2046_clk), .rst(f2046_rst), .rdata(f2046_rdata));
  assign f2046_clk = clk;
  assign f2046_rst = rst;
  // Bindings to f2046

  // f2048
  logic [0:0] f2048_wen;
  logic [31:0] f2048_wdata;
  logic [0:0] f2048_clk;
  logic [0:0] f2048_rst;
  logic [31:0] f2048_rdata;
  sr_buffer_32_1 f2048(.wen(f2048_wen), .wdata(f2048_wdata), .clk(f2048_clk), .rst(f2048_rst), .rdata(f2048_rdata));
  assign f2048_clk = clk;
  assign f2048_rst = rst;
  // Bindings to f2048

  // f2050
  logic [0:0] f2050_wen;
  logic [31:0] f2050_wdata;
  logic [0:0] f2050_clk;
  logic [0:0] f2050_rst;
  logic [31:0] f2050_rdata;
  sr_buffer_32_1 f2050(.wen(f2050_wen), .wdata(f2050_wdata), .clk(f2050_clk), .rst(f2050_rst), .rdata(f2050_rdata));
  assign f2050_clk = clk;
  assign f2050_rst = rst;
  // Bindings to f2050

  // f2052
  logic [0:0] f2052_wen;
  logic [31:0] f2052_wdata;
  logic [0:0] f2052_clk;
  logic [0:0] f2052_rst;
  logic [31:0] f2052_rdata;
  sr_buffer_32_1 f2052(.wen(f2052_wen), .wdata(f2052_wdata), .clk(f2052_clk), .rst(f2052_rst), .rdata(f2052_rdata));
  assign f2052_clk = clk;
  assign f2052_rst = rst;
  // Bindings to f2052

  // f2054
  logic [0:0] f2054_wen;
  logic [31:0] f2054_wdata;
  logic [0:0] f2054_clk;
  logic [0:0] f2054_rst;
  logic [31:0] f2054_rdata;
  sr_buffer_32_1 f2054(.wen(f2054_wen), .wdata(f2054_wdata), .clk(f2054_clk), .rst(f2054_rst), .rdata(f2054_rdata));
  assign f2054_clk = clk;
  assign f2054_rst = rst;
  // Bindings to f2054

  // f2056
  logic [0:0] f2056_wen;
  logic [31:0] f2056_wdata;
  logic [0:0] f2056_clk;
  logic [0:0] f2056_rst;
  logic [31:0] f2056_rdata;
  sr_buffer_32_1 f2056(.wen(f2056_wen), .wdata(f2056_wdata), .clk(f2056_clk), .rst(f2056_rst), .rdata(f2056_rdata));
  assign f2056_clk = clk;
  assign f2056_rst = rst;
  // Bindings to f2056

  // f2058
  logic [0:0] f2058_wen;
  logic [31:0] f2058_wdata;
  logic [0:0] f2058_clk;
  logic [0:0] f2058_rst;
  logic [31:0] f2058_rdata;
  sr_buffer_32_1 f2058(.wen(f2058_wen), .wdata(f2058_wdata), .clk(f2058_clk), .rst(f2058_rst), .rdata(f2058_rdata));
  assign f2058_clk = clk;
  assign f2058_rst = rst;
  // Bindings to f2058

  // f2060
  logic [0:0] f2060_wen;
  logic [31:0] f2060_wdata;
  logic [0:0] f2060_clk;
  logic [0:0] f2060_rst;
  logic [31:0] f2060_rdata;
  sr_buffer_32_1 f2060(.wen(f2060_wen), .wdata(f2060_wdata), .clk(f2060_clk), .rst(f2060_rst), .rdata(f2060_rdata));
  assign f2060_clk = clk;
  assign f2060_rst = rst;
  // Bindings to f2060

  // f2062
  logic [0:0] f2062_wen;
  logic [31:0] f2062_wdata;
  logic [0:0] f2062_clk;
  logic [0:0] f2062_rst;
  logic [31:0] f2062_rdata;
  sr_buffer_32_1 f2062(.wen(f2062_wen), .wdata(f2062_wdata), .clk(f2062_clk), .rst(f2062_rst), .rdata(f2062_rdata));
  assign f2062_clk = clk;
  assign f2062_rst = rst;
  // Bindings to f2062

  // f2064
  logic [0:0] f2064_wen;
  logic [31:0] f2064_wdata;
  logic [0:0] f2064_clk;
  logic [0:0] f2064_rst;
  logic [31:0] f2064_rdata;
  sr_buffer_32_1 f2064(.wen(f2064_wen), .wdata(f2064_wdata), .clk(f2064_clk), .rst(f2064_rst), .rdata(f2064_rdata));
  assign f2064_clk = clk;
  assign f2064_rst = rst;
  // Bindings to f2064

  // f2066
  logic [0:0] f2066_wen;
  logic [31:0] f2066_wdata;
  logic [0:0] f2066_clk;
  logic [0:0] f2066_rst;
  logic [31:0] f2066_rdata;
  sr_buffer_32_1 f2066(.wen(f2066_wen), .wdata(f2066_wdata), .clk(f2066_clk), .rst(f2066_rst), .rdata(f2066_rdata));
  assign f2066_clk = clk;
  assign f2066_rst = rst;
  // Bindings to f2066

  // f2068
  logic [0:0] f2068_wen;
  logic [31:0] f2068_wdata;
  logic [0:0] f2068_clk;
  logic [0:0] f2068_rst;
  logic [31:0] f2068_rdata;
  sr_buffer_32_1 f2068(.wen(f2068_wen), .wdata(f2068_wdata), .clk(f2068_clk), .rst(f2068_rst), .rdata(f2068_rdata));
  assign f2068_clk = clk;
  assign f2068_rst = rst;
  // Bindings to f2068

  // f2070
  logic [0:0] f2070_wen;
  logic [31:0] f2070_wdata;
  logic [0:0] f2070_clk;
  logic [0:0] f2070_rst;
  logic [31:0] f2070_rdata;
  sr_buffer_32_1 f2070(.wen(f2070_wen), .wdata(f2070_wdata), .clk(f2070_clk), .rst(f2070_rst), .rdata(f2070_rdata));
  assign f2070_clk = clk;
  assign f2070_rst = rst;
  // Bindings to f2070

  // f2072
  logic [0:0] f2072_wen;
  logic [31:0] f2072_wdata;
  logic [0:0] f2072_clk;
  logic [0:0] f2072_rst;
  logic [31:0] f2072_rdata;
  sr_buffer_32_1 f2072(.wen(f2072_wen), .wdata(f2072_wdata), .clk(f2072_clk), .rst(f2072_rst), .rdata(f2072_rdata));
  assign f2072_clk = clk;
  assign f2072_rst = rst;
  // Bindings to f2072

  // f2074
  logic [0:0] f2074_wen;
  logic [31:0] f2074_wdata;
  logic [0:0] f2074_clk;
  logic [0:0] f2074_rst;
  logic [31:0] f2074_rdata;
  sr_buffer_32_1 f2074(.wen(f2074_wen), .wdata(f2074_wdata), .clk(f2074_clk), .rst(f2074_rst), .rdata(f2074_rdata));
  assign f2074_clk = clk;
  assign f2074_rst = rst;
  // Bindings to f2074

  // f2076
  logic [0:0] f2076_wen;
  logic [31:0] f2076_wdata;
  logic [0:0] f2076_clk;
  logic [0:0] f2076_rst;
  logic [31:0] f2076_rdata;
  sr_buffer_32_1 f2076(.wen(f2076_wen), .wdata(f2076_wdata), .clk(f2076_clk), .rst(f2076_rst), .rdata(f2076_rdata));
  assign f2076_clk = clk;
  assign f2076_rst = rst;
  // Bindings to f2076

  // f2078
  logic [0:0] f2078_wen;
  logic [31:0] f2078_wdata;
  logic [0:0] f2078_clk;
  logic [0:0] f2078_rst;
  logic [31:0] f2078_rdata;
  sr_buffer_32_1 f2078(.wen(f2078_wen), .wdata(f2078_wdata), .clk(f2078_clk), .rst(f2078_rst), .rdata(f2078_rdata));
  assign f2078_clk = clk;
  assign f2078_rst = rst;
  // Bindings to f2078

  // f2080
  logic [0:0] f2080_wen;
  logic [31:0] f2080_wdata;
  logic [0:0] f2080_clk;
  logic [0:0] f2080_rst;
  logic [31:0] f2080_rdata;
  sr_buffer_32_1 f2080(.wen(f2080_wen), .wdata(f2080_wdata), .clk(f2080_clk), .rst(f2080_rst), .rdata(f2080_rdata));
  assign f2080_clk = clk;
  assign f2080_rst = rst;
  // Bindings to f2080

  // f2082
  logic [0:0] f2082_wen;
  logic [31:0] f2082_wdata;
  logic [0:0] f2082_clk;
  logic [0:0] f2082_rst;
  logic [31:0] f2082_rdata;
  sr_buffer_32_1 f2082(.wen(f2082_wen), .wdata(f2082_wdata), .clk(f2082_clk), .rst(f2082_rst), .rdata(f2082_rdata));
  assign f2082_clk = clk;
  assign f2082_rst = rst;
  // Bindings to f2082

  // f2084
  logic [0:0] f2084_wen;
  logic [31:0] f2084_wdata;
  logic [0:0] f2084_clk;
  logic [0:0] f2084_rst;
  logic [31:0] f2084_rdata;
  sr_buffer_32_1 f2084(.wen(f2084_wen), .wdata(f2084_wdata), .clk(f2084_clk), .rst(f2084_rst), .rdata(f2084_rdata));
  assign f2084_clk = clk;
  assign f2084_rst = rst;
  // Bindings to f2084

  // f2086
  logic [0:0] f2086_wen;
  logic [31:0] f2086_wdata;
  logic [0:0] f2086_clk;
  logic [0:0] f2086_rst;
  logic [31:0] f2086_rdata;
  sr_buffer_32_1 f2086(.wen(f2086_wen), .wdata(f2086_wdata), .clk(f2086_clk), .rst(f2086_rst), .rdata(f2086_rdata));
  assign f2086_clk = clk;
  assign f2086_rst = rst;
  // Bindings to f2086

  // f2088
  logic [0:0] f2088_wen;
  logic [31:0] f2088_wdata;
  logic [0:0] f2088_clk;
  logic [0:0] f2088_rst;
  logic [31:0] f2088_rdata;
  sr_buffer_32_1 f2088(.wen(f2088_wen), .wdata(f2088_wdata), .clk(f2088_clk), .rst(f2088_rst), .rdata(f2088_rdata));
  assign f2088_clk = clk;
  assign f2088_rst = rst;
  // Bindings to f2088

  // f2090
  logic [0:0] f2090_wen;
  logic [31:0] f2090_wdata;
  logic [0:0] f2090_clk;
  logic [0:0] f2090_rst;
  logic [31:0] f2090_rdata;
  sr_buffer_32_1 f2090(.wen(f2090_wen), .wdata(f2090_wdata), .clk(f2090_clk), .rst(f2090_rst), .rdata(f2090_rdata));
  assign f2090_clk = clk;
  assign f2090_rst = rst;
  // Bindings to f2090

  // f2092
  logic [0:0] f2092_wen;
  logic [31:0] f2092_wdata;
  logic [0:0] f2092_clk;
  logic [0:0] f2092_rst;
  logic [31:0] f2092_rdata;
  sr_buffer_32_1 f2092(.wen(f2092_wen), .wdata(f2092_wdata), .clk(f2092_clk), .rst(f2092_rst), .rdata(f2092_rdata));
  assign f2092_clk = clk;
  assign f2092_rst = rst;
  // Bindings to f2092

  // f2094
  logic [0:0] f2094_wen;
  logic [31:0] f2094_wdata;
  logic [0:0] f2094_clk;
  logic [0:0] f2094_rst;
  logic [31:0] f2094_rdata;
  sr_buffer_32_1 f2094(.wen(f2094_wen), .wdata(f2094_wdata), .clk(f2094_clk), .rst(f2094_rst), .rdata(f2094_rdata));
  assign f2094_clk = clk;
  assign f2094_rst = rst;
  // Bindings to f2094

  // f2096
  logic [0:0] f2096_wen;
  logic [31:0] f2096_wdata;
  logic [0:0] f2096_clk;
  logic [0:0] f2096_rst;
  logic [31:0] f2096_rdata;
  sr_buffer_32_1 f2096(.wen(f2096_wen), .wdata(f2096_wdata), .clk(f2096_clk), .rst(f2096_rst), .rdata(f2096_rdata));
  assign f2096_clk = clk;
  assign f2096_rst = rst;
  // Bindings to f2096

  // f2098
  logic [0:0] f2098_wen;
  logic [31:0] f2098_wdata;
  logic [0:0] f2098_clk;
  logic [0:0] f2098_rst;
  logic [31:0] f2098_rdata;
  sr_buffer_32_1 f2098(.wen(f2098_wen), .wdata(f2098_wdata), .clk(f2098_clk), .rst(f2098_rst), .rdata(f2098_rdata));
  assign f2098_clk = clk;
  assign f2098_rst = rst;
  // Bindings to f2098

  // f2100
  logic [0:0] f2100_wen;
  logic [31:0] f2100_wdata;
  logic [0:0] f2100_clk;
  logic [0:0] f2100_rst;
  logic [31:0] f2100_rdata;
  sr_buffer_32_1 f2100(.wen(f2100_wen), .wdata(f2100_wdata), .clk(f2100_clk), .rst(f2100_rst), .rdata(f2100_rdata));
  assign f2100_clk = clk;
  assign f2100_rst = rst;
  // Bindings to f2100

  // f2102
  logic [0:0] f2102_wen;
  logic [31:0] f2102_wdata;
  logic [0:0] f2102_clk;
  logic [0:0] f2102_rst;
  logic [31:0] f2102_rdata;
  sr_buffer_32_1 f2102(.wen(f2102_wen), .wdata(f2102_wdata), .clk(f2102_clk), .rst(f2102_rst), .rdata(f2102_rdata));
  assign f2102_clk = clk;
  assign f2102_rst = rst;
  // Bindings to f2102

  // f2104
  logic [0:0] f2104_wen;
  logic [31:0] f2104_wdata;
  logic [0:0] f2104_clk;
  logic [0:0] f2104_rst;
  logic [31:0] f2104_rdata;
  sr_buffer_32_1 f2104(.wen(f2104_wen), .wdata(f2104_wdata), .clk(f2104_clk), .rst(f2104_rst), .rdata(f2104_rdata));
  assign f2104_clk = clk;
  assign f2104_rst = rst;
  // Bindings to f2104

  // f2106
  logic [0:0] f2106_wen;
  logic [31:0] f2106_wdata;
  logic [0:0] f2106_clk;
  logic [0:0] f2106_rst;
  logic [31:0] f2106_rdata;
  sr_buffer_32_1 f2106(.wen(f2106_wen), .wdata(f2106_wdata), .clk(f2106_clk), .rst(f2106_rst), .rdata(f2106_rdata));
  assign f2106_clk = clk;
  assign f2106_rst = rst;
  // Bindings to f2106

  // f2108
  logic [0:0] f2108_wen;
  logic [31:0] f2108_wdata;
  logic [0:0] f2108_clk;
  logic [0:0] f2108_rst;
  logic [31:0] f2108_rdata;
  sr_buffer_32_1 f2108(.wen(f2108_wen), .wdata(f2108_wdata), .clk(f2108_clk), .rst(f2108_rst), .rdata(f2108_rdata));
  assign f2108_clk = clk;
  assign f2108_rst = rst;
  // Bindings to f2108

  // f2110
  logic [0:0] f2110_wen;
  logic [31:0] f2110_wdata;
  logic [0:0] f2110_clk;
  logic [0:0] f2110_rst;
  logic [31:0] f2110_rdata;
  sr_buffer_32_1 f2110(.wen(f2110_wen), .wdata(f2110_wdata), .clk(f2110_clk), .rst(f2110_rst), .rdata(f2110_rdata));
  assign f2110_clk = clk;
  assign f2110_rst = rst;
  // Bindings to f2110

  // f2112
  logic [0:0] f2112_wen;
  logic [31:0] f2112_wdata;
  logic [0:0] f2112_clk;
  logic [0:0] f2112_rst;
  logic [31:0] f2112_rdata;
  sr_buffer_32_1 f2112(.wen(f2112_wen), .wdata(f2112_wdata), .clk(f2112_clk), .rst(f2112_rst), .rdata(f2112_rdata));
  assign f2112_clk = clk;
  assign f2112_rst = rst;
  // Bindings to f2112

  // f2114
  logic [0:0] f2114_wen;
  logic [31:0] f2114_wdata;
  logic [0:0] f2114_clk;
  logic [0:0] f2114_rst;
  logic [31:0] f2114_rdata;
  sr_buffer_32_1 f2114(.wen(f2114_wen), .wdata(f2114_wdata), .clk(f2114_clk), .rst(f2114_rst), .rdata(f2114_rdata));
  assign f2114_clk = clk;
  assign f2114_rst = rst;
  // Bindings to f2114

  // f2116
  logic [0:0] f2116_wen;
  logic [31:0] f2116_wdata;
  logic [0:0] f2116_clk;
  logic [0:0] f2116_rst;
  logic [31:0] f2116_rdata;
  sr_buffer_32_1 f2116(.wen(f2116_wen), .wdata(f2116_wdata), .clk(f2116_clk), .rst(f2116_rst), .rdata(f2116_rdata));
  assign f2116_clk = clk;
  assign f2116_rst = rst;
  // Bindings to f2116

  // f2118
  logic [0:0] f2118_wen;
  logic [31:0] f2118_wdata;
  logic [0:0] f2118_clk;
  logic [0:0] f2118_rst;
  logic [31:0] f2118_rdata;
  sr_buffer_32_1 f2118(.wen(f2118_wen), .wdata(f2118_wdata), .clk(f2118_clk), .rst(f2118_rst), .rdata(f2118_rdata));
  assign f2118_clk = clk;
  assign f2118_rst = rst;
  // Bindings to f2118

  // f2120
  logic [0:0] f2120_wen;
  logic [31:0] f2120_wdata;
  logic [0:0] f2120_clk;
  logic [0:0] f2120_rst;
  logic [31:0] f2120_rdata;
  sr_buffer_32_1 f2120(.wen(f2120_wen), .wdata(f2120_wdata), .clk(f2120_clk), .rst(f2120_rst), .rdata(f2120_rdata));
  assign f2120_clk = clk;
  assign f2120_rst = rst;
  // Bindings to f2120

  // f2122
  logic [0:0] f2122_wen;
  logic [31:0] f2122_wdata;
  logic [0:0] f2122_clk;
  logic [0:0] f2122_rst;
  logic [31:0] f2122_rdata;
  sr_buffer_32_1 f2122(.wen(f2122_wen), .wdata(f2122_wdata), .clk(f2122_clk), .rst(f2122_rst), .rdata(f2122_rdata));
  assign f2122_clk = clk;
  assign f2122_rst = rst;
  // Bindings to f2122

  // f2124
  logic [0:0] f2124_wen;
  logic [31:0] f2124_wdata;
  logic [0:0] f2124_clk;
  logic [0:0] f2124_rst;
  logic [31:0] f2124_rdata;
  sr_buffer_32_1 f2124(.wen(f2124_wen), .wdata(f2124_wdata), .clk(f2124_clk), .rst(f2124_rst), .rdata(f2124_rdata));
  assign f2124_clk = clk;
  assign f2124_rst = rst;
  // Bindings to f2124

  // f2126
  logic [0:0] f2126_wen;
  logic [31:0] f2126_wdata;
  logic [0:0] f2126_clk;
  logic [0:0] f2126_rst;
  logic [31:0] f2126_rdata;
  sr_buffer_32_1 f2126(.wen(f2126_wen), .wdata(f2126_wdata), .clk(f2126_clk), .rst(f2126_rst), .rdata(f2126_rdata));
  assign f2126_clk = clk;
  assign f2126_rst = rst;
  // Bindings to f2126

  // f2128
  logic [0:0] f2128_wen;
  logic [31:0] f2128_wdata;
  logic [0:0] f2128_clk;
  logic [0:0] f2128_rst;
  logic [31:0] f2128_rdata;
  sr_buffer_32_1 f2128(.wen(f2128_wen), .wdata(f2128_wdata), .clk(f2128_clk), .rst(f2128_rst), .rdata(f2128_rdata));
  assign f2128_clk = clk;
  assign f2128_rst = rst;
  // Bindings to f2128

  // f2130
  logic [0:0] f2130_wen;
  logic [31:0] f2130_wdata;
  logic [0:0] f2130_clk;
  logic [0:0] f2130_rst;
  logic [31:0] f2130_rdata;
  sr_buffer_32_1 f2130(.wen(f2130_wen), .wdata(f2130_wdata), .clk(f2130_clk), .rst(f2130_rst), .rdata(f2130_rdata));
  assign f2130_clk = clk;
  assign f2130_rst = rst;
  // Bindings to f2130

  // f2132
  logic [0:0] f2132_wen;
  logic [31:0] f2132_wdata;
  logic [0:0] f2132_clk;
  logic [0:0] f2132_rst;
  logic [31:0] f2132_rdata;
  sr_buffer_32_1 f2132(.wen(f2132_wen), .wdata(f2132_wdata), .clk(f2132_clk), .rst(f2132_rst), .rdata(f2132_rdata));
  assign f2132_clk = clk;
  assign f2132_rst = rst;
  // Bindings to f2132

  // f2134
  logic [0:0] f2134_wen;
  logic [31:0] f2134_wdata;
  logic [0:0] f2134_clk;
  logic [0:0] f2134_rst;
  logic [31:0] f2134_rdata;
  sr_buffer_32_1 f2134(.wen(f2134_wen), .wdata(f2134_wdata), .clk(f2134_clk), .rst(f2134_rst), .rdata(f2134_rdata));
  assign f2134_clk = clk;
  assign f2134_rst = rst;
  // Bindings to f2134

  // f2136
  logic [0:0] f2136_wen;
  logic [31:0] f2136_wdata;
  logic [0:0] f2136_clk;
  logic [0:0] f2136_rst;
  logic [31:0] f2136_rdata;
  sr_buffer_32_1 f2136(.wen(f2136_wen), .wdata(f2136_wdata), .clk(f2136_clk), .rst(f2136_rst), .rdata(f2136_rdata));
  assign f2136_clk = clk;
  assign f2136_rst = rst;
  // Bindings to f2136

  // f2138
  logic [0:0] f2138_wen;
  logic [31:0] f2138_wdata;
  logic [0:0] f2138_clk;
  logic [0:0] f2138_rst;
  logic [31:0] f2138_rdata;
  sr_buffer_32_1 f2138(.wen(f2138_wen), .wdata(f2138_wdata), .clk(f2138_clk), .rst(f2138_rst), .rdata(f2138_rdata));
  assign f2138_clk = clk;
  assign f2138_rst = rst;
  // Bindings to f2138

  // f2140
  logic [0:0] f2140_wen;
  logic [31:0] f2140_wdata;
  logic [0:0] f2140_clk;
  logic [0:0] f2140_rst;
  logic [31:0] f2140_rdata;
  sr_buffer_32_1 f2140(.wen(f2140_wen), .wdata(f2140_wdata), .clk(f2140_clk), .rst(f2140_rst), .rdata(f2140_rdata));
  assign f2140_clk = clk;
  assign f2140_rst = rst;
  // Bindings to f2140

  // f2142
  logic [0:0] f2142_wen;
  logic [31:0] f2142_wdata;
  logic [0:0] f2142_clk;
  logic [0:0] f2142_rst;
  logic [31:0] f2142_rdata;
  sr_buffer_32_1 f2142(.wen(f2142_wen), .wdata(f2142_wdata), .clk(f2142_clk), .rst(f2142_rst), .rdata(f2142_rdata));
  assign f2142_clk = clk;
  assign f2142_rst = rst;
  // Bindings to f2142

  // f2144
  logic [0:0] f2144_wen;
  logic [31:0] f2144_wdata;
  logic [0:0] f2144_clk;
  logic [0:0] f2144_rst;
  logic [31:0] f2144_rdata;
  sr_buffer_32_1 f2144(.wen(f2144_wen), .wdata(f2144_wdata), .clk(f2144_clk), .rst(f2144_rst), .rdata(f2144_rdata));
  assign f2144_clk = clk;
  assign f2144_rst = rst;
  // Bindings to f2144

  // f2146
  logic [0:0] f2146_wen;
  logic [31:0] f2146_wdata;
  logic [0:0] f2146_clk;
  logic [0:0] f2146_rst;
  logic [31:0] f2146_rdata;
  sr_buffer_32_1 f2146(.wen(f2146_wen), .wdata(f2146_wdata), .clk(f2146_clk), .rst(f2146_rst), .rdata(f2146_rdata));
  assign f2146_clk = clk;
  assign f2146_rst = rst;
  // Bindings to f2146

  // f2148
  logic [0:0] f2148_wen;
  logic [31:0] f2148_wdata;
  logic [0:0] f2148_clk;
  logic [0:0] f2148_rst;
  logic [31:0] f2148_rdata;
  sr_buffer_32_1 f2148(.wen(f2148_wen), .wdata(f2148_wdata), .clk(f2148_clk), .rst(f2148_rst), .rdata(f2148_rdata));
  assign f2148_clk = clk;
  assign f2148_rst = rst;
  // Bindings to f2148

  // f2150
  logic [0:0] f2150_wen;
  logic [31:0] f2150_wdata;
  logic [0:0] f2150_clk;
  logic [0:0] f2150_rst;
  logic [31:0] f2150_rdata;
  sr_buffer_32_1 f2150(.wen(f2150_wen), .wdata(f2150_wdata), .clk(f2150_clk), .rst(f2150_rst), .rdata(f2150_rdata));
  assign f2150_clk = clk;
  assign f2150_rst = rst;
  // Bindings to f2150

  // f2152
  logic [0:0] f2152_wen;
  logic [31:0] f2152_wdata;
  logic [0:0] f2152_clk;
  logic [0:0] f2152_rst;
  logic [31:0] f2152_rdata;
  sr_buffer_32_1 f2152(.wen(f2152_wen), .wdata(f2152_wdata), .clk(f2152_clk), .rst(f2152_rst), .rdata(f2152_rdata));
  assign f2152_clk = clk;
  assign f2152_rst = rst;
  // Bindings to f2152

  // f2154
  logic [0:0] f2154_wen;
  logic [31:0] f2154_wdata;
  logic [0:0] f2154_clk;
  logic [0:0] f2154_rst;
  logic [31:0] f2154_rdata;
  sr_buffer_32_1 f2154(.wen(f2154_wen), .wdata(f2154_wdata), .clk(f2154_clk), .rst(f2154_rst), .rdata(f2154_rdata));
  assign f2154_clk = clk;
  assign f2154_rst = rst;
  // Bindings to f2154

  // f2156
  logic [0:0] f2156_wen;
  logic [31:0] f2156_wdata;
  logic [0:0] f2156_clk;
  logic [0:0] f2156_rst;
  logic [31:0] f2156_rdata;
  sr_buffer_32_1 f2156(.wen(f2156_wen), .wdata(f2156_wdata), .clk(f2156_clk), .rst(f2156_rst), .rdata(f2156_rdata));
  assign f2156_clk = clk;
  assign f2156_rst = rst;
  // Bindings to f2156

  // f2158
  logic [0:0] f2158_wen;
  logic [31:0] f2158_wdata;
  logic [0:0] f2158_clk;
  logic [0:0] f2158_rst;
  logic [31:0] f2158_rdata;
  sr_buffer_32_1 f2158(.wen(f2158_wen), .wdata(f2158_wdata), .clk(f2158_clk), .rst(f2158_rst), .rdata(f2158_rdata));
  assign f2158_clk = clk;
  assign f2158_rst = rst;
  // Bindings to f2158

  // f2160
  logic [0:0] f2160_wen;
  logic [31:0] f2160_wdata;
  logic [0:0] f2160_clk;
  logic [0:0] f2160_rst;
  logic [31:0] f2160_rdata;
  sr_buffer_32_1 f2160(.wen(f2160_wen), .wdata(f2160_wdata), .clk(f2160_clk), .rst(f2160_rst), .rdata(f2160_rdata));
  assign f2160_clk = clk;
  assign f2160_rst = rst;
  // Bindings to f2160

  // f2162
  logic [0:0] f2162_wen;
  logic [31:0] f2162_wdata;
  logic [0:0] f2162_clk;
  logic [0:0] f2162_rst;
  logic [31:0] f2162_rdata;
  sr_buffer_32_1 f2162(.wen(f2162_wen), .wdata(f2162_wdata), .clk(f2162_clk), .rst(f2162_rst), .rdata(f2162_rdata));
  assign f2162_clk = clk;
  assign f2162_rst = rst;
  // Bindings to f2162

  // f2164
  logic [0:0] f2164_wen;
  logic [31:0] f2164_wdata;
  logic [0:0] f2164_clk;
  logic [0:0] f2164_rst;
  logic [31:0] f2164_rdata;
  sr_buffer_32_1 f2164(.wen(f2164_wen), .wdata(f2164_wdata), .clk(f2164_clk), .rst(f2164_rst), .rdata(f2164_rdata));
  assign f2164_clk = clk;
  assign f2164_rst = rst;
  // Bindings to f2164

  // f2166
  logic [0:0] f2166_wen;
  logic [31:0] f2166_wdata;
  logic [0:0] f2166_clk;
  logic [0:0] f2166_rst;
  logic [31:0] f2166_rdata;
  sr_buffer_32_1 f2166(.wen(f2166_wen), .wdata(f2166_wdata), .clk(f2166_clk), .rst(f2166_rst), .rdata(f2166_rdata));
  assign f2166_clk = clk;
  assign f2166_rst = rst;
  // Bindings to f2166

  // f2168
  logic [0:0] f2168_wen;
  logic [31:0] f2168_wdata;
  logic [0:0] f2168_clk;
  logic [0:0] f2168_rst;
  logic [31:0] f2168_rdata;
  sr_buffer_32_1 f2168(.wen(f2168_wen), .wdata(f2168_wdata), .clk(f2168_clk), .rst(f2168_rst), .rdata(f2168_rdata));
  assign f2168_clk = clk;
  assign f2168_rst = rst;
  // Bindings to f2168

  // f2170
  logic [0:0] f2170_wen;
  logic [31:0] f2170_wdata;
  logic [0:0] f2170_clk;
  logic [0:0] f2170_rst;
  logic [31:0] f2170_rdata;
  sr_buffer_32_1 f2170(.wen(f2170_wen), .wdata(f2170_wdata), .clk(f2170_clk), .rst(f2170_rst), .rdata(f2170_rdata));
  assign f2170_clk = clk;
  assign f2170_rst = rst;
  // Bindings to f2170

  // f2172
  logic [0:0] f2172_wen;
  logic [31:0] f2172_wdata;
  logic [0:0] f2172_clk;
  logic [0:0] f2172_rst;
  logic [31:0] f2172_rdata;
  sr_buffer_32_1 f2172(.wen(f2172_wen), .wdata(f2172_wdata), .clk(f2172_clk), .rst(f2172_rst), .rdata(f2172_rdata));
  assign f2172_clk = clk;
  assign f2172_rst = rst;
  // Bindings to f2172

  // f2174
  logic [0:0] f2174_wen;
  logic [31:0] f2174_wdata;
  logic [0:0] f2174_clk;
  logic [0:0] f2174_rst;
  logic [31:0] f2174_rdata;
  sr_buffer_32_1 f2174(.wen(f2174_wen), .wdata(f2174_wdata), .clk(f2174_clk), .rst(f2174_rst), .rdata(f2174_rdata));
  assign f2174_clk = clk;
  assign f2174_rst = rst;
  // Bindings to f2174

  // f2176
  logic [0:0] f2176_wen;
  logic [31:0] f2176_wdata;
  logic [0:0] f2176_clk;
  logic [0:0] f2176_rst;
  logic [31:0] f2176_rdata;
  sr_buffer_32_1 f2176(.wen(f2176_wen), .wdata(f2176_wdata), .clk(f2176_clk), .rst(f2176_rst), .rdata(f2176_rdata));
  assign f2176_clk = clk;
  assign f2176_rst = rst;
  // Bindings to f2176

  // f2178
  logic [0:0] f2178_wen;
  logic [31:0] f2178_wdata;
  logic [0:0] f2178_clk;
  logic [0:0] f2178_rst;
  logic [31:0] f2178_rdata;
  sr_buffer_32_1 f2178(.wen(f2178_wen), .wdata(f2178_wdata), .clk(f2178_clk), .rst(f2178_rst), .rdata(f2178_rdata));
  assign f2178_clk = clk;
  assign f2178_rst = rst;
  // Bindings to f2178

  // f2180
  logic [0:0] f2180_wen;
  logic [31:0] f2180_wdata;
  logic [0:0] f2180_clk;
  logic [0:0] f2180_rst;
  logic [31:0] f2180_rdata;
  sr_buffer_32_1 f2180(.wen(f2180_wen), .wdata(f2180_wdata), .clk(f2180_clk), .rst(f2180_rst), .rdata(f2180_rdata));
  assign f2180_clk = clk;
  assign f2180_rst = rst;
  // Bindings to f2180

  // f2182
  logic [0:0] f2182_wen;
  logic [31:0] f2182_wdata;
  logic [0:0] f2182_clk;
  logic [0:0] f2182_rst;
  logic [31:0] f2182_rdata;
  sr_buffer_32_1 f2182(.wen(f2182_wen), .wdata(f2182_wdata), .clk(f2182_clk), .rst(f2182_rst), .rdata(f2182_rdata));
  assign f2182_clk = clk;
  assign f2182_rst = rst;
  // Bindings to f2182

  // f2184
  logic [0:0] f2184_wen;
  logic [31:0] f2184_wdata;
  logic [0:0] f2184_clk;
  logic [0:0] f2184_rst;
  logic [31:0] f2184_rdata;
  sr_buffer_32_1 f2184(.wen(f2184_wen), .wdata(f2184_wdata), .clk(f2184_clk), .rst(f2184_rst), .rdata(f2184_rdata));
  assign f2184_clk = clk;
  assign f2184_rst = rst;
  // Bindings to f2184

  // f2186
  logic [0:0] f2186_wen;
  logic [31:0] f2186_wdata;
  logic [0:0] f2186_clk;
  logic [0:0] f2186_rst;
  logic [31:0] f2186_rdata;
  sr_buffer_32_1 f2186(.wen(f2186_wen), .wdata(f2186_wdata), .clk(f2186_clk), .rst(f2186_rst), .rdata(f2186_rdata));
  assign f2186_clk = clk;
  assign f2186_rst = rst;
  // Bindings to f2186

  // f2188
  logic [0:0] f2188_wen;
  logic [31:0] f2188_wdata;
  logic [0:0] f2188_clk;
  logic [0:0] f2188_rst;
  logic [31:0] f2188_rdata;
  sr_buffer_32_1 f2188(.wen(f2188_wen), .wdata(f2188_wdata), .clk(f2188_clk), .rst(f2188_rst), .rdata(f2188_rdata));
  assign f2188_clk = clk;
  assign f2188_rst = rst;
  // Bindings to f2188

  // f2190
  logic [0:0] f2190_wen;
  logic [31:0] f2190_wdata;
  logic [0:0] f2190_clk;
  logic [0:0] f2190_rst;
  logic [31:0] f2190_rdata;
  sr_buffer_32_1 f2190(.wen(f2190_wen), .wdata(f2190_wdata), .clk(f2190_clk), .rst(f2190_rst), .rdata(f2190_rdata));
  assign f2190_clk = clk;
  assign f2190_rst = rst;
  // Bindings to f2190

  // f2192
  logic [0:0] f2192_wen;
  logic [31:0] f2192_wdata;
  logic [0:0] f2192_clk;
  logic [0:0] f2192_rst;
  logic [31:0] f2192_rdata;
  sr_buffer_32_1 f2192(.wen(f2192_wen), .wdata(f2192_wdata), .clk(f2192_clk), .rst(f2192_rst), .rdata(f2192_rdata));
  assign f2192_clk = clk;
  assign f2192_rst = rst;
  // Bindings to f2192

  // f2194
  logic [0:0] f2194_wen;
  logic [31:0] f2194_wdata;
  logic [0:0] f2194_clk;
  logic [0:0] f2194_rst;
  logic [31:0] f2194_rdata;
  sr_buffer_32_1 f2194(.wen(f2194_wen), .wdata(f2194_wdata), .clk(f2194_clk), .rst(f2194_rst), .rdata(f2194_rdata));
  assign f2194_clk = clk;
  assign f2194_rst = rst;
  // Bindings to f2194

  // f2196
  logic [0:0] f2196_wen;
  logic [31:0] f2196_wdata;
  logic [0:0] f2196_clk;
  logic [0:0] f2196_rst;
  logic [31:0] f2196_rdata;
  sr_buffer_32_1 f2196(.wen(f2196_wen), .wdata(f2196_wdata), .clk(f2196_clk), .rst(f2196_rst), .rdata(f2196_rdata));
  assign f2196_clk = clk;
  assign f2196_rst = rst;
  // Bindings to f2196

  // f2198
  logic [0:0] f2198_wen;
  logic [31:0] f2198_wdata;
  logic [0:0] f2198_clk;
  logic [0:0] f2198_rst;
  logic [31:0] f2198_rdata;
  sr_buffer_32_1 f2198(.wen(f2198_wen), .wdata(f2198_wdata), .clk(f2198_clk), .rst(f2198_rst), .rdata(f2198_rdata));
  assign f2198_clk = clk;
  assign f2198_rst = rst;
  // Bindings to f2198

  // f2200
  logic [0:0] f2200_wen;
  logic [31:0] f2200_wdata;
  logic [0:0] f2200_clk;
  logic [0:0] f2200_rst;
  logic [31:0] f2200_rdata;
  sr_buffer_32_1 f2200(.wen(f2200_wen), .wdata(f2200_wdata), .clk(f2200_clk), .rst(f2200_rst), .rdata(f2200_rdata));
  assign f2200_clk = clk;
  assign f2200_rst = rst;
  // Bindings to f2200

  // f2202
  logic [0:0] f2202_wen;
  logic [31:0] f2202_wdata;
  logic [0:0] f2202_clk;
  logic [0:0] f2202_rst;
  logic [31:0] f2202_rdata;
  sr_buffer_32_1 f2202(.wen(f2202_wen), .wdata(f2202_wdata), .clk(f2202_clk), .rst(f2202_rst), .rdata(f2202_rdata));
  assign f2202_clk = clk;
  assign f2202_rst = rst;
  // Bindings to f2202

  // f2204
  logic [0:0] f2204_wen;
  logic [31:0] f2204_wdata;
  logic [0:0] f2204_clk;
  logic [0:0] f2204_rst;
  logic [31:0] f2204_rdata;
  sr_buffer_32_1 f2204(.wen(f2204_wen), .wdata(f2204_wdata), .clk(f2204_clk), .rst(f2204_rst), .rdata(f2204_rdata));
  assign f2204_clk = clk;
  assign f2204_rst = rst;
  // Bindings to f2204

  // f2206
  logic [0:0] f2206_wen;
  logic [31:0] f2206_wdata;
  logic [0:0] f2206_clk;
  logic [0:0] f2206_rst;
  logic [31:0] f2206_rdata;
  sr_buffer_32_1 f2206(.wen(f2206_wen), .wdata(f2206_wdata), .clk(f2206_clk), .rst(f2206_rst), .rdata(f2206_rdata));
  assign f2206_clk = clk;
  assign f2206_rst = rst;
  // Bindings to f2206

  // f2208
  logic [0:0] f2208_wen;
  logic [31:0] f2208_wdata;
  logic [0:0] f2208_clk;
  logic [0:0] f2208_rst;
  logic [31:0] f2208_rdata;
  sr_buffer_32_1 f2208(.wen(f2208_wen), .wdata(f2208_wdata), .clk(f2208_clk), .rst(f2208_rst), .rdata(f2208_rdata));
  assign f2208_clk = clk;
  assign f2208_rst = rst;
  // Bindings to f2208

  // f2210
  logic [0:0] f2210_wen;
  logic [31:0] f2210_wdata;
  logic [0:0] f2210_clk;
  logic [0:0] f2210_rst;
  logic [31:0] f2210_rdata;
  sr_buffer_32_1 f2210(.wen(f2210_wen), .wdata(f2210_wdata), .clk(f2210_clk), .rst(f2210_rst), .rdata(f2210_rdata));
  assign f2210_clk = clk;
  assign f2210_rst = rst;
  // Bindings to f2210

  // f2212
  logic [0:0] f2212_wen;
  logic [31:0] f2212_wdata;
  logic [0:0] f2212_clk;
  logic [0:0] f2212_rst;
  logic [31:0] f2212_rdata;
  sr_buffer_32_1 f2212(.wen(f2212_wen), .wdata(f2212_wdata), .clk(f2212_clk), .rst(f2212_rst), .rdata(f2212_rdata));
  assign f2212_clk = clk;
  assign f2212_rst = rst;
  // Bindings to f2212

  // f2214
  logic [0:0] f2214_wen;
  logic [31:0] f2214_wdata;
  logic [0:0] f2214_clk;
  logic [0:0] f2214_rst;
  logic [31:0] f2214_rdata;
  sr_buffer_32_1 f2214(.wen(f2214_wen), .wdata(f2214_wdata), .clk(f2214_clk), .rst(f2214_rst), .rdata(f2214_rdata));
  assign f2214_clk = clk;
  assign f2214_rst = rst;
  // Bindings to f2214

  // f2216
  logic [0:0] f2216_wen;
  logic [31:0] f2216_wdata;
  logic [0:0] f2216_clk;
  logic [0:0] f2216_rst;
  logic [31:0] f2216_rdata;
  sr_buffer_32_1 f2216(.wen(f2216_wen), .wdata(f2216_wdata), .clk(f2216_clk), .rst(f2216_rst), .rdata(f2216_rdata));
  assign f2216_clk = clk;
  assign f2216_rst = rst;
  // Bindings to f2216

  // f2218
  logic [0:0] f2218_wen;
  logic [31:0] f2218_wdata;
  logic [0:0] f2218_clk;
  logic [0:0] f2218_rst;
  logic [31:0] f2218_rdata;
  sr_buffer_32_1 f2218(.wen(f2218_wen), .wdata(f2218_wdata), .clk(f2218_clk), .rst(f2218_rst), .rdata(f2218_rdata));
  assign f2218_clk = clk;
  assign f2218_rst = rst;
  // Bindings to f2218

  // f2220
  logic [0:0] f2220_wen;
  logic [31:0] f2220_wdata;
  logic [0:0] f2220_clk;
  logic [0:0] f2220_rst;
  logic [31:0] f2220_rdata;
  sr_buffer_32_1 f2220(.wen(f2220_wen), .wdata(f2220_wdata), .clk(f2220_clk), .rst(f2220_rst), .rdata(f2220_rdata));
  assign f2220_clk = clk;
  assign f2220_rst = rst;
  // Bindings to f2220

  // f2222
  logic [0:0] f2222_wen;
  logic [31:0] f2222_wdata;
  logic [0:0] f2222_clk;
  logic [0:0] f2222_rst;
  logic [31:0] f2222_rdata;
  sr_buffer_32_1 f2222(.wen(f2222_wen), .wdata(f2222_wdata), .clk(f2222_clk), .rst(f2222_rst), .rdata(f2222_rdata));
  assign f2222_clk = clk;
  assign f2222_rst = rst;
  // Bindings to f2222

  // f2224
  logic [0:0] f2224_wen;
  logic [31:0] f2224_wdata;
  logic [0:0] f2224_clk;
  logic [0:0] f2224_rst;
  logic [31:0] f2224_rdata;
  sr_buffer_32_1 f2224(.wen(f2224_wen), .wdata(f2224_wdata), .clk(f2224_clk), .rst(f2224_rst), .rdata(f2224_rdata));
  assign f2224_clk = clk;
  assign f2224_rst = rst;
  // Bindings to f2224

  // f2226
  logic [0:0] f2226_wen;
  logic [31:0] f2226_wdata;
  logic [0:0] f2226_clk;
  logic [0:0] f2226_rst;
  logic [31:0] f2226_rdata;
  sr_buffer_32_1 f2226(.wen(f2226_wen), .wdata(f2226_wdata), .clk(f2226_clk), .rst(f2226_rst), .rdata(f2226_rdata));
  assign f2226_clk = clk;
  assign f2226_rst = rst;
  // Bindings to f2226

  // f2228
  logic [0:0] f2228_wen;
  logic [31:0] f2228_wdata;
  logic [0:0] f2228_clk;
  logic [0:0] f2228_rst;
  logic [31:0] f2228_rdata;
  sr_buffer_32_1 f2228(.wen(f2228_wen), .wdata(f2228_wdata), .clk(f2228_clk), .rst(f2228_rst), .rdata(f2228_rdata));
  assign f2228_clk = clk;
  assign f2228_rst = rst;
  // Bindings to f2228

  // f2230
  logic [0:0] f2230_wen;
  logic [31:0] f2230_wdata;
  logic [0:0] f2230_clk;
  logic [0:0] f2230_rst;
  logic [31:0] f2230_rdata;
  sr_buffer_32_1 f2230(.wen(f2230_wen), .wdata(f2230_wdata), .clk(f2230_clk), .rst(f2230_rst), .rdata(f2230_rdata));
  assign f2230_clk = clk;
  assign f2230_rst = rst;
  // Bindings to f2230

  // f2232
  logic [0:0] f2232_wen;
  logic [31:0] f2232_wdata;
  logic [0:0] f2232_clk;
  logic [0:0] f2232_rst;
  logic [31:0] f2232_rdata;
  sr_buffer_32_1 f2232(.wen(f2232_wen), .wdata(f2232_wdata), .clk(f2232_clk), .rst(f2232_rst), .rdata(f2232_rdata));
  assign f2232_clk = clk;
  assign f2232_rst = rst;
  // Bindings to f2232

  // f2234
  logic [0:0] f2234_wen;
  logic [31:0] f2234_wdata;
  logic [0:0] f2234_clk;
  logic [0:0] f2234_rst;
  logic [31:0] f2234_rdata;
  sr_buffer_32_1 f2234(.wen(f2234_wen), .wdata(f2234_wdata), .clk(f2234_clk), .rst(f2234_rst), .rdata(f2234_rdata));
  assign f2234_clk = clk;
  assign f2234_rst = rst;
  // Bindings to f2234

  // f2236
  logic [0:0] f2236_wen;
  logic [31:0] f2236_wdata;
  logic [0:0] f2236_clk;
  logic [0:0] f2236_rst;
  logic [31:0] f2236_rdata;
  sr_buffer_32_1 f2236(.wen(f2236_wen), .wdata(f2236_wdata), .clk(f2236_clk), .rst(f2236_rst), .rdata(f2236_rdata));
  assign f2236_clk = clk;
  assign f2236_rst = rst;
  // Bindings to f2236

  // f2238
  logic [0:0] f2238_wen;
  logic [31:0] f2238_wdata;
  logic [0:0] f2238_clk;
  logic [0:0] f2238_rst;
  logic [31:0] f2238_rdata;
  sr_buffer_32_1 f2238(.wen(f2238_wen), .wdata(f2238_wdata), .clk(f2238_clk), .rst(f2238_rst), .rdata(f2238_rdata));
  assign f2238_clk = clk;
  assign f2238_rst = rst;
  // Bindings to f2238

  // f2240
  logic [0:0] f2240_wen;
  logic [31:0] f2240_wdata;
  logic [0:0] f2240_clk;
  logic [0:0] f2240_rst;
  logic [31:0] f2240_rdata;
  sr_buffer_32_1 f2240(.wen(f2240_wen), .wdata(f2240_wdata), .clk(f2240_clk), .rst(f2240_rst), .rdata(f2240_rdata));
  assign f2240_clk = clk;
  assign f2240_rst = rst;
  // Bindings to f2240

  // f2242
  logic [0:0] f2242_wen;
  logic [31:0] f2242_wdata;
  logic [0:0] f2242_clk;
  logic [0:0] f2242_rst;
  logic [31:0] f2242_rdata;
  sr_buffer_32_1 f2242(.wen(f2242_wen), .wdata(f2242_wdata), .clk(f2242_clk), .rst(f2242_rst), .rdata(f2242_rdata));
  assign f2242_clk = clk;
  assign f2242_rst = rst;
  // Bindings to f2242

  // f2244
  logic [0:0] f2244_wen;
  logic [31:0] f2244_wdata;
  logic [0:0] f2244_clk;
  logic [0:0] f2244_rst;
  logic [31:0] f2244_rdata;
  sr_buffer_32_1 f2244(.wen(f2244_wen), .wdata(f2244_wdata), .clk(f2244_clk), .rst(f2244_rst), .rdata(f2244_rdata));
  assign f2244_clk = clk;
  assign f2244_rst = rst;
  // Bindings to f2244

  // f2246
  logic [0:0] f2246_wen;
  logic [31:0] f2246_wdata;
  logic [0:0] f2246_clk;
  logic [0:0] f2246_rst;
  logic [31:0] f2246_rdata;
  sr_buffer_32_1 f2246(.wen(f2246_wen), .wdata(f2246_wdata), .clk(f2246_clk), .rst(f2246_rst), .rdata(f2246_rdata));
  assign f2246_clk = clk;
  assign f2246_rst = rst;
  // Bindings to f2246

  // f2248
  logic [0:0] f2248_wen;
  logic [31:0] f2248_wdata;
  logic [0:0] f2248_clk;
  logic [0:0] f2248_rst;
  logic [31:0] f2248_rdata;
  sr_buffer_32_1 f2248(.wen(f2248_wen), .wdata(f2248_wdata), .clk(f2248_clk), .rst(f2248_rst), .rdata(f2248_rdata));
  assign f2248_clk = clk;
  assign f2248_rst = rst;
  // Bindings to f2248

  // f2250
  logic [0:0] f2250_wen;
  logic [31:0] f2250_wdata;
  logic [0:0] f2250_clk;
  logic [0:0] f2250_rst;
  logic [31:0] f2250_rdata;
  sr_buffer_32_1 f2250(.wen(f2250_wen), .wdata(f2250_wdata), .clk(f2250_clk), .rst(f2250_rst), .rdata(f2250_rdata));
  assign f2250_clk = clk;
  assign f2250_rst = rst;
  // Bindings to f2250

  // f2252
  logic [0:0] f2252_wen;
  logic [31:0] f2252_wdata;
  logic [0:0] f2252_clk;
  logic [0:0] f2252_rst;
  logic [31:0] f2252_rdata;
  sr_buffer_32_1 f2252(.wen(f2252_wen), .wdata(f2252_wdata), .clk(f2252_clk), .rst(f2252_rst), .rdata(f2252_rdata));
  assign f2252_clk = clk;
  assign f2252_rst = rst;
  // Bindings to f2252

  // f2254
  logic [0:0] f2254_wen;
  logic [31:0] f2254_wdata;
  logic [0:0] f2254_clk;
  logic [0:0] f2254_rst;
  logic [31:0] f2254_rdata;
  sr_buffer_32_1 f2254(.wen(f2254_wen), .wdata(f2254_wdata), .clk(f2254_clk), .rst(f2254_rst), .rdata(f2254_rdata));
  assign f2254_clk = clk;
  assign f2254_rst = rst;
  // Bindings to f2254

  // f2256
  logic [0:0] f2256_wen;
  logic [31:0] f2256_wdata;
  logic [0:0] f2256_clk;
  logic [0:0] f2256_rst;
  logic [31:0] f2256_rdata;
  sr_buffer_32_1 f2256(.wen(f2256_wen), .wdata(f2256_wdata), .clk(f2256_clk), .rst(f2256_rst), .rdata(f2256_rdata));
  assign f2256_clk = clk;
  assign f2256_rst = rst;
  // Bindings to f2256

  // f2258
  logic [0:0] f2258_wen;
  logic [31:0] f2258_wdata;
  logic [0:0] f2258_clk;
  logic [0:0] f2258_rst;
  logic [31:0] f2258_rdata;
  sr_buffer_32_1 f2258(.wen(f2258_wen), .wdata(f2258_wdata), .clk(f2258_clk), .rst(f2258_rst), .rdata(f2258_rdata));
  assign f2258_clk = clk;
  assign f2258_rst = rst;
  // Bindings to f2258

  // f2260
  logic [0:0] f2260_wen;
  logic [31:0] f2260_wdata;
  logic [0:0] f2260_clk;
  logic [0:0] f2260_rst;
  logic [31:0] f2260_rdata;
  sr_buffer_32_1 f2260(.wen(f2260_wen), .wdata(f2260_wdata), .clk(f2260_clk), .rst(f2260_rst), .rdata(f2260_rdata));
  assign f2260_clk = clk;
  assign f2260_rst = rst;
  // Bindings to f2260

  // f2262
  logic [0:0] f2262_wen;
  logic [31:0] f2262_wdata;
  logic [0:0] f2262_clk;
  logic [0:0] f2262_rst;
  logic [31:0] f2262_rdata;
  sr_buffer_32_1 f2262(.wen(f2262_wen), .wdata(f2262_wdata), .clk(f2262_clk), .rst(f2262_rst), .rdata(f2262_rdata));
  assign f2262_clk = clk;
  assign f2262_rst = rst;
  // Bindings to f2262

  // f2264
  logic [0:0] f2264_wen;
  logic [31:0] f2264_wdata;
  logic [0:0] f2264_clk;
  logic [0:0] f2264_rst;
  logic [31:0] f2264_rdata;
  sr_buffer_32_1 f2264(.wen(f2264_wen), .wdata(f2264_wdata), .clk(f2264_clk), .rst(f2264_rst), .rdata(f2264_rdata));
  assign f2264_clk = clk;
  assign f2264_rst = rst;
  // Bindings to f2264

  // f2266
  logic [0:0] f2266_wen;
  logic [31:0] f2266_wdata;
  logic [0:0] f2266_clk;
  logic [0:0] f2266_rst;
  logic [31:0] f2266_rdata;
  sr_buffer_32_1 f2266(.wen(f2266_wen), .wdata(f2266_wdata), .clk(f2266_clk), .rst(f2266_rst), .rdata(f2266_rdata));
  assign f2266_clk = clk;
  assign f2266_rst = rst;
  // Bindings to f2266

  // f2268
  logic [0:0] f2268_wen;
  logic [31:0] f2268_wdata;
  logic [0:0] f2268_clk;
  logic [0:0] f2268_rst;
  logic [31:0] f2268_rdata;
  sr_buffer_32_1 f2268(.wen(f2268_wen), .wdata(f2268_wdata), .clk(f2268_clk), .rst(f2268_rst), .rdata(f2268_rdata));
  assign f2268_clk = clk;
  assign f2268_rst = rst;
  // Bindings to f2268

  // f2270
  logic [0:0] f2270_wen;
  logic [31:0] f2270_wdata;
  logic [0:0] f2270_clk;
  logic [0:0] f2270_rst;
  logic [31:0] f2270_rdata;
  sr_buffer_32_1 f2270(.wen(f2270_wen), .wdata(f2270_wdata), .clk(f2270_clk), .rst(f2270_rst), .rdata(f2270_rdata));
  assign f2270_clk = clk;
  assign f2270_rst = rst;
  // Bindings to f2270

  // f2272
  logic [0:0] f2272_wen;
  logic [31:0] f2272_wdata;
  logic [0:0] f2272_clk;
  logic [0:0] f2272_rst;
  logic [31:0] f2272_rdata;
  sr_buffer_32_1 f2272(.wen(f2272_wen), .wdata(f2272_wdata), .clk(f2272_clk), .rst(f2272_rst), .rdata(f2272_rdata));
  assign f2272_clk = clk;
  assign f2272_rst = rst;
  // Bindings to f2272

  // f2274
  logic [0:0] f2274_wen;
  logic [31:0] f2274_wdata;
  logic [0:0] f2274_clk;
  logic [0:0] f2274_rst;
  logic [31:0] f2274_rdata;
  sr_buffer_32_1 f2274(.wen(f2274_wen), .wdata(f2274_wdata), .clk(f2274_clk), .rst(f2274_rst), .rdata(f2274_rdata));
  assign f2274_clk = clk;
  assign f2274_rst = rst;
  // Bindings to f2274

  // f2276
  logic [0:0] f2276_wen;
  logic [31:0] f2276_wdata;
  logic [0:0] f2276_clk;
  logic [0:0] f2276_rst;
  logic [31:0] f2276_rdata;
  sr_buffer_32_1 f2276(.wen(f2276_wen), .wdata(f2276_wdata), .clk(f2276_clk), .rst(f2276_rst), .rdata(f2276_rdata));
  assign f2276_clk = clk;
  assign f2276_rst = rst;
  // Bindings to f2276

  // f2278
  logic [0:0] f2278_wen;
  logic [31:0] f2278_wdata;
  logic [0:0] f2278_clk;
  logic [0:0] f2278_rst;
  logic [31:0] f2278_rdata;
  sr_buffer_32_1 f2278(.wen(f2278_wen), .wdata(f2278_wdata), .clk(f2278_clk), .rst(f2278_rst), .rdata(f2278_rdata));
  assign f2278_clk = clk;
  assign f2278_rst = rst;
  // Bindings to f2278

  // f2280
  logic [0:0] f2280_wen;
  logic [31:0] f2280_wdata;
  logic [0:0] f2280_clk;
  logic [0:0] f2280_rst;
  logic [31:0] f2280_rdata;
  sr_buffer_32_1 f2280(.wen(f2280_wen), .wdata(f2280_wdata), .clk(f2280_clk), .rst(f2280_rst), .rdata(f2280_rdata));
  assign f2280_clk = clk;
  assign f2280_rst = rst;
  // Bindings to f2280

  // f2282
  logic [0:0] f2282_wen;
  logic [31:0] f2282_wdata;
  logic [0:0] f2282_clk;
  logic [0:0] f2282_rst;
  logic [31:0] f2282_rdata;
  sr_buffer_32_1 f2282(.wen(f2282_wen), .wdata(f2282_wdata), .clk(f2282_clk), .rst(f2282_rst), .rdata(f2282_rdata));
  assign f2282_clk = clk;
  assign f2282_rst = rst;
  // Bindings to f2282

  // f2284
  logic [0:0] f2284_wen;
  logic [31:0] f2284_wdata;
  logic [0:0] f2284_clk;
  logic [0:0] f2284_rst;
  logic [31:0] f2284_rdata;
  sr_buffer_32_1 f2284(.wen(f2284_wen), .wdata(f2284_wdata), .clk(f2284_clk), .rst(f2284_rst), .rdata(f2284_rdata));
  assign f2284_clk = clk;
  assign f2284_rst = rst;
  // Bindings to f2284

  // f2286
  logic [0:0] f2286_wen;
  logic [31:0] f2286_wdata;
  logic [0:0] f2286_clk;
  logic [0:0] f2286_rst;
  logic [31:0] f2286_rdata;
  sr_buffer_32_1 f2286(.wen(f2286_wen), .wdata(f2286_wdata), .clk(f2286_clk), .rst(f2286_rst), .rdata(f2286_rdata));
  assign f2286_clk = clk;
  assign f2286_rst = rst;
  // Bindings to f2286

  // f2288
  logic [0:0] f2288_wen;
  logic [31:0] f2288_wdata;
  logic [0:0] f2288_clk;
  logic [0:0] f2288_rst;
  logic [31:0] f2288_rdata;
  sr_buffer_32_1 f2288(.wen(f2288_wen), .wdata(f2288_wdata), .clk(f2288_clk), .rst(f2288_rst), .rdata(f2288_rdata));
  assign f2288_clk = clk;
  assign f2288_rst = rst;
  // Bindings to f2288

  // f2290
  logic [0:0] f2290_wen;
  logic [31:0] f2290_wdata;
  logic [0:0] f2290_clk;
  logic [0:0] f2290_rst;
  logic [31:0] f2290_rdata;
  sr_buffer_32_1 f2290(.wen(f2290_wen), .wdata(f2290_wdata), .clk(f2290_clk), .rst(f2290_rst), .rdata(f2290_rdata));
  assign f2290_clk = clk;
  assign f2290_rst = rst;
  // Bindings to f2290

  // f2292
  logic [0:0] f2292_wen;
  logic [31:0] f2292_wdata;
  logic [0:0] f2292_clk;
  logic [0:0] f2292_rst;
  logic [31:0] f2292_rdata;
  sr_buffer_32_1 f2292(.wen(f2292_wen), .wdata(f2292_wdata), .clk(f2292_clk), .rst(f2292_rst), .rdata(f2292_rdata));
  assign f2292_clk = clk;
  assign f2292_rst = rst;
  // Bindings to f2292

  // f2294
  logic [0:0] f2294_wen;
  logic [31:0] f2294_wdata;
  logic [0:0] f2294_clk;
  logic [0:0] f2294_rst;
  logic [31:0] f2294_rdata;
  sr_buffer_32_1 f2294(.wen(f2294_wen), .wdata(f2294_wdata), .clk(f2294_clk), .rst(f2294_rst), .rdata(f2294_rdata));
  assign f2294_clk = clk;
  assign f2294_rst = rst;
  // Bindings to f2294

  // f2296
  logic [0:0] f2296_wen;
  logic [31:0] f2296_wdata;
  logic [0:0] f2296_clk;
  logic [0:0] f2296_rst;
  logic [31:0] f2296_rdata;
  sr_buffer_32_1 f2296(.wen(f2296_wen), .wdata(f2296_wdata), .clk(f2296_clk), .rst(f2296_rst), .rdata(f2296_rdata));
  assign f2296_clk = clk;
  assign f2296_rst = rst;
  // Bindings to f2296

  // f2298
  logic [0:0] f2298_wen;
  logic [31:0] f2298_wdata;
  logic [0:0] f2298_clk;
  logic [0:0] f2298_rst;
  logic [31:0] f2298_rdata;
  sr_buffer_32_1 f2298(.wen(f2298_wen), .wdata(f2298_wdata), .clk(f2298_clk), .rst(f2298_rst), .rdata(f2298_rdata));
  assign f2298_clk = clk;
  assign f2298_rst = rst;
  // Bindings to f2298

  // f2300
  logic [0:0] f2300_wen;
  logic [31:0] f2300_wdata;
  logic [0:0] f2300_clk;
  logic [0:0] f2300_rst;
  logic [31:0] f2300_rdata;
  sr_buffer_32_1 f2300(.wen(f2300_wen), .wdata(f2300_wdata), .clk(f2300_clk), .rst(f2300_rst), .rdata(f2300_rdata));
  assign f2300_clk = clk;
  assign f2300_rst = rst;
  // Bindings to f2300

  // f2302
  logic [0:0] f2302_wen;
  logic [31:0] f2302_wdata;
  logic [0:0] f2302_clk;
  logic [0:0] f2302_rst;
  logic [31:0] f2302_rdata;
  sr_buffer_32_1 f2302(.wen(f2302_wen), .wdata(f2302_wdata), .clk(f2302_clk), .rst(f2302_rst), .rdata(f2302_rdata));
  assign f2302_clk = clk;
  assign f2302_rst = rst;
  // Bindings to f2302

  // f2304
  logic [0:0] f2304_wen;
  logic [31:0] f2304_wdata;
  logic [0:0] f2304_clk;
  logic [0:0] f2304_rst;
  logic [31:0] f2304_rdata;
  sr_buffer_32_1 f2304(.wen(f2304_wen), .wdata(f2304_wdata), .clk(f2304_clk), .rst(f2304_rst), .rdata(f2304_rdata));
  assign f2304_clk = clk;
  assign f2304_rst = rst;
  // Bindings to f2304

  // f2306
  logic [0:0] f2306_wen;
  logic [31:0] f2306_wdata;
  logic [0:0] f2306_clk;
  logic [0:0] f2306_rst;
  logic [31:0] f2306_rdata;
  sr_buffer_32_1 f2306(.wen(f2306_wen), .wdata(f2306_wdata), .clk(f2306_clk), .rst(f2306_rst), .rdata(f2306_rdata));
  assign f2306_clk = clk;
  assign f2306_rst = rst;
  // Bindings to f2306

  // f2308
  logic [0:0] f2308_wen;
  logic [31:0] f2308_wdata;
  logic [0:0] f2308_clk;
  logic [0:0] f2308_rst;
  logic [31:0] f2308_rdata;
  sr_buffer_32_1 f2308(.wen(f2308_wen), .wdata(f2308_wdata), .clk(f2308_clk), .rst(f2308_rst), .rdata(f2308_rdata));
  assign f2308_clk = clk;
  assign f2308_rst = rst;
  // Bindings to f2308

  // f2310
  logic [0:0] f2310_wen;
  logic [31:0] f2310_wdata;
  logic [0:0] f2310_clk;
  logic [0:0] f2310_rst;
  logic [31:0] f2310_rdata;
  sr_buffer_32_1 f2310(.wen(f2310_wen), .wdata(f2310_wdata), .clk(f2310_clk), .rst(f2310_rst), .rdata(f2310_rdata));
  assign f2310_clk = clk;
  assign f2310_rst = rst;
  // Bindings to f2310

  // f2312
  logic [0:0] f2312_wen;
  logic [31:0] f2312_wdata;
  logic [0:0] f2312_clk;
  logic [0:0] f2312_rst;
  logic [31:0] f2312_rdata;
  sr_buffer_32_1 f2312(.wen(f2312_wen), .wdata(f2312_wdata), .clk(f2312_clk), .rst(f2312_rst), .rdata(f2312_rdata));
  assign f2312_clk = clk;
  assign f2312_rst = rst;
  // Bindings to f2312

  // f2314
  logic [0:0] f2314_wen;
  logic [31:0] f2314_wdata;
  logic [0:0] f2314_clk;
  logic [0:0] f2314_rst;
  logic [31:0] f2314_rdata;
  sr_buffer_32_1 f2314(.wen(f2314_wen), .wdata(f2314_wdata), .clk(f2314_clk), .rst(f2314_rst), .rdata(f2314_rdata));
  assign f2314_clk = clk;
  assign f2314_rst = rst;
  // Bindings to f2314

  // f2316
  logic [0:0] f2316_wen;
  logic [31:0] f2316_wdata;
  logic [0:0] f2316_clk;
  logic [0:0] f2316_rst;
  logic [31:0] f2316_rdata;
  sr_buffer_32_1 f2316(.wen(f2316_wen), .wdata(f2316_wdata), .clk(f2316_clk), .rst(f2316_rst), .rdata(f2316_rdata));
  assign f2316_clk = clk;
  assign f2316_rst = rst;
  // Bindings to f2316

  // f2318
  logic [0:0] f2318_wen;
  logic [31:0] f2318_wdata;
  logic [0:0] f2318_clk;
  logic [0:0] f2318_rst;
  logic [31:0] f2318_rdata;
  sr_buffer_32_1 f2318(.wen(f2318_wen), .wdata(f2318_wdata), .clk(f2318_clk), .rst(f2318_rst), .rdata(f2318_rdata));
  assign f2318_clk = clk;
  assign f2318_rst = rst;
  // Bindings to f2318

  // f2320
  logic [0:0] f2320_wen;
  logic [31:0] f2320_wdata;
  logic [0:0] f2320_clk;
  logic [0:0] f2320_rst;
  logic [31:0] f2320_rdata;
  sr_buffer_32_1 f2320(.wen(f2320_wen), .wdata(f2320_wdata), .clk(f2320_clk), .rst(f2320_rst), .rdata(f2320_rdata));
  assign f2320_clk = clk;
  assign f2320_rst = rst;
  // Bindings to f2320

  // f2322
  logic [0:0] f2322_wen;
  logic [31:0] f2322_wdata;
  logic [0:0] f2322_clk;
  logic [0:0] f2322_rst;
  logic [31:0] f2322_rdata;
  sr_buffer_32_1 f2322(.wen(f2322_wen), .wdata(f2322_wdata), .clk(f2322_clk), .rst(f2322_rst), .rdata(f2322_rdata));
  assign f2322_clk = clk;
  assign f2322_rst = rst;
  // Bindings to f2322

  // f2324
  logic [0:0] f2324_wen;
  logic [31:0] f2324_wdata;
  logic [0:0] f2324_clk;
  logic [0:0] f2324_rst;
  logic [31:0] f2324_rdata;
  sr_buffer_32_1 f2324(.wen(f2324_wen), .wdata(f2324_wdata), .clk(f2324_clk), .rst(f2324_rst), .rdata(f2324_rdata));
  assign f2324_clk = clk;
  assign f2324_rst = rst;
  // Bindings to f2324

  // f2326
  logic [0:0] f2326_wen;
  logic [31:0] f2326_wdata;
  logic [0:0] f2326_clk;
  logic [0:0] f2326_rst;
  logic [31:0] f2326_rdata;
  sr_buffer_32_1 f2326(.wen(f2326_wen), .wdata(f2326_wdata), .clk(f2326_clk), .rst(f2326_rst), .rdata(f2326_rdata));
  assign f2326_clk = clk;
  assign f2326_rst = rst;
  // Bindings to f2326

  // f2328
  logic [0:0] f2328_wen;
  logic [31:0] f2328_wdata;
  logic [0:0] f2328_clk;
  logic [0:0] f2328_rst;
  logic [31:0] f2328_rdata;
  sr_buffer_32_1 f2328(.wen(f2328_wen), .wdata(f2328_wdata), .clk(f2328_clk), .rst(f2328_rst), .rdata(f2328_rdata));
  assign f2328_clk = clk;
  assign f2328_rst = rst;
  // Bindings to f2328

  // f2330
  logic [0:0] f2330_wen;
  logic [31:0] f2330_wdata;
  logic [0:0] f2330_clk;
  logic [0:0] f2330_rst;
  logic [31:0] f2330_rdata;
  sr_buffer_32_1 f2330(.wen(f2330_wen), .wdata(f2330_wdata), .clk(f2330_clk), .rst(f2330_rst), .rdata(f2330_rdata));
  assign f2330_clk = clk;
  assign f2330_rst = rst;
  // Bindings to f2330

  // f2332
  logic [0:0] f2332_wen;
  logic [31:0] f2332_wdata;
  logic [0:0] f2332_clk;
  logic [0:0] f2332_rst;
  logic [31:0] f2332_rdata;
  sr_buffer_32_1 f2332(.wen(f2332_wen), .wdata(f2332_wdata), .clk(f2332_clk), .rst(f2332_rst), .rdata(f2332_rdata));
  assign f2332_clk = clk;
  assign f2332_rst = rst;
  // Bindings to f2332

  // f2334
  logic [0:0] f2334_wen;
  logic [31:0] f2334_wdata;
  logic [0:0] f2334_clk;
  logic [0:0] f2334_rst;
  logic [31:0] f2334_rdata;
  sr_buffer_32_1 f2334(.wen(f2334_wen), .wdata(f2334_wdata), .clk(f2334_clk), .rst(f2334_rst), .rdata(f2334_rdata));
  assign f2334_clk = clk;
  assign f2334_rst = rst;
  // Bindings to f2334

  // f2336
  logic [0:0] f2336_wen;
  logic [31:0] f2336_wdata;
  logic [0:0] f2336_clk;
  logic [0:0] f2336_rst;
  logic [31:0] f2336_rdata;
  sr_buffer_32_1 f2336(.wen(f2336_wen), .wdata(f2336_wdata), .clk(f2336_clk), .rst(f2336_rst), .rdata(f2336_rdata));
  assign f2336_clk = clk;
  assign f2336_rst = rst;
  // Bindings to f2336

  // f2338
  logic [0:0] f2338_wen;
  logic [31:0] f2338_wdata;
  logic [0:0] f2338_clk;
  logic [0:0] f2338_rst;
  logic [31:0] f2338_rdata;
  sr_buffer_32_1 f2338(.wen(f2338_wen), .wdata(f2338_wdata), .clk(f2338_clk), .rst(f2338_rst), .rdata(f2338_rdata));
  assign f2338_clk = clk;
  assign f2338_rst = rst;
  // Bindings to f2338

  // f2340
  logic [0:0] f2340_wen;
  logic [31:0] f2340_wdata;
  logic [0:0] f2340_clk;
  logic [0:0] f2340_rst;
  logic [31:0] f2340_rdata;
  sr_buffer_32_1 f2340(.wen(f2340_wen), .wdata(f2340_wdata), .clk(f2340_clk), .rst(f2340_rst), .rdata(f2340_rdata));
  assign f2340_clk = clk;
  assign f2340_rst = rst;
  // Bindings to f2340

  // f2342
  logic [0:0] f2342_wen;
  logic [31:0] f2342_wdata;
  logic [0:0] f2342_clk;
  logic [0:0] f2342_rst;
  logic [31:0] f2342_rdata;
  sr_buffer_32_1 f2342(.wen(f2342_wen), .wdata(f2342_wdata), .clk(f2342_clk), .rst(f2342_rst), .rdata(f2342_rdata));
  assign f2342_clk = clk;
  assign f2342_rst = rst;
  // Bindings to f2342

  // f2344
  logic [0:0] f2344_wen;
  logic [31:0] f2344_wdata;
  logic [0:0] f2344_clk;
  logic [0:0] f2344_rst;
  logic [31:0] f2344_rdata;
  sr_buffer_32_1 f2344(.wen(f2344_wen), .wdata(f2344_wdata), .clk(f2344_clk), .rst(f2344_rst), .rdata(f2344_rdata));
  assign f2344_clk = clk;
  assign f2344_rst = rst;
  // Bindings to f2344

  // f2346
  logic [0:0] f2346_wen;
  logic [31:0] f2346_wdata;
  logic [0:0] f2346_clk;
  logic [0:0] f2346_rst;
  logic [31:0] f2346_rdata;
  sr_buffer_32_1 f2346(.wen(f2346_wen), .wdata(f2346_wdata), .clk(f2346_clk), .rst(f2346_rst), .rdata(f2346_rdata));
  assign f2346_clk = clk;
  assign f2346_rst = rst;
  // Bindings to f2346

  // f2348
  logic [0:0] f2348_wen;
  logic [31:0] f2348_wdata;
  logic [0:0] f2348_clk;
  logic [0:0] f2348_rst;
  logic [31:0] f2348_rdata;
  sr_buffer_32_1 f2348(.wen(f2348_wen), .wdata(f2348_wdata), .clk(f2348_clk), .rst(f2348_rst), .rdata(f2348_rdata));
  assign f2348_clk = clk;
  assign f2348_rst = rst;
  // Bindings to f2348

  // f2350
  logic [0:0] f2350_wen;
  logic [31:0] f2350_wdata;
  logic [0:0] f2350_clk;
  logic [0:0] f2350_rst;
  logic [31:0] f2350_rdata;
  sr_buffer_32_1 f2350(.wen(f2350_wen), .wdata(f2350_wdata), .clk(f2350_clk), .rst(f2350_rst), .rdata(f2350_rdata));
  assign f2350_clk = clk;
  assign f2350_rst = rst;
  // Bindings to f2350

  // f2352
  logic [0:0] f2352_wen;
  logic [31:0] f2352_wdata;
  logic [0:0] f2352_clk;
  logic [0:0] f2352_rst;
  logic [31:0] f2352_rdata;
  sr_buffer_32_1 f2352(.wen(f2352_wen), .wdata(f2352_wdata), .clk(f2352_clk), .rst(f2352_rst), .rdata(f2352_rdata));
  assign f2352_clk = clk;
  assign f2352_rst = rst;
  // Bindings to f2352

  // f2354
  logic [0:0] f2354_wen;
  logic [31:0] f2354_wdata;
  logic [0:0] f2354_clk;
  logic [0:0] f2354_rst;
  logic [31:0] f2354_rdata;
  sr_buffer_32_1 f2354(.wen(f2354_wen), .wdata(f2354_wdata), .clk(f2354_clk), .rst(f2354_rst), .rdata(f2354_rdata));
  assign f2354_clk = clk;
  assign f2354_rst = rst;
  // Bindings to f2354

  // f2356
  logic [0:0] f2356_wen;
  logic [31:0] f2356_wdata;
  logic [0:0] f2356_clk;
  logic [0:0] f2356_rst;
  logic [31:0] f2356_rdata;
  sr_buffer_32_1 f2356(.wen(f2356_wen), .wdata(f2356_wdata), .clk(f2356_clk), .rst(f2356_rst), .rdata(f2356_rdata));
  assign f2356_clk = clk;
  assign f2356_rst = rst;
  // Bindings to f2356

  // f2358
  logic [0:0] f2358_wen;
  logic [31:0] f2358_wdata;
  logic [0:0] f2358_clk;
  logic [0:0] f2358_rst;
  logic [31:0] f2358_rdata;
  sr_buffer_32_1 f2358(.wen(f2358_wen), .wdata(f2358_wdata), .clk(f2358_clk), .rst(f2358_rst), .rdata(f2358_rdata));
  assign f2358_clk = clk;
  assign f2358_rst = rst;
  // Bindings to f2358

  // f2360
  logic [0:0] f2360_wen;
  logic [31:0] f2360_wdata;
  logic [0:0] f2360_clk;
  logic [0:0] f2360_rst;
  logic [31:0] f2360_rdata;
  sr_buffer_32_1 f2360(.wen(f2360_wen), .wdata(f2360_wdata), .clk(f2360_clk), .rst(f2360_rst), .rdata(f2360_rdata));
  assign f2360_clk = clk;
  assign f2360_rst = rst;
  // Bindings to f2360

  // f2362
  logic [0:0] f2362_wen;
  logic [31:0] f2362_wdata;
  logic [0:0] f2362_clk;
  logic [0:0] f2362_rst;
  logic [31:0] f2362_rdata;
  sr_buffer_32_1 f2362(.wen(f2362_wen), .wdata(f2362_wdata), .clk(f2362_clk), .rst(f2362_rst), .rdata(f2362_rdata));
  assign f2362_clk = clk;
  assign f2362_rst = rst;
  // Bindings to f2362

  // f2364
  logic [0:0] f2364_wen;
  logic [31:0] f2364_wdata;
  logic [0:0] f2364_clk;
  logic [0:0] f2364_rst;
  logic [31:0] f2364_rdata;
  sr_buffer_32_1 f2364(.wen(f2364_wen), .wdata(f2364_wdata), .clk(f2364_clk), .rst(f2364_rst), .rdata(f2364_rdata));
  assign f2364_clk = clk;
  assign f2364_rst = rst;
  // Bindings to f2364

  // f2366
  logic [0:0] f2366_wen;
  logic [31:0] f2366_wdata;
  logic [0:0] f2366_clk;
  logic [0:0] f2366_rst;
  logic [31:0] f2366_rdata;
  sr_buffer_32_1 f2366(.wen(f2366_wen), .wdata(f2366_wdata), .clk(f2366_clk), .rst(f2366_rst), .rdata(f2366_rdata));
  assign f2366_clk = clk;
  assign f2366_rst = rst;
  // Bindings to f2366

  // f2368
  logic [0:0] f2368_wen;
  logic [31:0] f2368_wdata;
  logic [0:0] f2368_clk;
  logic [0:0] f2368_rst;
  logic [31:0] f2368_rdata;
  sr_buffer_32_1 f2368(.wen(f2368_wen), .wdata(f2368_wdata), .clk(f2368_clk), .rst(f2368_rst), .rdata(f2368_rdata));
  assign f2368_clk = clk;
  assign f2368_rst = rst;
  // Bindings to f2368

  // f2370
  logic [0:0] f2370_wen;
  logic [31:0] f2370_wdata;
  logic [0:0] f2370_clk;
  logic [0:0] f2370_rst;
  logic [31:0] f2370_rdata;
  sr_buffer_32_1 f2370(.wen(f2370_wen), .wdata(f2370_wdata), .clk(f2370_clk), .rst(f2370_rst), .rdata(f2370_rdata));
  assign f2370_clk = clk;
  assign f2370_rst = rst;
  // Bindings to f2370

  // f2372
  logic [0:0] f2372_wen;
  logic [31:0] f2372_wdata;
  logic [0:0] f2372_clk;
  logic [0:0] f2372_rst;
  logic [31:0] f2372_rdata;
  sr_buffer_32_1 f2372(.wen(f2372_wen), .wdata(f2372_wdata), .clk(f2372_clk), .rst(f2372_rst), .rdata(f2372_rdata));
  assign f2372_clk = clk;
  assign f2372_rst = rst;
  // Bindings to f2372

  // f2374
  logic [0:0] f2374_wen;
  logic [31:0] f2374_wdata;
  logic [0:0] f2374_clk;
  logic [0:0] f2374_rst;
  logic [31:0] f2374_rdata;
  sr_buffer_32_1 f2374(.wen(f2374_wen), .wdata(f2374_wdata), .clk(f2374_clk), .rst(f2374_rst), .rdata(f2374_rdata));
  assign f2374_clk = clk;
  assign f2374_rst = rst;
  // Bindings to f2374

  // f2376
  logic [0:0] f2376_wen;
  logic [31:0] f2376_wdata;
  logic [0:0] f2376_clk;
  logic [0:0] f2376_rst;
  logic [31:0] f2376_rdata;
  sr_buffer_32_1 f2376(.wen(f2376_wen), .wdata(f2376_wdata), .clk(f2376_clk), .rst(f2376_rst), .rdata(f2376_rdata));
  assign f2376_clk = clk;
  assign f2376_rst = rst;
  // Bindings to f2376

  // f2378
  logic [0:0] f2378_wen;
  logic [31:0] f2378_wdata;
  logic [0:0] f2378_clk;
  logic [0:0] f2378_rst;
  logic [31:0] f2378_rdata;
  sr_buffer_32_1 f2378(.wen(f2378_wen), .wdata(f2378_wdata), .clk(f2378_clk), .rst(f2378_rst), .rdata(f2378_rdata));
  assign f2378_clk = clk;
  assign f2378_rst = rst;
  // Bindings to f2378

  // f2380
  logic [0:0] f2380_wen;
  logic [31:0] f2380_wdata;
  logic [0:0] f2380_clk;
  logic [0:0] f2380_rst;
  logic [31:0] f2380_rdata;
  sr_buffer_32_1 f2380(.wen(f2380_wen), .wdata(f2380_wdata), .clk(f2380_clk), .rst(f2380_rst), .rdata(f2380_rdata));
  assign f2380_clk = clk;
  assign f2380_rst = rst;
  // Bindings to f2380

  // f2382
  logic [0:0] f2382_wen;
  logic [31:0] f2382_wdata;
  logic [0:0] f2382_clk;
  logic [0:0] f2382_rst;
  logic [31:0] f2382_rdata;
  sr_buffer_32_1 f2382(.wen(f2382_wen), .wdata(f2382_wdata), .clk(f2382_clk), .rst(f2382_rst), .rdata(f2382_rdata));
  assign f2382_clk = clk;
  assign f2382_rst = rst;
  // Bindings to f2382

  // f2384
  logic [0:0] f2384_wen;
  logic [31:0] f2384_wdata;
  logic [0:0] f2384_clk;
  logic [0:0] f2384_rst;
  logic [31:0] f2384_rdata;
  sr_buffer_32_1 f2384(.wen(f2384_wen), .wdata(f2384_wdata), .clk(f2384_clk), .rst(f2384_rst), .rdata(f2384_rdata));
  assign f2384_clk = clk;
  assign f2384_rst = rst;
  // Bindings to f2384

  // f2386
  logic [0:0] f2386_wen;
  logic [31:0] f2386_wdata;
  logic [0:0] f2386_clk;
  logic [0:0] f2386_rst;
  logic [31:0] f2386_rdata;
  sr_buffer_32_1 f2386(.wen(f2386_wen), .wdata(f2386_wdata), .clk(f2386_clk), .rst(f2386_rst), .rdata(f2386_rdata));
  assign f2386_clk = clk;
  assign f2386_rst = rst;
  // Bindings to f2386

  // f2388
  logic [0:0] f2388_wen;
  logic [31:0] f2388_wdata;
  logic [0:0] f2388_clk;
  logic [0:0] f2388_rst;
  logic [31:0] f2388_rdata;
  sr_buffer_32_1 f2388(.wen(f2388_wen), .wdata(f2388_wdata), .clk(f2388_clk), .rst(f2388_rst), .rdata(f2388_rdata));
  assign f2388_clk = clk;
  assign f2388_rst = rst;
  // Bindings to f2388

  // f2390
  logic [0:0] f2390_wen;
  logic [31:0] f2390_wdata;
  logic [0:0] f2390_clk;
  logic [0:0] f2390_rst;
  logic [31:0] f2390_rdata;
  sr_buffer_32_1 f2390(.wen(f2390_wen), .wdata(f2390_wdata), .clk(f2390_clk), .rst(f2390_rst), .rdata(f2390_rdata));
  assign f2390_clk = clk;
  assign f2390_rst = rst;
  // Bindings to f2390

  // f2392
  logic [0:0] f2392_wen;
  logic [31:0] f2392_wdata;
  logic [0:0] f2392_clk;
  logic [0:0] f2392_rst;
  logic [31:0] f2392_rdata;
  sr_buffer_32_1 f2392(.wen(f2392_wen), .wdata(f2392_wdata), .clk(f2392_clk), .rst(f2392_rst), .rdata(f2392_rdata));
  assign f2392_clk = clk;
  assign f2392_rst = rst;
  // Bindings to f2392

  // f2394
  logic [0:0] f2394_wen;
  logic [31:0] f2394_wdata;
  logic [0:0] f2394_clk;
  logic [0:0] f2394_rst;
  logic [31:0] f2394_rdata;
  sr_buffer_32_1 f2394(.wen(f2394_wen), .wdata(f2394_wdata), .clk(f2394_clk), .rst(f2394_rst), .rdata(f2394_rdata));
  assign f2394_clk = clk;
  assign f2394_rst = rst;
  // Bindings to f2394

  // f2396
  logic [0:0] f2396_wen;
  logic [31:0] f2396_wdata;
  logic [0:0] f2396_clk;
  logic [0:0] f2396_rst;
  logic [31:0] f2396_rdata;
  sr_buffer_32_1 f2396(.wen(f2396_wen), .wdata(f2396_wdata), .clk(f2396_clk), .rst(f2396_rst), .rdata(f2396_rdata));
  assign f2396_clk = clk;
  assign f2396_rst = rst;
  // Bindings to f2396

  // f2398
  logic [0:0] f2398_wen;
  logic [31:0] f2398_wdata;
  logic [0:0] f2398_clk;
  logic [0:0] f2398_rst;
  logic [31:0] f2398_rdata;
  sr_buffer_32_1 f2398(.wen(f2398_wen), .wdata(f2398_wdata), .clk(f2398_clk), .rst(f2398_rst), .rdata(f2398_rdata));
  assign f2398_clk = clk;
  assign f2398_rst = rst;
  // Bindings to f2398

  // f2400
  logic [0:0] f2400_wen;
  logic [31:0] f2400_wdata;
  logic [0:0] f2400_clk;
  logic [0:0] f2400_rst;
  logic [31:0] f2400_rdata;
  sr_buffer_32_1 f2400(.wen(f2400_wen), .wdata(f2400_wdata), .clk(f2400_clk), .rst(f2400_rst), .rdata(f2400_rdata));
  assign f2400_clk = clk;
  assign f2400_rst = rst;
  // Bindings to f2400

  // f2402
  logic [0:0] f2402_wen;
  logic [31:0] f2402_wdata;
  logic [0:0] f2402_clk;
  logic [0:0] f2402_rst;
  logic [31:0] f2402_rdata;
  sr_buffer_32_1 f2402(.wen(f2402_wen), .wdata(f2402_wdata), .clk(f2402_clk), .rst(f2402_rst), .rdata(f2402_rdata));
  assign f2402_clk = clk;
  assign f2402_rst = rst;
  // Bindings to f2402

  // f2404
  logic [0:0] f2404_wen;
  logic [31:0] f2404_wdata;
  logic [0:0] f2404_clk;
  logic [0:0] f2404_rst;
  logic [31:0] f2404_rdata;
  sr_buffer_32_1 f2404(.wen(f2404_wen), .wdata(f2404_wdata), .clk(f2404_clk), .rst(f2404_rst), .rdata(f2404_rdata));
  assign f2404_clk = clk;
  assign f2404_rst = rst;
  // Bindings to f2404

  // f2406
  logic [0:0] f2406_wen;
  logic [31:0] f2406_wdata;
  logic [0:0] f2406_clk;
  logic [0:0] f2406_rst;
  logic [31:0] f2406_rdata;
  sr_buffer_32_1 f2406(.wen(f2406_wen), .wdata(f2406_wdata), .clk(f2406_clk), .rst(f2406_rst), .rdata(f2406_rdata));
  assign f2406_clk = clk;
  assign f2406_rst = rst;
  // Bindings to f2406

  // f2408
  logic [0:0] f2408_wen;
  logic [31:0] f2408_wdata;
  logic [0:0] f2408_clk;
  logic [0:0] f2408_rst;
  logic [31:0] f2408_rdata;
  sr_buffer_32_1 f2408(.wen(f2408_wen), .wdata(f2408_wdata), .clk(f2408_clk), .rst(f2408_rst), .rdata(f2408_rdata));
  assign f2408_clk = clk;
  assign f2408_rst = rst;
  // Bindings to f2408

  // f2410
  logic [0:0] f2410_wen;
  logic [31:0] f2410_wdata;
  logic [0:0] f2410_clk;
  logic [0:0] f2410_rst;
  logic [31:0] f2410_rdata;
  sr_buffer_32_1 f2410(.wen(f2410_wen), .wdata(f2410_wdata), .clk(f2410_clk), .rst(f2410_rst), .rdata(f2410_rdata));
  assign f2410_clk = clk;
  assign f2410_rst = rst;
  // Bindings to f2410

  // f2412
  logic [0:0] f2412_wen;
  logic [31:0] f2412_wdata;
  logic [0:0] f2412_clk;
  logic [0:0] f2412_rst;
  logic [31:0] f2412_rdata;
  sr_buffer_32_1 f2412(.wen(f2412_wen), .wdata(f2412_wdata), .clk(f2412_clk), .rst(f2412_rst), .rdata(f2412_rdata));
  assign f2412_clk = clk;
  assign f2412_rst = rst;
  // Bindings to f2412

  // f2414
  logic [0:0] f2414_wen;
  logic [31:0] f2414_wdata;
  logic [0:0] f2414_clk;
  logic [0:0] f2414_rst;
  logic [31:0] f2414_rdata;
  sr_buffer_32_1 f2414(.wen(f2414_wen), .wdata(f2414_wdata), .clk(f2414_clk), .rst(f2414_rst), .rdata(f2414_rdata));
  assign f2414_clk = clk;
  assign f2414_rst = rst;
  // Bindings to f2414

  // f2416
  logic [0:0] f2416_wen;
  logic [31:0] f2416_wdata;
  logic [0:0] f2416_clk;
  logic [0:0] f2416_rst;
  logic [31:0] f2416_rdata;
  sr_buffer_32_1 f2416(.wen(f2416_wen), .wdata(f2416_wdata), .clk(f2416_clk), .rst(f2416_rst), .rdata(f2416_rdata));
  assign f2416_clk = clk;
  assign f2416_rst = rst;
  // Bindings to f2416

  // f2418
  logic [0:0] f2418_wen;
  logic [31:0] f2418_wdata;
  logic [0:0] f2418_clk;
  logic [0:0] f2418_rst;
  logic [31:0] f2418_rdata;
  sr_buffer_32_1 f2418(.wen(f2418_wen), .wdata(f2418_wdata), .clk(f2418_clk), .rst(f2418_rst), .rdata(f2418_rdata));
  assign f2418_clk = clk;
  assign f2418_rst = rst;
  // Bindings to f2418

  // f2420
  logic [0:0] f2420_wen;
  logic [31:0] f2420_wdata;
  logic [0:0] f2420_clk;
  logic [0:0] f2420_rst;
  logic [31:0] f2420_rdata;
  sr_buffer_32_1 f2420(.wen(f2420_wen), .wdata(f2420_wdata), .clk(f2420_clk), .rst(f2420_rst), .rdata(f2420_rdata));
  assign f2420_clk = clk;
  assign f2420_rst = rst;
  // Bindings to f2420

  // f2422
  logic [0:0] f2422_wen;
  logic [31:0] f2422_wdata;
  logic [0:0] f2422_clk;
  logic [0:0] f2422_rst;
  logic [31:0] f2422_rdata;
  sr_buffer_32_1 f2422(.wen(f2422_wen), .wdata(f2422_wdata), .clk(f2422_clk), .rst(f2422_rst), .rdata(f2422_rdata));
  assign f2422_clk = clk;
  assign f2422_rst = rst;
  // Bindings to f2422

  // f2424
  logic [0:0] f2424_wen;
  logic [31:0] f2424_wdata;
  logic [0:0] f2424_clk;
  logic [0:0] f2424_rst;
  logic [31:0] f2424_rdata;
  sr_buffer_32_1 f2424(.wen(f2424_wen), .wdata(f2424_wdata), .clk(f2424_clk), .rst(f2424_rst), .rdata(f2424_rdata));
  assign f2424_clk = clk;
  assign f2424_rst = rst;
  // Bindings to f2424

  // f2426
  logic [0:0] f2426_wen;
  logic [31:0] f2426_wdata;
  logic [0:0] f2426_clk;
  logic [0:0] f2426_rst;
  logic [31:0] f2426_rdata;
  sr_buffer_32_1 f2426(.wen(f2426_wen), .wdata(f2426_wdata), .clk(f2426_clk), .rst(f2426_rst), .rdata(f2426_rdata));
  assign f2426_clk = clk;
  assign f2426_rst = rst;
  // Bindings to f2426

  // f2428
  logic [0:0] f2428_wen;
  logic [31:0] f2428_wdata;
  logic [0:0] f2428_clk;
  logic [0:0] f2428_rst;
  logic [31:0] f2428_rdata;
  sr_buffer_32_1 f2428(.wen(f2428_wen), .wdata(f2428_wdata), .clk(f2428_clk), .rst(f2428_rst), .rdata(f2428_rdata));
  assign f2428_clk = clk;
  assign f2428_rst = rst;
  // Bindings to f2428

  // f2430
  logic [0:0] f2430_wen;
  logic [31:0] f2430_wdata;
  logic [0:0] f2430_clk;
  logic [0:0] f2430_rst;
  logic [31:0] f2430_rdata;
  sr_buffer_32_1 f2430(.wen(f2430_wen), .wdata(f2430_wdata), .clk(f2430_clk), .rst(f2430_rst), .rdata(f2430_rdata));
  assign f2430_clk = clk;
  assign f2430_rst = rst;
  // Bindings to f2430

  // f2432
  logic [0:0] f2432_wen;
  logic [31:0] f2432_wdata;
  logic [0:0] f2432_clk;
  logic [0:0] f2432_rst;
  logic [31:0] f2432_rdata;
  sr_buffer_32_1 f2432(.wen(f2432_wen), .wdata(f2432_wdata), .clk(f2432_clk), .rst(f2432_rst), .rdata(f2432_rdata));
  assign f2432_clk = clk;
  assign f2432_rst = rst;
  // Bindings to f2432

  // f2434
  logic [0:0] f2434_wen;
  logic [31:0] f2434_wdata;
  logic [0:0] f2434_clk;
  logic [0:0] f2434_rst;
  logic [31:0] f2434_rdata;
  sr_buffer_32_1 f2434(.wen(f2434_wen), .wdata(f2434_wdata), .clk(f2434_clk), .rst(f2434_rst), .rdata(f2434_rdata));
  assign f2434_clk = clk;
  assign f2434_rst = rst;
  // Bindings to f2434

  // f2436
  logic [0:0] f2436_wen;
  logic [31:0] f2436_wdata;
  logic [0:0] f2436_clk;
  logic [0:0] f2436_rst;
  logic [31:0] f2436_rdata;
  sr_buffer_32_1 f2436(.wen(f2436_wen), .wdata(f2436_wdata), .clk(f2436_clk), .rst(f2436_rst), .rdata(f2436_rdata));
  assign f2436_clk = clk;
  assign f2436_rst = rst;
  // Bindings to f2436

  // f2438
  logic [0:0] f2438_wen;
  logic [31:0] f2438_wdata;
  logic [0:0] f2438_clk;
  logic [0:0] f2438_rst;
  logic [31:0] f2438_rdata;
  sr_buffer_32_1 f2438(.wen(f2438_wen), .wdata(f2438_wdata), .clk(f2438_clk), .rst(f2438_rst), .rdata(f2438_rdata));
  assign f2438_clk = clk;
  assign f2438_rst = rst;
  // Bindings to f2438

  // f2440
  logic [0:0] f2440_wen;
  logic [31:0] f2440_wdata;
  logic [0:0] f2440_clk;
  logic [0:0] f2440_rst;
  logic [31:0] f2440_rdata;
  sr_buffer_32_1 f2440(.wen(f2440_wen), .wdata(f2440_wdata), .clk(f2440_clk), .rst(f2440_rst), .rdata(f2440_rdata));
  assign f2440_clk = clk;
  assign f2440_rst = rst;
  // Bindings to f2440

  // f2442
  logic [0:0] f2442_wen;
  logic [31:0] f2442_wdata;
  logic [0:0] f2442_clk;
  logic [0:0] f2442_rst;
  logic [31:0] f2442_rdata;
  sr_buffer_32_1 f2442(.wen(f2442_wen), .wdata(f2442_wdata), .clk(f2442_clk), .rst(f2442_rst), .rdata(f2442_rdata));
  assign f2442_clk = clk;
  assign f2442_rst = rst;
  // Bindings to f2442

  // f2444
  logic [0:0] f2444_wen;
  logic [31:0] f2444_wdata;
  logic [0:0] f2444_clk;
  logic [0:0] f2444_rst;
  logic [31:0] f2444_rdata;
  sr_buffer_32_1 f2444(.wen(f2444_wen), .wdata(f2444_wdata), .clk(f2444_clk), .rst(f2444_rst), .rdata(f2444_rdata));
  assign f2444_clk = clk;
  assign f2444_rst = rst;
  // Bindings to f2444

  // f2446
  logic [0:0] f2446_wen;
  logic [31:0] f2446_wdata;
  logic [0:0] f2446_clk;
  logic [0:0] f2446_rst;
  logic [31:0] f2446_rdata;
  sr_buffer_32_1 f2446(.wen(f2446_wen), .wdata(f2446_wdata), .clk(f2446_clk), .rst(f2446_rst), .rdata(f2446_rdata));
  assign f2446_clk = clk;
  assign f2446_rst = rst;
  // Bindings to f2446

  // f2448
  logic [0:0] f2448_wen;
  logic [31:0] f2448_wdata;
  logic [0:0] f2448_clk;
  logic [0:0] f2448_rst;
  logic [31:0] f2448_rdata;
  sr_buffer_32_1 f2448(.wen(f2448_wen), .wdata(f2448_wdata), .clk(f2448_clk), .rst(f2448_rst), .rdata(f2448_rdata));
  assign f2448_clk = clk;
  assign f2448_rst = rst;
  // Bindings to f2448

  // f2450
  logic [0:0] f2450_wen;
  logic [31:0] f2450_wdata;
  logic [0:0] f2450_clk;
  logic [0:0] f2450_rst;
  logic [31:0] f2450_rdata;
  sr_buffer_32_1 f2450(.wen(f2450_wen), .wdata(f2450_wdata), .clk(f2450_clk), .rst(f2450_rst), .rdata(f2450_rdata));
  assign f2450_clk = clk;
  assign f2450_rst = rst;
  // Bindings to f2450

  // f2452
  logic [0:0] f2452_wen;
  logic [31:0] f2452_wdata;
  logic [0:0] f2452_clk;
  logic [0:0] f2452_rst;
  logic [31:0] f2452_rdata;
  sr_buffer_32_1 f2452(.wen(f2452_wen), .wdata(f2452_wdata), .clk(f2452_clk), .rst(f2452_rst), .rdata(f2452_rdata));
  assign f2452_clk = clk;
  assign f2452_rst = rst;
  // Bindings to f2452

  // f2454
  logic [0:0] f2454_wen;
  logic [31:0] f2454_wdata;
  logic [0:0] f2454_clk;
  logic [0:0] f2454_rst;
  logic [31:0] f2454_rdata;
  sr_buffer_32_1 f2454(.wen(f2454_wen), .wdata(f2454_wdata), .clk(f2454_clk), .rst(f2454_rst), .rdata(f2454_rdata));
  assign f2454_clk = clk;
  assign f2454_rst = rst;
  // Bindings to f2454

  // f2456
  logic [0:0] f2456_wen;
  logic [31:0] f2456_wdata;
  logic [0:0] f2456_clk;
  logic [0:0] f2456_rst;
  logic [31:0] f2456_rdata;
  sr_buffer_32_1 f2456(.wen(f2456_wen), .wdata(f2456_wdata), .clk(f2456_clk), .rst(f2456_rst), .rdata(f2456_rdata));
  assign f2456_clk = clk;
  assign f2456_rst = rst;
  // Bindings to f2456

  // f2458
  logic [0:0] f2458_wen;
  logic [31:0] f2458_wdata;
  logic [0:0] f2458_clk;
  logic [0:0] f2458_rst;
  logic [31:0] f2458_rdata;
  sr_buffer_32_1 f2458(.wen(f2458_wen), .wdata(f2458_wdata), .clk(f2458_clk), .rst(f2458_rst), .rdata(f2458_rdata));
  assign f2458_clk = clk;
  assign f2458_rst = rst;
  // Bindings to f2458

  // f2460
  logic [0:0] f2460_wen;
  logic [31:0] f2460_wdata;
  logic [0:0] f2460_clk;
  logic [0:0] f2460_rst;
  logic [31:0] f2460_rdata;
  sr_buffer_32_1 f2460(.wen(f2460_wen), .wdata(f2460_wdata), .clk(f2460_clk), .rst(f2460_rst), .rdata(f2460_rdata));
  assign f2460_clk = clk;
  assign f2460_rst = rst;
  // Bindings to f2460

  // f2462
  logic [0:0] f2462_wen;
  logic [31:0] f2462_wdata;
  logic [0:0] f2462_clk;
  logic [0:0] f2462_rst;
  logic [31:0] f2462_rdata;
  sr_buffer_32_1 f2462(.wen(f2462_wen), .wdata(f2462_wdata), .clk(f2462_clk), .rst(f2462_rst), .rdata(f2462_rdata));
  assign f2462_clk = clk;
  assign f2462_rst = rst;
  // Bindings to f2462

  // f2464
  logic [0:0] f2464_wen;
  logic [31:0] f2464_wdata;
  logic [0:0] f2464_clk;
  logic [0:0] f2464_rst;
  logic [31:0] f2464_rdata;
  sr_buffer_32_1 f2464(.wen(f2464_wen), .wdata(f2464_wdata), .clk(f2464_clk), .rst(f2464_rst), .rdata(f2464_rdata));
  assign f2464_clk = clk;
  assign f2464_rst = rst;
  // Bindings to f2464

  // f2466
  logic [0:0] f2466_wen;
  logic [31:0] f2466_wdata;
  logic [0:0] f2466_clk;
  logic [0:0] f2466_rst;
  logic [31:0] f2466_rdata;
  sr_buffer_32_1 f2466(.wen(f2466_wen), .wdata(f2466_wdata), .clk(f2466_clk), .rst(f2466_rst), .rdata(f2466_rdata));
  assign f2466_clk = clk;
  assign f2466_rst = rst;
  // Bindings to f2466

  // f2468
  logic [0:0] f2468_wen;
  logic [31:0] f2468_wdata;
  logic [0:0] f2468_clk;
  logic [0:0] f2468_rst;
  logic [31:0] f2468_rdata;
  sr_buffer_32_1 f2468(.wen(f2468_wen), .wdata(f2468_wdata), .clk(f2468_clk), .rst(f2468_rst), .rdata(f2468_rdata));
  assign f2468_clk = clk;
  assign f2468_rst = rst;
  // Bindings to f2468

  // f2470
  logic [0:0] f2470_wen;
  logic [31:0] f2470_wdata;
  logic [0:0] f2470_clk;
  logic [0:0] f2470_rst;
  logic [31:0] f2470_rdata;
  sr_buffer_32_1 f2470(.wen(f2470_wen), .wdata(f2470_wdata), .clk(f2470_clk), .rst(f2470_rst), .rdata(f2470_rdata));
  assign f2470_clk = clk;
  assign f2470_rst = rst;
  // Bindings to f2470

  // f2472
  logic [0:0] f2472_wen;
  logic [31:0] f2472_wdata;
  logic [0:0] f2472_clk;
  logic [0:0] f2472_rst;
  logic [31:0] f2472_rdata;
  sr_buffer_32_1 f2472(.wen(f2472_wen), .wdata(f2472_wdata), .clk(f2472_clk), .rst(f2472_rst), .rdata(f2472_rdata));
  assign f2472_clk = clk;
  assign f2472_rst = rst;
  // Bindings to f2472

  // f2474
  logic [0:0] f2474_wen;
  logic [31:0] f2474_wdata;
  logic [0:0] f2474_clk;
  logic [0:0] f2474_rst;
  logic [31:0] f2474_rdata;
  sr_buffer_32_1 f2474(.wen(f2474_wen), .wdata(f2474_wdata), .clk(f2474_clk), .rst(f2474_rst), .rdata(f2474_rdata));
  assign f2474_clk = clk;
  assign f2474_rst = rst;
  // Bindings to f2474

  // f2476
  logic [0:0] f2476_wen;
  logic [31:0] f2476_wdata;
  logic [0:0] f2476_clk;
  logic [0:0] f2476_rst;
  logic [31:0] f2476_rdata;
  sr_buffer_32_1 f2476(.wen(f2476_wen), .wdata(f2476_wdata), .clk(f2476_clk), .rst(f2476_rst), .rdata(f2476_rdata));
  assign f2476_clk = clk;
  assign f2476_rst = rst;
  // Bindings to f2476

  // f2478
  logic [0:0] f2478_wen;
  logic [31:0] f2478_wdata;
  logic [0:0] f2478_clk;
  logic [0:0] f2478_rst;
  logic [31:0] f2478_rdata;
  sr_buffer_32_1 f2478(.wen(f2478_wen), .wdata(f2478_wdata), .clk(f2478_clk), .rst(f2478_rst), .rdata(f2478_rdata));
  assign f2478_clk = clk;
  assign f2478_rst = rst;
  // Bindings to f2478

  // f2480
  logic [0:0] f2480_wen;
  logic [31:0] f2480_wdata;
  logic [0:0] f2480_clk;
  logic [0:0] f2480_rst;
  logic [31:0] f2480_rdata;
  sr_buffer_32_1 f2480(.wen(f2480_wen), .wdata(f2480_wdata), .clk(f2480_clk), .rst(f2480_rst), .rdata(f2480_rdata));
  assign f2480_clk = clk;
  assign f2480_rst = rst;
  // Bindings to f2480

  // f2482
  logic [0:0] f2482_wen;
  logic [31:0] f2482_wdata;
  logic [0:0] f2482_clk;
  logic [0:0] f2482_rst;
  logic [31:0] f2482_rdata;
  sr_buffer_32_1 f2482(.wen(f2482_wen), .wdata(f2482_wdata), .clk(f2482_clk), .rst(f2482_rst), .rdata(f2482_rdata));
  assign f2482_clk = clk;
  assign f2482_rst = rst;
  // Bindings to f2482

  // f2484
  logic [0:0] f2484_wen;
  logic [31:0] f2484_wdata;
  logic [0:0] f2484_clk;
  logic [0:0] f2484_rst;
  logic [31:0] f2484_rdata;
  sr_buffer_32_1 f2484(.wen(f2484_wen), .wdata(f2484_wdata), .clk(f2484_clk), .rst(f2484_rst), .rdata(f2484_rdata));
  assign f2484_clk = clk;
  assign f2484_rst = rst;
  // Bindings to f2484

  // f2486
  logic [0:0] f2486_wen;
  logic [31:0] f2486_wdata;
  logic [0:0] f2486_clk;
  logic [0:0] f2486_rst;
  logic [31:0] f2486_rdata;
  sr_buffer_32_1 f2486(.wen(f2486_wen), .wdata(f2486_wdata), .clk(f2486_clk), .rst(f2486_rst), .rdata(f2486_rdata));
  assign f2486_clk = clk;
  assign f2486_rst = rst;
  // Bindings to f2486

  // f2488
  logic [0:0] f2488_wen;
  logic [31:0] f2488_wdata;
  logic [0:0] f2488_clk;
  logic [0:0] f2488_rst;
  logic [31:0] f2488_rdata;
  sr_buffer_32_1 f2488(.wen(f2488_wen), .wdata(f2488_wdata), .clk(f2488_clk), .rst(f2488_rst), .rdata(f2488_rdata));
  assign f2488_clk = clk;
  assign f2488_rst = rst;
  // Bindings to f2488

  // f2490
  logic [0:0] f2490_wen;
  logic [31:0] f2490_wdata;
  logic [0:0] f2490_clk;
  logic [0:0] f2490_rst;
  logic [31:0] f2490_rdata;
  sr_buffer_32_1 f2490(.wen(f2490_wen), .wdata(f2490_wdata), .clk(f2490_clk), .rst(f2490_rst), .rdata(f2490_rdata));
  assign f2490_clk = clk;
  assign f2490_rst = rst;
  // Bindings to f2490

  // f2492
  logic [0:0] f2492_wen;
  logic [31:0] f2492_wdata;
  logic [0:0] f2492_clk;
  logic [0:0] f2492_rst;
  logic [31:0] f2492_rdata;
  sr_buffer_32_1 f2492(.wen(f2492_wen), .wdata(f2492_wdata), .clk(f2492_clk), .rst(f2492_rst), .rdata(f2492_rdata));
  assign f2492_clk = clk;
  assign f2492_rst = rst;
  // Bindings to f2492

  // f2494
  logic [0:0] f2494_wen;
  logic [31:0] f2494_wdata;
  logic [0:0] f2494_clk;
  logic [0:0] f2494_rst;
  logic [31:0] f2494_rdata;
  sr_buffer_32_1 f2494(.wen(f2494_wen), .wdata(f2494_wdata), .clk(f2494_clk), .rst(f2494_rst), .rdata(f2494_rdata));
  assign f2494_clk = clk;
  assign f2494_rst = rst;
  // Bindings to f2494

  // f2496
  logic [0:0] f2496_wen;
  logic [31:0] f2496_wdata;
  logic [0:0] f2496_clk;
  logic [0:0] f2496_rst;
  logic [31:0] f2496_rdata;
  sr_buffer_32_1 f2496(.wen(f2496_wen), .wdata(f2496_wdata), .clk(f2496_clk), .rst(f2496_rst), .rdata(f2496_rdata));
  assign f2496_clk = clk;
  assign f2496_rst = rst;
  // Bindings to f2496

  // f2498
  logic [0:0] f2498_wen;
  logic [31:0] f2498_wdata;
  logic [0:0] f2498_clk;
  logic [0:0] f2498_rst;
  logic [31:0] f2498_rdata;
  sr_buffer_32_1 f2498(.wen(f2498_wen), .wdata(f2498_wdata), .clk(f2498_clk), .rst(f2498_rst), .rdata(f2498_rdata));
  assign f2498_clk = clk;
  assign f2498_rst = rst;
  // Bindings to f2498

  // f2500
  logic [0:0] f2500_wen;
  logic [31:0] f2500_wdata;
  logic [0:0] f2500_clk;
  logic [0:0] f2500_rst;
  logic [31:0] f2500_rdata;
  sr_buffer_32_1 f2500(.wen(f2500_wen), .wdata(f2500_wdata), .clk(f2500_clk), .rst(f2500_rst), .rdata(f2500_rdata));
  assign f2500_clk = clk;
  assign f2500_rst = rst;
  // Bindings to f2500

  // f2502
  logic [0:0] f2502_wen;
  logic [31:0] f2502_wdata;
  logic [0:0] f2502_clk;
  logic [0:0] f2502_rst;
  logic [31:0] f2502_rdata;
  sr_buffer_32_1 f2502(.wen(f2502_wen), .wdata(f2502_wdata), .clk(f2502_clk), .rst(f2502_rst), .rdata(f2502_rdata));
  assign f2502_clk = clk;
  assign f2502_rst = rst;
  // Bindings to f2502

  // f2504
  logic [0:0] f2504_wen;
  logic [31:0] f2504_wdata;
  logic [0:0] f2504_clk;
  logic [0:0] f2504_rst;
  logic [31:0] f2504_rdata;
  sr_buffer_32_1 f2504(.wen(f2504_wen), .wdata(f2504_wdata), .clk(f2504_clk), .rst(f2504_rst), .rdata(f2504_rdata));
  assign f2504_clk = clk;
  assign f2504_rst = rst;
  // Bindings to f2504

  // f2506
  logic [0:0] f2506_wen;
  logic [31:0] f2506_wdata;
  logic [0:0] f2506_clk;
  logic [0:0] f2506_rst;
  logic [31:0] f2506_rdata;
  sr_buffer_32_1 f2506(.wen(f2506_wen), .wdata(f2506_wdata), .clk(f2506_clk), .rst(f2506_rst), .rdata(f2506_rdata));
  assign f2506_clk = clk;
  assign f2506_rst = rst;
  // Bindings to f2506

  // f2508
  logic [0:0] f2508_wen;
  logic [31:0] f2508_wdata;
  logic [0:0] f2508_clk;
  logic [0:0] f2508_rst;
  logic [31:0] f2508_rdata;
  sr_buffer_32_1 f2508(.wen(f2508_wen), .wdata(f2508_wdata), .clk(f2508_clk), .rst(f2508_rst), .rdata(f2508_rdata));
  assign f2508_clk = clk;
  assign f2508_rst = rst;
  // Bindings to f2508

  // f2510
  logic [0:0] f2510_wen;
  logic [31:0] f2510_wdata;
  logic [0:0] f2510_clk;
  logic [0:0] f2510_rst;
  logic [31:0] f2510_rdata;
  sr_buffer_32_1 f2510(.wen(f2510_wen), .wdata(f2510_wdata), .clk(f2510_clk), .rst(f2510_rst), .rdata(f2510_rdata));
  assign f2510_clk = clk;
  assign f2510_rst = rst;
  // Bindings to f2510

  // f2512
  logic [0:0] f2512_wen;
  logic [31:0] f2512_wdata;
  logic [0:0] f2512_clk;
  logic [0:0] f2512_rst;
  logic [31:0] f2512_rdata;
  sr_buffer_32_1 f2512(.wen(f2512_wen), .wdata(f2512_wdata), .clk(f2512_clk), .rst(f2512_rst), .rdata(f2512_rdata));
  assign f2512_clk = clk;
  assign f2512_rst = rst;
  // Bindings to f2512

  // f2514
  logic [0:0] f2514_wen;
  logic [31:0] f2514_wdata;
  logic [0:0] f2514_clk;
  logic [0:0] f2514_rst;
  logic [31:0] f2514_rdata;
  sr_buffer_32_1 f2514(.wen(f2514_wen), .wdata(f2514_wdata), .clk(f2514_clk), .rst(f2514_rst), .rdata(f2514_rdata));
  assign f2514_clk = clk;
  assign f2514_rst = rst;
  // Bindings to f2514

  // f2516
  logic [0:0] f2516_wen;
  logic [31:0] f2516_wdata;
  logic [0:0] f2516_clk;
  logic [0:0] f2516_rst;
  logic [31:0] f2516_rdata;
  sr_buffer_32_1 f2516(.wen(f2516_wen), .wdata(f2516_wdata), .clk(f2516_clk), .rst(f2516_rst), .rdata(f2516_rdata));
  assign f2516_clk = clk;
  assign f2516_rst = rst;
  // Bindings to f2516

  // f2518
  logic [0:0] f2518_wen;
  logic [31:0] f2518_wdata;
  logic [0:0] f2518_clk;
  logic [0:0] f2518_rst;
  logic [31:0] f2518_rdata;
  sr_buffer_32_1 f2518(.wen(f2518_wen), .wdata(f2518_wdata), .clk(f2518_clk), .rst(f2518_rst), .rdata(f2518_rdata));
  assign f2518_clk = clk;
  assign f2518_rst = rst;
  // Bindings to f2518

  // f2520
  logic [0:0] f2520_wen;
  logic [31:0] f2520_wdata;
  logic [0:0] f2520_clk;
  logic [0:0] f2520_rst;
  logic [31:0] f2520_rdata;
  sr_buffer_32_1 f2520(.wen(f2520_wen), .wdata(f2520_wdata), .clk(f2520_clk), .rst(f2520_rst), .rdata(f2520_rdata));
  assign f2520_clk = clk;
  assign f2520_rst = rst;
  // Bindings to f2520

  // f2522
  logic [0:0] f2522_wen;
  logic [31:0] f2522_wdata;
  logic [0:0] f2522_clk;
  logic [0:0] f2522_rst;
  logic [31:0] f2522_rdata;
  sr_buffer_32_1 f2522(.wen(f2522_wen), .wdata(f2522_wdata), .clk(f2522_clk), .rst(f2522_rst), .rdata(f2522_rdata));
  assign f2522_clk = clk;
  assign f2522_rst = rst;
  // Bindings to f2522

  // f2524
  logic [0:0] f2524_wen;
  logic [31:0] f2524_wdata;
  logic [0:0] f2524_clk;
  logic [0:0] f2524_rst;
  logic [31:0] f2524_rdata;
  sr_buffer_32_1 f2524(.wen(f2524_wen), .wdata(f2524_wdata), .clk(f2524_clk), .rst(f2524_rst), .rdata(f2524_rdata));
  assign f2524_clk = clk;
  assign f2524_rst = rst;
  // Bindings to f2524

  // f2526
  logic [0:0] f2526_wen;
  logic [31:0] f2526_wdata;
  logic [0:0] f2526_clk;
  logic [0:0] f2526_rst;
  logic [31:0] f2526_rdata;
  sr_buffer_32_1 f2526(.wen(f2526_wen), .wdata(f2526_wdata), .clk(f2526_clk), .rst(f2526_rst), .rdata(f2526_rdata));
  assign f2526_clk = clk;
  assign f2526_rst = rst;
  // Bindings to f2526

  // f2528
  logic [0:0] f2528_wen;
  logic [31:0] f2528_wdata;
  logic [0:0] f2528_clk;
  logic [0:0] f2528_rst;
  logic [31:0] f2528_rdata;
  sr_buffer_32_1 f2528(.wen(f2528_wen), .wdata(f2528_wdata), .clk(f2528_clk), .rst(f2528_rst), .rdata(f2528_rdata));
  assign f2528_clk = clk;
  assign f2528_rst = rst;
  // Bindings to f2528

  // f2530
  logic [0:0] f2530_wen;
  logic [31:0] f2530_wdata;
  logic [0:0] f2530_clk;
  logic [0:0] f2530_rst;
  logic [31:0] f2530_rdata;
  sr_buffer_32_1 f2530(.wen(f2530_wen), .wdata(f2530_wdata), .clk(f2530_clk), .rst(f2530_rst), .rdata(f2530_rdata));
  assign f2530_clk = clk;
  assign f2530_rst = rst;
  // Bindings to f2530

  // f722
  logic [0:0] f722_wen;
  logic [31:0] f722_wdata;
  logic [0:0] f722_clk;
  logic [0:0] f722_rst;
  logic [31:0] f722_rdata;
  sr_buffer_32_1 f722(.wen(f722_wen), .wdata(f722_wdata), .clk(f722_clk), .rst(f722_rst), .rdata(f722_rdata));
  assign f722_clk = clk;
  assign f722_rst = rst;
  // Bindings to f722

  // f728
  logic [0:0] f728_wen;
  logic [31:0] f728_wdata;
  logic [0:0] f728_clk;
  logic [0:0] f728_rst;
  logic [31:0] f728_rdata;
  sr_buffer_32_1 f728(.wen(f728_wen), .wdata(f728_wdata), .clk(f728_clk), .rst(f728_rst), .rdata(f728_rdata));
  assign f728_clk = clk;
  assign f728_rst = rst;
  // Bindings to f728

  // f730
  logic [0:0] f730_wen;
  logic [31:0] f730_wdata;
  logic [0:0] f730_clk;
  logic [0:0] f730_rst;
  logic [31:0] f730_rdata;
  sr_buffer_32_1 f730(.wen(f730_wen), .wdata(f730_wdata), .clk(f730_clk), .rst(f730_rst), .rdata(f730_rdata));
  assign f730_clk = clk;
  assign f730_rst = rst;
  // Bindings to f730

  // f732
  logic [0:0] f732_wen;
  logic [31:0] f732_wdata;
  logic [0:0] f732_clk;
  logic [0:0] f732_rst;
  logic [31:0] f732_rdata;
  sr_buffer_32_1 f732(.wen(f732_wen), .wdata(f732_wdata), .clk(f732_clk), .rst(f732_rst), .rdata(f732_rdata));
  assign f732_clk = clk;
  assign f732_rst = rst;
  // Bindings to f732

  // f734
  logic [0:0] f734_wen;
  logic [31:0] f734_wdata;
  logic [0:0] f734_clk;
  logic [0:0] f734_rst;
  logic [31:0] f734_rdata;
  sr_buffer_32_1 f734(.wen(f734_wen), .wdata(f734_wdata), .clk(f734_clk), .rst(f734_rst), .rdata(f734_rdata));
  assign f734_clk = clk;
  assign f734_rst = rst;
  // Bindings to f734

  // f736
  logic [0:0] f736_wen;
  logic [31:0] f736_wdata;
  logic [0:0] f736_clk;
  logic [0:0] f736_rst;
  logic [31:0] f736_rdata;
  sr_buffer_32_1 f736(.wen(f736_wen), .wdata(f736_wdata), .clk(f736_clk), .rst(f736_rst), .rdata(f736_rdata));
  assign f736_clk = clk;
  assign f736_rst = rst;
  // Bindings to f736

  // f724
  logic [0:0] f724_wen;
  logic [31:0] f724_wdata;
  logic [0:0] f724_clk;
  logic [0:0] f724_rst;
  logic [31:0] f724_rdata;
  sr_buffer_32_1 f724(.wen(f724_wen), .wdata(f724_wdata), .clk(f724_clk), .rst(f724_rst), .rdata(f724_rdata));
  assign f724_clk = clk;
  assign f724_rst = rst;
  // Bindings to f724

  // f726
  logic [0:0] f726_wen;
  logic [31:0] f726_wdata;
  logic [0:0] f726_clk;
  logic [0:0] f726_rst;
  logic [31:0] f726_rdata;
  sr_buffer_32_1 f726(.wen(f726_wen), .wdata(f726_wdata), .clk(f726_clk), .rst(f726_rst), .rdata(f726_rdata));
  assign f726_clk = clk;
  assign f726_rst = rst;
  // Bindings to f726

  // f738
  logic [0:0] f738_wen;
  logic [31:0] f738_wdata;
  logic [0:0] f738_clk;
  logic [0:0] f738_rst;
  logic [31:0] f738_rdata;
  sr_buffer_32_1 f738(.wen(f738_wen), .wdata(f738_wdata), .clk(f738_clk), .rst(f738_rst), .rdata(f738_rdata));
  assign f738_clk = clk;
  assign f738_rst = rst;
  // Bindings to f738

  // f740
  logic [0:0] f740_wen;
  logic [31:0] f740_wdata;
  logic [0:0] f740_clk;
  logic [0:0] f740_rst;
  logic [31:0] f740_rdata;
  sr_buffer_32_1 f740(.wen(f740_wen), .wdata(f740_wdata), .clk(f740_clk), .rst(f740_rst), .rdata(f740_rdata));
  assign f740_clk = clk;
  assign f740_rst = rst;
  // Bindings to f740

  // f742
  logic [0:0] f742_wen;
  logic [31:0] f742_wdata;
  logic [0:0] f742_clk;
  logic [0:0] f742_rst;
  logic [31:0] f742_rdata;
  sr_buffer_32_1 f742(.wen(f742_wen), .wdata(f742_wdata), .clk(f742_clk), .rst(f742_rst), .rdata(f742_rdata));
  assign f742_clk = clk;
  assign f742_rst = rst;
  // Bindings to f742

  // f744
  logic [0:0] f744_wen;
  logic [31:0] f744_wdata;
  logic [0:0] f744_clk;
  logic [0:0] f744_rst;
  logic [31:0] f744_rdata;
  sr_buffer_32_1 f744(.wen(f744_wen), .wdata(f744_wdata), .clk(f744_clk), .rst(f744_rst), .rdata(f744_rdata));
  assign f744_clk = clk;
  assign f744_rst = rst;
  // Bindings to f744

  // f746
  logic [0:0] f746_wen;
  logic [31:0] f746_wdata;
  logic [0:0] f746_clk;
  logic [0:0] f746_rst;
  logic [31:0] f746_rdata;
  sr_buffer_32_1 f746(.wen(f746_wen), .wdata(f746_wdata), .clk(f746_clk), .rst(f746_rst), .rdata(f746_rdata));
  assign f746_clk = clk;
  assign f746_rst = rst;
  // Bindings to f746

  // f748
  logic [0:0] f748_wen;
  logic [31:0] f748_wdata;
  logic [0:0] f748_clk;
  logic [0:0] f748_rst;
  logic [31:0] f748_rdata;
  sr_buffer_32_1 f748(.wen(f748_wen), .wdata(f748_wdata), .clk(f748_clk), .rst(f748_rst), .rdata(f748_rdata));
  assign f748_clk = clk;
  assign f748_rst = rst;
  // Bindings to f748

  // f750
  logic [0:0] f750_wen;
  logic [31:0] f750_wdata;
  logic [0:0] f750_clk;
  logic [0:0] f750_rst;
  logic [31:0] f750_rdata;
  sr_buffer_32_1 f750(.wen(f750_wen), .wdata(f750_wdata), .clk(f750_clk), .rst(f750_rst), .rdata(f750_rdata));
  assign f750_clk = clk;
  assign f750_rst = rst;
  // Bindings to f750

  // f752
  logic [0:0] f752_wen;
  logic [31:0] f752_wdata;
  logic [0:0] f752_clk;
  logic [0:0] f752_rst;
  logic [31:0] f752_rdata;
  sr_buffer_32_1 f752(.wen(f752_wen), .wdata(f752_wdata), .clk(f752_clk), .rst(f752_rst), .rdata(f752_rdata));
  assign f752_clk = clk;
  assign f752_rst = rst;
  // Bindings to f752

  // f754
  logic [0:0] f754_wen;
  logic [31:0] f754_wdata;
  logic [0:0] f754_clk;
  logic [0:0] f754_rst;
  logic [31:0] f754_rdata;
  sr_buffer_32_1 f754(.wen(f754_wen), .wdata(f754_wdata), .clk(f754_clk), .rst(f754_rst), .rdata(f754_rdata));
  assign f754_clk = clk;
  assign f754_rst = rst;
  // Bindings to f754

  // f756
  logic [0:0] f756_wen;
  logic [31:0] f756_wdata;
  logic [0:0] f756_clk;
  logic [0:0] f756_rst;
  logic [31:0] f756_rdata;
  sr_buffer_32_1 f756(.wen(f756_wen), .wdata(f756_wdata), .clk(f756_clk), .rst(f756_rst), .rdata(f756_rdata));
  assign f756_clk = clk;
  assign f756_rst = rst;
  // Bindings to f756

  // f758
  logic [0:0] f758_wen;
  logic [31:0] f758_wdata;
  logic [0:0] f758_clk;
  logic [0:0] f758_rst;
  logic [31:0] f758_rdata;
  sr_buffer_32_1 f758(.wen(f758_wen), .wdata(f758_wdata), .clk(f758_clk), .rst(f758_rst), .rdata(f758_rdata));
  assign f758_clk = clk;
  assign f758_rst = rst;
  // Bindings to f758

  // f760
  logic [0:0] f760_wen;
  logic [31:0] f760_wdata;
  logic [0:0] f760_clk;
  logic [0:0] f760_rst;
  logic [31:0] f760_rdata;
  sr_buffer_32_1 f760(.wen(f760_wen), .wdata(f760_wdata), .clk(f760_clk), .rst(f760_rst), .rdata(f760_rdata));
  assign f760_clk = clk;
  assign f760_rst = rst;
  // Bindings to f760

  // f762
  logic [0:0] f762_wen;
  logic [31:0] f762_wdata;
  logic [0:0] f762_clk;
  logic [0:0] f762_rst;
  logic [31:0] f762_rdata;
  sr_buffer_32_1 f762(.wen(f762_wen), .wdata(f762_wdata), .clk(f762_clk), .rst(f762_rst), .rdata(f762_rdata));
  assign f762_clk = clk;
  assign f762_rst = rst;
  // Bindings to f762

  // f764
  logic [0:0] f764_wen;
  logic [31:0] f764_wdata;
  logic [0:0] f764_clk;
  logic [0:0] f764_rst;
  logic [31:0] f764_rdata;
  sr_buffer_32_1 f764(.wen(f764_wen), .wdata(f764_wdata), .clk(f764_clk), .rst(f764_rst), .rdata(f764_rdata));
  assign f764_clk = clk;
  assign f764_rst = rst;
  // Bindings to f764

  // f766
  logic [0:0] f766_wen;
  logic [31:0] f766_wdata;
  logic [0:0] f766_clk;
  logic [0:0] f766_rst;
  logic [31:0] f766_rdata;
  sr_buffer_32_1 f766(.wen(f766_wen), .wdata(f766_wdata), .clk(f766_clk), .rst(f766_rst), .rdata(f766_rdata));
  assign f766_clk = clk;
  assign f766_rst = rst;
  // Bindings to f766

  // f768
  logic [0:0] f768_wen;
  logic [31:0] f768_wdata;
  logic [0:0] f768_clk;
  logic [0:0] f768_rst;
  logic [31:0] f768_rdata;
  sr_buffer_32_1 f768(.wen(f768_wen), .wdata(f768_wdata), .clk(f768_clk), .rst(f768_rst), .rdata(f768_rdata));
  assign f768_clk = clk;
  assign f768_rst = rst;
  // Bindings to f768

  // f770
  logic [0:0] f770_wen;
  logic [31:0] f770_wdata;
  logic [0:0] f770_clk;
  logic [0:0] f770_rst;
  logic [31:0] f770_rdata;
  sr_buffer_32_1 f770(.wen(f770_wen), .wdata(f770_wdata), .clk(f770_clk), .rst(f770_rst), .rdata(f770_rdata));
  assign f770_clk = clk;
  assign f770_rst = rst;
  // Bindings to f770

  // f772
  logic [0:0] f772_wen;
  logic [31:0] f772_wdata;
  logic [0:0] f772_clk;
  logic [0:0] f772_rst;
  logic [31:0] f772_rdata;
  sr_buffer_32_1 f772(.wen(f772_wen), .wdata(f772_wdata), .clk(f772_clk), .rst(f772_rst), .rdata(f772_rdata));
  assign f772_clk = clk;
  assign f772_rst = rst;
  // Bindings to f772

  // f774
  logic [0:0] f774_wen;
  logic [31:0] f774_wdata;
  logic [0:0] f774_clk;
  logic [0:0] f774_rst;
  logic [31:0] f774_rdata;
  sr_buffer_32_1 f774(.wen(f774_wen), .wdata(f774_wdata), .clk(f774_clk), .rst(f774_rst), .rdata(f774_rdata));
  assign f774_clk = clk;
  assign f774_rst = rst;
  // Bindings to f774

  // f776
  logic [0:0] f776_wen;
  logic [31:0] f776_wdata;
  logic [0:0] f776_clk;
  logic [0:0] f776_rst;
  logic [31:0] f776_rdata;
  sr_buffer_32_1 f776(.wen(f776_wen), .wdata(f776_wdata), .clk(f776_clk), .rst(f776_rst), .rdata(f776_rdata));
  assign f776_clk = clk;
  assign f776_rst = rst;
  // Bindings to f776

  // f778
  logic [0:0] f778_wen;
  logic [31:0] f778_wdata;
  logic [0:0] f778_clk;
  logic [0:0] f778_rst;
  logic [31:0] f778_rdata;
  sr_buffer_32_1 f778(.wen(f778_wen), .wdata(f778_wdata), .clk(f778_clk), .rst(f778_rst), .rdata(f778_rdata));
  assign f778_clk = clk;
  assign f778_rst = rst;
  // Bindings to f778

  // f780
  logic [0:0] f780_wen;
  logic [31:0] f780_wdata;
  logic [0:0] f780_clk;
  logic [0:0] f780_rst;
  logic [31:0] f780_rdata;
  sr_buffer_32_1 f780(.wen(f780_wen), .wdata(f780_wdata), .clk(f780_clk), .rst(f780_rst), .rdata(f780_rdata));
  assign f780_clk = clk;
  assign f780_rst = rst;
  // Bindings to f780

  // f782
  logic [0:0] f782_wen;
  logic [31:0] f782_wdata;
  logic [0:0] f782_clk;
  logic [0:0] f782_rst;
  logic [31:0] f782_rdata;
  sr_buffer_32_1 f782(.wen(f782_wen), .wdata(f782_wdata), .clk(f782_clk), .rst(f782_rst), .rdata(f782_rdata));
  assign f782_clk = clk;
  assign f782_rst = rst;
  // Bindings to f782

  // f784
  logic [0:0] f784_wen;
  logic [31:0] f784_wdata;
  logic [0:0] f784_clk;
  logic [0:0] f784_rst;
  logic [31:0] f784_rdata;
  sr_buffer_32_1 f784(.wen(f784_wen), .wdata(f784_wdata), .clk(f784_clk), .rst(f784_rst), .rdata(f784_rdata));
  assign f784_clk = clk;
  assign f784_rst = rst;
  // Bindings to f784

  // f786
  logic [0:0] f786_wen;
  logic [31:0] f786_wdata;
  logic [0:0] f786_clk;
  logic [0:0] f786_rst;
  logic [31:0] f786_rdata;
  sr_buffer_32_1 f786(.wen(f786_wen), .wdata(f786_wdata), .clk(f786_clk), .rst(f786_rst), .rdata(f786_rdata));
  assign f786_clk = clk;
  assign f786_rst = rst;
  // Bindings to f786

  // f788
  logic [0:0] f788_wen;
  logic [31:0] f788_wdata;
  logic [0:0] f788_clk;
  logic [0:0] f788_rst;
  logic [31:0] f788_rdata;
  sr_buffer_32_1 f788(.wen(f788_wen), .wdata(f788_wdata), .clk(f788_clk), .rst(f788_rst), .rdata(f788_rdata));
  assign f788_clk = clk;
  assign f788_rst = rst;
  // Bindings to f788

  // f790
  logic [0:0] f790_wen;
  logic [31:0] f790_wdata;
  logic [0:0] f790_clk;
  logic [0:0] f790_rst;
  logic [31:0] f790_rdata;
  sr_buffer_32_1 f790(.wen(f790_wen), .wdata(f790_wdata), .clk(f790_clk), .rst(f790_rst), .rdata(f790_rdata));
  assign f790_clk = clk;
  assign f790_rst = rst;
  // Bindings to f790

  // f792
  logic [0:0] f792_wen;
  logic [31:0] f792_wdata;
  logic [0:0] f792_clk;
  logic [0:0] f792_rst;
  logic [31:0] f792_rdata;
  sr_buffer_32_1 f792(.wen(f792_wen), .wdata(f792_wdata), .clk(f792_clk), .rst(f792_rst), .rdata(f792_rdata));
  assign f792_clk = clk;
  assign f792_rst = rst;
  // Bindings to f792

  // f794
  logic [0:0] f794_wen;
  logic [31:0] f794_wdata;
  logic [0:0] f794_clk;
  logic [0:0] f794_rst;
  logic [31:0] f794_rdata;
  sr_buffer_32_1 f794(.wen(f794_wen), .wdata(f794_wdata), .clk(f794_clk), .rst(f794_rst), .rdata(f794_rdata));
  assign f794_clk = clk;
  assign f794_rst = rst;
  // Bindings to f794

  // f796
  logic [0:0] f796_wen;
  logic [31:0] f796_wdata;
  logic [0:0] f796_clk;
  logic [0:0] f796_rst;
  logic [31:0] f796_rdata;
  sr_buffer_32_1 f796(.wen(f796_wen), .wdata(f796_wdata), .clk(f796_clk), .rst(f796_rst), .rdata(f796_rdata));
  assign f796_clk = clk;
  assign f796_rst = rst;
  // Bindings to f796

  // f798
  logic [0:0] f798_wen;
  logic [31:0] f798_wdata;
  logic [0:0] f798_clk;
  logic [0:0] f798_rst;
  logic [31:0] f798_rdata;
  sr_buffer_32_1 f798(.wen(f798_wen), .wdata(f798_wdata), .clk(f798_clk), .rst(f798_rst), .rdata(f798_rdata));
  assign f798_clk = clk;
  assign f798_rst = rst;
  // Bindings to f798

  // f800
  logic [0:0] f800_wen;
  logic [31:0] f800_wdata;
  logic [0:0] f800_clk;
  logic [0:0] f800_rst;
  logic [31:0] f800_rdata;
  sr_buffer_32_1 f800(.wen(f800_wen), .wdata(f800_wdata), .clk(f800_clk), .rst(f800_rst), .rdata(f800_rdata));
  assign f800_clk = clk;
  assign f800_rst = rst;
  // Bindings to f800

  // f802
  logic [0:0] f802_wen;
  logic [31:0] f802_wdata;
  logic [0:0] f802_clk;
  logic [0:0] f802_rst;
  logic [31:0] f802_rdata;
  sr_buffer_32_1 f802(.wen(f802_wen), .wdata(f802_wdata), .clk(f802_clk), .rst(f802_rst), .rdata(f802_rdata));
  assign f802_clk = clk;
  assign f802_rst = rst;
  // Bindings to f802

  // f806
  logic [0:0] f806_wen;
  logic [31:0] f806_wdata;
  logic [0:0] f806_clk;
  logic [0:0] f806_rst;
  logic [31:0] f806_rdata;
  sr_buffer_32_1 f806(.wen(f806_wen), .wdata(f806_wdata), .clk(f806_clk), .rst(f806_rst), .rdata(f806_rdata));
  assign f806_clk = clk;
  assign f806_rst = rst;
  // Bindings to f806

  // f808
  logic [0:0] f808_wen;
  logic [31:0] f808_wdata;
  logic [0:0] f808_clk;
  logic [0:0] f808_rst;
  logic [31:0] f808_rdata;
  sr_buffer_32_1 f808(.wen(f808_wen), .wdata(f808_wdata), .clk(f808_clk), .rst(f808_rst), .rdata(f808_rdata));
  assign f808_clk = clk;
  assign f808_rst = rst;
  // Bindings to f808

  // f810
  logic [0:0] f810_wen;
  logic [31:0] f810_wdata;
  logic [0:0] f810_clk;
  logic [0:0] f810_rst;
  logic [31:0] f810_rdata;
  sr_buffer_32_1 f810(.wen(f810_wen), .wdata(f810_wdata), .clk(f810_clk), .rst(f810_rst), .rdata(f810_rdata));
  assign f810_clk = clk;
  assign f810_rst = rst;
  // Bindings to f810

  // f812
  logic [0:0] f812_wen;
  logic [31:0] f812_wdata;
  logic [0:0] f812_clk;
  logic [0:0] f812_rst;
  logic [31:0] f812_rdata;
  sr_buffer_32_1 f812(.wen(f812_wen), .wdata(f812_wdata), .clk(f812_clk), .rst(f812_rst), .rdata(f812_rdata));
  assign f812_clk = clk;
  assign f812_rst = rst;
  // Bindings to f812

  // f814
  logic [0:0] f814_wen;
  logic [31:0] f814_wdata;
  logic [0:0] f814_clk;
  logic [0:0] f814_rst;
  logic [31:0] f814_rdata;
  sr_buffer_32_1 f814(.wen(f814_wen), .wdata(f814_wdata), .clk(f814_clk), .rst(f814_rst), .rdata(f814_rdata));
  assign f814_clk = clk;
  assign f814_rst = rst;
  // Bindings to f814

  // f816
  logic [0:0] f816_wen;
  logic [31:0] f816_wdata;
  logic [0:0] f816_clk;
  logic [0:0] f816_rst;
  logic [31:0] f816_rdata;
  sr_buffer_32_1 f816(.wen(f816_wen), .wdata(f816_wdata), .clk(f816_clk), .rst(f816_rst), .rdata(f816_rdata));
  assign f816_clk = clk;
  assign f816_rst = rst;
  // Bindings to f816

  // f818
  logic [0:0] f818_wen;
  logic [31:0] f818_wdata;
  logic [0:0] f818_clk;
  logic [0:0] f818_rst;
  logic [31:0] f818_rdata;
  sr_buffer_32_1 f818(.wen(f818_wen), .wdata(f818_wdata), .clk(f818_clk), .rst(f818_rst), .rdata(f818_rdata));
  assign f818_clk = clk;
  assign f818_rst = rst;
  // Bindings to f818

  // f820
  logic [0:0] f820_wen;
  logic [31:0] f820_wdata;
  logic [0:0] f820_clk;
  logic [0:0] f820_rst;
  logic [31:0] f820_rdata;
  sr_buffer_32_1 f820(.wen(f820_wen), .wdata(f820_wdata), .clk(f820_clk), .rst(f820_rst), .rdata(f820_rdata));
  assign f820_clk = clk;
  assign f820_rst = rst;
  // Bindings to f820

  // f822
  logic [0:0] f822_wen;
  logic [31:0] f822_wdata;
  logic [0:0] f822_clk;
  logic [0:0] f822_rst;
  logic [31:0] f822_rdata;
  sr_buffer_32_1 f822(.wen(f822_wen), .wdata(f822_wdata), .clk(f822_clk), .rst(f822_rst), .rdata(f822_rdata));
  assign f822_clk = clk;
  assign f822_rst = rst;
  // Bindings to f822

  // f824
  logic [0:0] f824_wen;
  logic [31:0] f824_wdata;
  logic [0:0] f824_clk;
  logic [0:0] f824_rst;
  logic [31:0] f824_rdata;
  sr_buffer_32_1 f824(.wen(f824_wen), .wdata(f824_wdata), .clk(f824_clk), .rst(f824_rst), .rdata(f824_rdata));
  assign f824_clk = clk;
  assign f824_rst = rst;
  // Bindings to f824

  // f826
  logic [0:0] f826_wen;
  logic [31:0] f826_wdata;
  logic [0:0] f826_clk;
  logic [0:0] f826_rst;
  logic [31:0] f826_rdata;
  sr_buffer_32_1 f826(.wen(f826_wen), .wdata(f826_wdata), .clk(f826_clk), .rst(f826_rst), .rdata(f826_rdata));
  assign f826_clk = clk;
  assign f826_rst = rst;
  // Bindings to f826

  // f828
  logic [0:0] f828_wen;
  logic [31:0] f828_wdata;
  logic [0:0] f828_clk;
  logic [0:0] f828_rst;
  logic [31:0] f828_rdata;
  sr_buffer_32_1 f828(.wen(f828_wen), .wdata(f828_wdata), .clk(f828_clk), .rst(f828_rst), .rdata(f828_rdata));
  assign f828_clk = clk;
  assign f828_rst = rst;
  // Bindings to f828

  // f830
  logic [0:0] f830_wen;
  logic [31:0] f830_wdata;
  logic [0:0] f830_clk;
  logic [0:0] f830_rst;
  logic [31:0] f830_rdata;
  sr_buffer_32_1 f830(.wen(f830_wen), .wdata(f830_wdata), .clk(f830_clk), .rst(f830_rst), .rdata(f830_rdata));
  assign f830_clk = clk;
  assign f830_rst = rst;
  // Bindings to f830

  // f832
  logic [0:0] f832_wen;
  logic [31:0] f832_wdata;
  logic [0:0] f832_clk;
  logic [0:0] f832_rst;
  logic [31:0] f832_rdata;
  sr_buffer_32_1 f832(.wen(f832_wen), .wdata(f832_wdata), .clk(f832_clk), .rst(f832_rst), .rdata(f832_rdata));
  assign f832_clk = clk;
  assign f832_rst = rst;
  // Bindings to f832

  // f834
  logic [0:0] f834_wen;
  logic [31:0] f834_wdata;
  logic [0:0] f834_clk;
  logic [0:0] f834_rst;
  logic [31:0] f834_rdata;
  sr_buffer_32_1 f834(.wen(f834_wen), .wdata(f834_wdata), .clk(f834_clk), .rst(f834_rst), .rdata(f834_rdata));
  assign f834_clk = clk;
  assign f834_rst = rst;
  // Bindings to f834

  // f836
  logic [0:0] f836_wen;
  logic [31:0] f836_wdata;
  logic [0:0] f836_clk;
  logic [0:0] f836_rst;
  logic [31:0] f836_rdata;
  sr_buffer_32_1 f836(.wen(f836_wen), .wdata(f836_wdata), .clk(f836_clk), .rst(f836_rst), .rdata(f836_rdata));
  assign f836_clk = clk;
  assign f836_rst = rst;
  // Bindings to f836

  // f840
  logic [0:0] f840_wen;
  logic [31:0] f840_wdata;
  logic [0:0] f840_clk;
  logic [0:0] f840_rst;
  logic [31:0] f840_rdata;
  sr_buffer_32_1 f840(.wen(f840_wen), .wdata(f840_wdata), .clk(f840_clk), .rst(f840_rst), .rdata(f840_rdata));
  assign f840_clk = clk;
  assign f840_rst = rst;
  // Bindings to f840

  // f846
  logic [0:0] f846_wen;
  logic [31:0] f846_wdata;
  logic [0:0] f846_clk;
  logic [0:0] f846_rst;
  logic [31:0] f846_rdata;
  sr_buffer_32_1 f846(.wen(f846_wen), .wdata(f846_wdata), .clk(f846_clk), .rst(f846_rst), .rdata(f846_rdata));
  assign f846_clk = clk;
  assign f846_rst = rst;
  // Bindings to f846

  // f848
  logic [0:0] f848_wen;
  logic [31:0] f848_wdata;
  logic [0:0] f848_clk;
  logic [0:0] f848_rst;
  logic [31:0] f848_rdata;
  sr_buffer_32_1 f848(.wen(f848_wen), .wdata(f848_wdata), .clk(f848_clk), .rst(f848_rst), .rdata(f848_rdata));
  assign f848_clk = clk;
  assign f848_rst = rst;
  // Bindings to f848

  // f852
  logic [0:0] f852_wen;
  logic [31:0] f852_wdata;
  logic [0:0] f852_clk;
  logic [0:0] f852_rst;
  logic [31:0] f852_rdata;
  sr_buffer_32_1 f852(.wen(f852_wen), .wdata(f852_wdata), .clk(f852_clk), .rst(f852_rst), .rdata(f852_rdata));
  assign f852_clk = clk;
  assign f852_rst = rst;
  // Bindings to f852

  // f854
  logic [0:0] f854_wen;
  logic [31:0] f854_wdata;
  logic [0:0] f854_clk;
  logic [0:0] f854_rst;
  logic [31:0] f854_rdata;
  sr_buffer_32_1 f854(.wen(f854_wen), .wdata(f854_wdata), .clk(f854_clk), .rst(f854_rst), .rdata(f854_rdata));
  assign f854_clk = clk;
  assign f854_rst = rst;
  // Bindings to f854

  // f856
  logic [0:0] f856_wen;
  logic [31:0] f856_wdata;
  logic [0:0] f856_clk;
  logic [0:0] f856_rst;
  logic [31:0] f856_rdata;
  sr_buffer_32_1 f856(.wen(f856_wen), .wdata(f856_wdata), .clk(f856_clk), .rst(f856_rst), .rdata(f856_rdata));
  assign f856_clk = clk;
  assign f856_rst = rst;
  // Bindings to f856

  // f858
  logic [0:0] f858_wen;
  logic [31:0] f858_wdata;
  logic [0:0] f858_clk;
  logic [0:0] f858_rst;
  logic [31:0] f858_rdata;
  sr_buffer_32_1 f858(.wen(f858_wen), .wdata(f858_wdata), .clk(f858_clk), .rst(f858_rst), .rdata(f858_rdata));
  assign f858_clk = clk;
  assign f858_rst = rst;
  // Bindings to f858

  // f860
  logic [0:0] f860_wen;
  logic [31:0] f860_wdata;
  logic [0:0] f860_clk;
  logic [0:0] f860_rst;
  logic [31:0] f860_rdata;
  sr_buffer_32_1 f860(.wen(f860_wen), .wdata(f860_wdata), .clk(f860_clk), .rst(f860_rst), .rdata(f860_rdata));
  assign f860_clk = clk;
  assign f860_rst = rst;
  // Bindings to f860

  // f862
  logic [0:0] f862_wen;
  logic [31:0] f862_wdata;
  logic [0:0] f862_clk;
  logic [0:0] f862_rst;
  logic [31:0] f862_rdata;
  sr_buffer_32_1 f862(.wen(f862_wen), .wdata(f862_wdata), .clk(f862_clk), .rst(f862_rst), .rdata(f862_rdata));
  assign f862_clk = clk;
  assign f862_rst = rst;
  // Bindings to f862

  // f864
  logic [0:0] f864_wen;
  logic [31:0] f864_wdata;
  logic [0:0] f864_clk;
  logic [0:0] f864_rst;
  logic [31:0] f864_rdata;
  sr_buffer_32_1 f864(.wen(f864_wen), .wdata(f864_wdata), .clk(f864_clk), .rst(f864_rst), .rdata(f864_rdata));
  assign f864_clk = clk;
  assign f864_rst = rst;
  // Bindings to f864

  // f866
  logic [0:0] f866_wen;
  logic [31:0] f866_wdata;
  logic [0:0] f866_clk;
  logic [0:0] f866_rst;
  logic [31:0] f866_rdata;
  sr_buffer_32_1 f866(.wen(f866_wen), .wdata(f866_wdata), .clk(f866_clk), .rst(f866_rst), .rdata(f866_rdata));
  assign f866_clk = clk;
  assign f866_rst = rst;
  // Bindings to f866

  // f868
  logic [0:0] f868_wen;
  logic [31:0] f868_wdata;
  logic [0:0] f868_clk;
  logic [0:0] f868_rst;
  logic [31:0] f868_rdata;
  sr_buffer_32_1 f868(.wen(f868_wen), .wdata(f868_wdata), .clk(f868_clk), .rst(f868_rst), .rdata(f868_rdata));
  assign f868_clk = clk;
  assign f868_rst = rst;
  // Bindings to f868

  // f870
  logic [0:0] f870_wen;
  logic [31:0] f870_wdata;
  logic [0:0] f870_clk;
  logic [0:0] f870_rst;
  logic [31:0] f870_rdata;
  sr_buffer_32_1 f870(.wen(f870_wen), .wdata(f870_wdata), .clk(f870_clk), .rst(f870_rst), .rdata(f870_rdata));
  assign f870_clk = clk;
  assign f870_rst = rst;
  // Bindings to f870

  // f872
  logic [0:0] f872_wen;
  logic [31:0] f872_wdata;
  logic [0:0] f872_clk;
  logic [0:0] f872_rst;
  logic [31:0] f872_rdata;
  sr_buffer_32_1 f872(.wen(f872_wen), .wdata(f872_wdata), .clk(f872_clk), .rst(f872_rst), .rdata(f872_rdata));
  assign f872_clk = clk;
  assign f872_rst = rst;
  // Bindings to f872

  // f874
  logic [0:0] f874_wen;
  logic [31:0] f874_wdata;
  logic [0:0] f874_clk;
  logic [0:0] f874_rst;
  logic [31:0] f874_rdata;
  sr_buffer_32_1 f874(.wen(f874_wen), .wdata(f874_wdata), .clk(f874_clk), .rst(f874_rst), .rdata(f874_rdata));
  assign f874_clk = clk;
  assign f874_rst = rst;
  // Bindings to f874

  // f876
  logic [0:0] f876_wen;
  logic [31:0] f876_wdata;
  logic [0:0] f876_clk;
  logic [0:0] f876_rst;
  logic [31:0] f876_rdata;
  sr_buffer_32_1 f876(.wen(f876_wen), .wdata(f876_wdata), .clk(f876_clk), .rst(f876_rst), .rdata(f876_rdata));
  assign f876_clk = clk;
  assign f876_rst = rst;
  // Bindings to f876

  // f878
  logic [0:0] f878_wen;
  logic [31:0] f878_wdata;
  logic [0:0] f878_clk;
  logic [0:0] f878_rst;
  logic [31:0] f878_rdata;
  sr_buffer_32_1 f878(.wen(f878_wen), .wdata(f878_wdata), .clk(f878_clk), .rst(f878_rst), .rdata(f878_rdata));
  assign f878_clk = clk;
  assign f878_rst = rst;
  // Bindings to f878

  // f880
  logic [0:0] f880_wen;
  logic [31:0] f880_wdata;
  logic [0:0] f880_clk;
  logic [0:0] f880_rst;
  logic [31:0] f880_rdata;
  sr_buffer_32_1 f880(.wen(f880_wen), .wdata(f880_wdata), .clk(f880_clk), .rst(f880_rst), .rdata(f880_rdata));
  assign f880_clk = clk;
  assign f880_rst = rst;
  // Bindings to f880

  // f882
  logic [0:0] f882_wen;
  logic [31:0] f882_wdata;
  logic [0:0] f882_clk;
  logic [0:0] f882_rst;
  logic [31:0] f882_rdata;
  sr_buffer_32_1 f882(.wen(f882_wen), .wdata(f882_wdata), .clk(f882_clk), .rst(f882_rst), .rdata(f882_rdata));
  assign f882_clk = clk;
  assign f882_rst = rst;
  // Bindings to f882

  // f884
  logic [0:0] f884_wen;
  logic [31:0] f884_wdata;
  logic [0:0] f884_clk;
  logic [0:0] f884_rst;
  logic [31:0] f884_rdata;
  sr_buffer_32_1 f884(.wen(f884_wen), .wdata(f884_wdata), .clk(f884_clk), .rst(f884_rst), .rdata(f884_rdata));
  assign f884_clk = clk;
  assign f884_rst = rst;
  // Bindings to f884

  // f886
  logic [0:0] f886_wen;
  logic [31:0] f886_wdata;
  logic [0:0] f886_clk;
  logic [0:0] f886_rst;
  logic [31:0] f886_rdata;
  sr_buffer_32_1 f886(.wen(f886_wen), .wdata(f886_wdata), .clk(f886_clk), .rst(f886_rst), .rdata(f886_rdata));
  assign f886_clk = clk;
  assign f886_rst = rst;
  // Bindings to f886

  // f888
  logic [0:0] f888_wen;
  logic [31:0] f888_wdata;
  logic [0:0] f888_clk;
  logic [0:0] f888_rst;
  logic [31:0] f888_rdata;
  sr_buffer_32_1 f888(.wen(f888_wen), .wdata(f888_wdata), .clk(f888_clk), .rst(f888_rst), .rdata(f888_rdata));
  assign f888_clk = clk;
  assign f888_rst = rst;
  // Bindings to f888

  // f890
  logic [0:0] f890_wen;
  logic [31:0] f890_wdata;
  logic [0:0] f890_clk;
  logic [0:0] f890_rst;
  logic [31:0] f890_rdata;
  sr_buffer_32_1 f890(.wen(f890_wen), .wdata(f890_wdata), .clk(f890_clk), .rst(f890_rst), .rdata(f890_rdata));
  assign f890_clk = clk;
  assign f890_rst = rst;
  // Bindings to f890

  // f892
  logic [0:0] f892_wen;
  logic [31:0] f892_wdata;
  logic [0:0] f892_clk;
  logic [0:0] f892_rst;
  logic [31:0] f892_rdata;
  sr_buffer_32_1 f892(.wen(f892_wen), .wdata(f892_wdata), .clk(f892_clk), .rst(f892_rst), .rdata(f892_rdata));
  assign f892_clk = clk;
  assign f892_rst = rst;
  // Bindings to f892

  // f894
  logic [0:0] f894_wen;
  logic [31:0] f894_wdata;
  logic [0:0] f894_clk;
  logic [0:0] f894_rst;
  logic [31:0] f894_rdata;
  sr_buffer_32_1 f894(.wen(f894_wen), .wdata(f894_wdata), .clk(f894_clk), .rst(f894_rst), .rdata(f894_rdata));
  assign f894_clk = clk;
  assign f894_rst = rst;
  // Bindings to f894

  // f896
  logic [0:0] f896_wen;
  logic [31:0] f896_wdata;
  logic [0:0] f896_clk;
  logic [0:0] f896_rst;
  logic [31:0] f896_rdata;
  sr_buffer_32_1 f896(.wen(f896_wen), .wdata(f896_wdata), .clk(f896_clk), .rst(f896_rst), .rdata(f896_rdata));
  assign f896_clk = clk;
  assign f896_rst = rst;
  // Bindings to f896

  // f898
  logic [0:0] f898_wen;
  logic [31:0] f898_wdata;
  logic [0:0] f898_clk;
  logic [0:0] f898_rst;
  logic [31:0] f898_rdata;
  sr_buffer_32_1 f898(.wen(f898_wen), .wdata(f898_wdata), .clk(f898_clk), .rst(f898_rst), .rdata(f898_rdata));
  assign f898_clk = clk;
  assign f898_rst = rst;
  // Bindings to f898

  // f900
  logic [0:0] f900_wen;
  logic [31:0] f900_wdata;
  logic [0:0] f900_clk;
  logic [0:0] f900_rst;
  logic [31:0] f900_rdata;
  sr_buffer_32_1 f900(.wen(f900_wen), .wdata(f900_wdata), .clk(f900_clk), .rst(f900_rst), .rdata(f900_rdata));
  assign f900_clk = clk;
  assign f900_rst = rst;
  // Bindings to f900

  // f902
  logic [0:0] f902_wen;
  logic [31:0] f902_wdata;
  logic [0:0] f902_clk;
  logic [0:0] f902_rst;
  logic [31:0] f902_rdata;
  sr_buffer_32_1 f902(.wen(f902_wen), .wdata(f902_wdata), .clk(f902_clk), .rst(f902_rst), .rdata(f902_rdata));
  assign f902_clk = clk;
  assign f902_rst = rst;
  // Bindings to f902

  // f904
  logic [0:0] f904_wen;
  logic [31:0] f904_wdata;
  logic [0:0] f904_clk;
  logic [0:0] f904_rst;
  logic [31:0] f904_rdata;
  sr_buffer_32_1 f904(.wen(f904_wen), .wdata(f904_wdata), .clk(f904_clk), .rst(f904_rst), .rdata(f904_rdata));
  assign f904_clk = clk;
  assign f904_rst = rst;
  // Bindings to f904

  // f906
  logic [0:0] f906_wen;
  logic [31:0] f906_wdata;
  logic [0:0] f906_clk;
  logic [0:0] f906_rst;
  logic [31:0] f906_rdata;
  sr_buffer_32_1 f906(.wen(f906_wen), .wdata(f906_wdata), .clk(f906_clk), .rst(f906_rst), .rdata(f906_rdata));
  assign f906_clk = clk;
  assign f906_rst = rst;
  // Bindings to f906

  // f908
  logic [0:0] f908_wen;
  logic [31:0] f908_wdata;
  logic [0:0] f908_clk;
  logic [0:0] f908_rst;
  logic [31:0] f908_rdata;
  sr_buffer_32_1 f908(.wen(f908_wen), .wdata(f908_wdata), .clk(f908_clk), .rst(f908_rst), .rdata(f908_rdata));
  assign f908_clk = clk;
  assign f908_rst = rst;
  // Bindings to f908

  // f910
  logic [0:0] f910_wen;
  logic [31:0] f910_wdata;
  logic [0:0] f910_clk;
  logic [0:0] f910_rst;
  logic [31:0] f910_rdata;
  sr_buffer_32_1 f910(.wen(f910_wen), .wdata(f910_wdata), .clk(f910_clk), .rst(f910_rst), .rdata(f910_rdata));
  assign f910_clk = clk;
  assign f910_rst = rst;
  // Bindings to f910

  // f912
  logic [0:0] f912_wen;
  logic [31:0] f912_wdata;
  logic [0:0] f912_clk;
  logic [0:0] f912_rst;
  logic [31:0] f912_rdata;
  sr_buffer_32_1 f912(.wen(f912_wen), .wdata(f912_wdata), .clk(f912_clk), .rst(f912_rst), .rdata(f912_rdata));
  assign f912_clk = clk;
  assign f912_rst = rst;
  // Bindings to f912

  // f914
  logic [0:0] f914_wen;
  logic [31:0] f914_wdata;
  logic [0:0] f914_clk;
  logic [0:0] f914_rst;
  logic [31:0] f914_rdata;
  sr_buffer_32_1 f914(.wen(f914_wen), .wdata(f914_wdata), .clk(f914_clk), .rst(f914_rst), .rdata(f914_rdata));
  assign f914_clk = clk;
  assign f914_rst = rst;
  // Bindings to f914

  // f916
  logic [0:0] f916_wen;
  logic [31:0] f916_wdata;
  logic [0:0] f916_clk;
  logic [0:0] f916_rst;
  logic [31:0] f916_rdata;
  sr_buffer_32_1 f916(.wen(f916_wen), .wdata(f916_wdata), .clk(f916_clk), .rst(f916_rst), .rdata(f916_rdata));
  assign f916_clk = clk;
  assign f916_rst = rst;
  // Bindings to f916

  // f918
  logic [0:0] f918_wen;
  logic [31:0] f918_wdata;
  logic [0:0] f918_clk;
  logic [0:0] f918_rst;
  logic [31:0] f918_rdata;
  sr_buffer_32_1 f918(.wen(f918_wen), .wdata(f918_wdata), .clk(f918_clk), .rst(f918_rst), .rdata(f918_rdata));
  assign f918_clk = clk;
  assign f918_rst = rst;
  // Bindings to f918

  // f920
  logic [0:0] f920_wen;
  logic [31:0] f920_wdata;
  logic [0:0] f920_clk;
  logic [0:0] f920_rst;
  logic [31:0] f920_rdata;
  sr_buffer_32_1 f920(.wen(f920_wen), .wdata(f920_wdata), .clk(f920_clk), .rst(f920_rst), .rdata(f920_rdata));
  assign f920_clk = clk;
  assign f920_rst = rst;
  // Bindings to f920

  // f922
  logic [0:0] f922_wen;
  logic [31:0] f922_wdata;
  logic [0:0] f922_clk;
  logic [0:0] f922_rst;
  logic [31:0] f922_rdata;
  sr_buffer_32_1 f922(.wen(f922_wen), .wdata(f922_wdata), .clk(f922_clk), .rst(f922_rst), .rdata(f922_rdata));
  assign f922_clk = clk;
  assign f922_rst = rst;
  // Bindings to f922

  // f924
  logic [0:0] f924_wen;
  logic [31:0] f924_wdata;
  logic [0:0] f924_clk;
  logic [0:0] f924_rst;
  logic [31:0] f924_rdata;
  sr_buffer_32_1 f924(.wen(f924_wen), .wdata(f924_wdata), .clk(f924_clk), .rst(f924_rst), .rdata(f924_rdata));
  assign f924_clk = clk;
  assign f924_rst = rst;
  // Bindings to f924

  // f926
  logic [0:0] f926_wen;
  logic [31:0] f926_wdata;
  logic [0:0] f926_clk;
  logic [0:0] f926_rst;
  logic [31:0] f926_rdata;
  sr_buffer_32_1 f926(.wen(f926_wen), .wdata(f926_wdata), .clk(f926_clk), .rst(f926_rst), .rdata(f926_rdata));
  assign f926_clk = clk;
  assign f926_rst = rst;
  // Bindings to f926

  // f928
  logic [0:0] f928_wen;
  logic [31:0] f928_wdata;
  logic [0:0] f928_clk;
  logic [0:0] f928_rst;
  logic [31:0] f928_rdata;
  sr_buffer_32_1 f928(.wen(f928_wen), .wdata(f928_wdata), .clk(f928_clk), .rst(f928_rst), .rdata(f928_rdata));
  assign f928_clk = clk;
  assign f928_rst = rst;
  // Bindings to f928

  // f930
  logic [0:0] f930_wen;
  logic [31:0] f930_wdata;
  logic [0:0] f930_clk;
  logic [0:0] f930_rst;
  logic [31:0] f930_rdata;
  sr_buffer_32_1 f930(.wen(f930_wen), .wdata(f930_wdata), .clk(f930_clk), .rst(f930_rst), .rdata(f930_rdata));
  assign f930_clk = clk;
  assign f930_rst = rst;
  // Bindings to f930

  // f932
  logic [0:0] f932_wen;
  logic [31:0] f932_wdata;
  logic [0:0] f932_clk;
  logic [0:0] f932_rst;
  logic [31:0] f932_rdata;
  sr_buffer_32_1 f932(.wen(f932_wen), .wdata(f932_wdata), .clk(f932_clk), .rst(f932_rst), .rdata(f932_rdata));
  assign f932_clk = clk;
  assign f932_rst = rst;
  // Bindings to f932

  // f934
  logic [0:0] f934_wen;
  logic [31:0] f934_wdata;
  logic [0:0] f934_clk;
  logic [0:0] f934_rst;
  logic [31:0] f934_rdata;
  sr_buffer_32_1 f934(.wen(f934_wen), .wdata(f934_wdata), .clk(f934_clk), .rst(f934_rst), .rdata(f934_rdata));
  assign f934_clk = clk;
  assign f934_rst = rst;
  // Bindings to f934

  // f936
  logic [0:0] f936_wen;
  logic [31:0] f936_wdata;
  logic [0:0] f936_clk;
  logic [0:0] f936_rst;
  logic [31:0] f936_rdata;
  sr_buffer_32_1 f936(.wen(f936_wen), .wdata(f936_wdata), .clk(f936_clk), .rst(f936_rst), .rdata(f936_rdata));
  assign f936_clk = clk;
  assign f936_rst = rst;
  // Bindings to f936

  // f938
  logic [0:0] f938_wen;
  logic [31:0] f938_wdata;
  logic [0:0] f938_clk;
  logic [0:0] f938_rst;
  logic [31:0] f938_rdata;
  sr_buffer_32_1 f938(.wen(f938_wen), .wdata(f938_wdata), .clk(f938_clk), .rst(f938_rst), .rdata(f938_rdata));
  assign f938_clk = clk;
  assign f938_rst = rst;
  // Bindings to f938

  // f844
  logic [0:0] f844_wen;
  logic [31:0] f844_wdata;
  logic [0:0] f844_clk;
  logic [0:0] f844_rst;
  logic [31:0] f844_rdata;
  sr_buffer_32_1 f844(.wen(f844_wen), .wdata(f844_wdata), .clk(f844_clk), .rst(f844_rst), .rdata(f844_rdata));
  assign f844_clk = clk;
  assign f844_rst = rst;
  // Bindings to f844

  // f710
  logic [0:0] f710_wen;
  logic [31:0] f710_wdata;
  logic [0:0] f710_clk;
  logic [0:0] f710_rst;
  logic [31:0] f710_rdata;
  sr_buffer_32_1 f710(.wen(f710_wen), .wdata(f710_wdata), .clk(f710_clk), .rst(f710_rst), .rdata(f710_rdata));
  assign f710_clk = clk;
  assign f710_rst = rst;
  // Bindings to f710

  // f712
  logic [0:0] f712_wen;
  logic [31:0] f712_wdata;
  logic [0:0] f712_clk;
  logic [0:0] f712_rst;
  logic [31:0] f712_rdata;
  sr_buffer_32_1 f712(.wen(f712_wen), .wdata(f712_wdata), .clk(f712_clk), .rst(f712_rst), .rdata(f712_rdata));
  assign f712_clk = clk;
  assign f712_rst = rst;
  // Bindings to f712

  // f850
  logic [0:0] f850_wen;
  logic [31:0] f850_wdata;
  logic [0:0] f850_clk;
  logic [0:0] f850_rst;
  logic [31:0] f850_rdata;
  sr_buffer_32_1 f850(.wen(f850_wen), .wdata(f850_wdata), .clk(f850_clk), .rst(f850_rst), .rdata(f850_rdata));
  assign f850_clk = clk;
  assign f850_rst = rst;
  // Bindings to f850

  // f716
  logic [0:0] f716_wen;
  logic [31:0] f716_wdata;
  logic [0:0] f716_clk;
  logic [0:0] f716_rst;
  logic [31:0] f716_rdata;
  sr_buffer_32_1 f716(.wen(f716_wen), .wdata(f716_wdata), .clk(f716_clk), .rst(f716_rst), .rdata(f716_rdata));
  assign f716_clk = clk;
  assign f716_rst = rst;
  // Bindings to f716

  // f720
  logic [0:0] f720_wen;
  logic [31:0] f720_wdata;
  logic [0:0] f720_clk;
  logic [0:0] f720_rst;
  logic [31:0] f720_rdata;
  sr_buffer_32_1 f720(.wen(f720_wen), .wdata(f720_wdata), .clk(f720_clk), .rst(f720_rst), .rdata(f720_rdata));
  assign f720_clk = clk;
  assign f720_rst = rst;
  // Bindings to f720

  // f842
  logic [0:0] f842_wen;
  logic [31:0] f842_wdata;
  logic [0:0] f842_clk;
  logic [0:0] f842_rst;
  logic [31:0] f842_rdata;
  sr_buffer_32_1 f842(.wen(f842_wen), .wdata(f842_wdata), .clk(f842_clk), .rst(f842_rst), .rdata(f842_rdata));
  assign f842_clk = clk;
  assign f842_rst = rst;
  // Bindings to f842

  // f718
  logic [0:0] f718_wen;
  logic [31:0] f718_wdata;
  logic [0:0] f718_clk;
  logic [0:0] f718_rst;
  logic [31:0] f718_rdata;
  sr_buffer_32_1 f718(.wen(f718_wen), .wdata(f718_wdata), .clk(f718_clk), .rst(f718_rst), .rdata(f718_rdata));
  assign f718_clk = clk;
  assign f718_rst = rst;
  // Bindings to f718

  // f714
  logic [0:0] f714_wen;
  logic [31:0] f714_wdata;
  logic [0:0] f714_clk;
  logic [0:0] f714_rst;
  logic [31:0] f714_rdata;
  sr_buffer_32_1 f714(.wen(f714_wen), .wdata(f714_wdata), .clk(f714_clk), .rst(f714_rst), .rdata(f714_rdata));
  assign f714_clk = clk;
  assign f714_rst = rst;
  // Bindings to f714

  // f708
  logic [0:0] f708_wen;
  logic [31:0] f708_wdata;
  logic [0:0] f708_clk;
  logic [0:0] f708_rst;
  logic [31:0] f708_rdata;
  sr_buffer_32_1 f708(.wen(f708_wen), .wdata(f708_wdata), .clk(f708_clk), .rst(f708_rst), .rdata(f708_rdata));
  assign f708_clk = clk;
  assign f708_rst = rst;
  // Bindings to f708



endmodule


module bright_weights_normed_gauss_blur_1_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1265;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_1_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_1_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2527;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_1_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1264;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_1_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_1_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_weights_normed_update_0_write_wen(output [0:0] bright_weights_normed_update_0_write_wen);

endmodule


module bright_weights_normed_gauss_blur_1_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (1259 - d0 >= 0) ? (1263) : (-1260 + d0 == 0) ? (1263) : 0;
    end
  end

endmodule


module out_wire_bright_weights_normed_gauss_blur_1_update_0_read_rdata(input [287:0] bright_weights_normed_gauss_blur_1_update_0_read_rdata);

endmodule


module bright_weights_normed(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_weights_normed_update_0_write_wen, input [31:0] fused_level_0_update_0_read_dummy, output [287:0] bright_weights_normed_gauss_blur_1_update_0_read_rdata, input [31:0] bright_weights_normed_update_0_write_wdata, input [287:0] bright_weights_normed_gauss_blur_1_update_0_read_dummy, output [31:0] fused_level_0_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_4;
  logic [31:0] rd_1;
  logic [287:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_4_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_4_stage_1 <= rd_4;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_clk;
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_rst;
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_start;
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_done;
  bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9 bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9(.clk(bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_clk), .rst(bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_rst), .start(bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_start), .done(bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_done));
  assign bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_clk = clk;
  assign bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9_rst = rst;
  // Bindings to bright_weights_normed_bright_weights_normed_update_0_write0_merged_banks_9

  // Bindings to bright_weights_normed_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_normed_update_0_write_wen;

  // selector_bright_weights_normed_gauss_blur_1_rd6_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd6_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd6_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd6_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd6_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd6_select_out;
  bright_weights_normed_gauss_blur_1_rd6_select selector_bright_weights_normed_gauss_blur_1_rd6_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd6_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd6_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd6_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd6_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd6_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd6_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd6_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd6_select

  // selector_bright_weights_normed_gauss_blur_1_rd5_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd5_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd5_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd5_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd5_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd5_select_out;
  bright_weights_normed_gauss_blur_1_rd5_select selector_bright_weights_normed_gauss_blur_1_rd5_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd5_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd5_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd5_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd5_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd5_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd5_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd5_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd5_select

  // selector_bright_weights_normed_gauss_blur_1_rd4_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd4_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd4_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd4_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd4_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd4_select_out;
  bright_weights_normed_gauss_blur_1_rd4_select selector_bright_weights_normed_gauss_blur_1_rd4_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd4_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd4_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd4_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd4_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd4_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd4_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd4_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd4_select

  // Bindings to fused_level_0_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_0_update_0_read_dummy;

  // Bindings to bright_weights_normed_gauss_blur_1_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_gauss_blur_1_update_0_read_rdata = rd_2;

  // Bindings to bright_weights_normed_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_normed_update_0_write_wdata;

  // selector_bright_weights_normed_gauss_blur_1_rd8_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd8_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd8_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd8_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd8_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd8_select_out;
  bright_weights_normed_gauss_blur_1_rd8_select selector_bright_weights_normed_gauss_blur_1_rd8_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd8_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd8_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd8_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd8_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd8_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd8_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd8_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd8_select

  // selector_bright_weights_normed_gauss_blur_1_rd7_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd7_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd7_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd7_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd7_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd7_select_out;
  bright_weights_normed_gauss_blur_1_rd7_select selector_bright_weights_normed_gauss_blur_1_rd7_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd7_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd7_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd7_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd7_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd7_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd7_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd7_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd7_select

  // selector_bright_weights_normed_gauss_blur_1_rd0_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd0_select_out;
  bright_weights_normed_gauss_blur_1_rd0_select selector_bright_weights_normed_gauss_blur_1_rd0_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd0_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd0_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd0_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd0_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd0_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd0_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd0_select

  // selector_fused_level_0_rd0_select
  logic [0:0] selector_fused_level_0_rd0_select_clk;
  logic [0:0] selector_fused_level_0_rd0_select_rst;
  logic [31:0] selector_fused_level_0_rd0_select_d0;
  logic [31:0] selector_fused_level_0_rd0_select_d1;
  logic [31:0] selector_fused_level_0_rd0_select_out;
  fused_level_0_rd0_select selector_fused_level_0_rd0_select(.clk(selector_fused_level_0_rd0_select_clk), .rst(selector_fused_level_0_rd0_select_rst), .d0(selector_fused_level_0_rd0_select_d0), .d1(selector_fused_level_0_rd0_select_d1), .out(selector_fused_level_0_rd0_select_out));
  assign selector_fused_level_0_rd0_select_clk = clk;
  assign selector_fused_level_0_rd0_select_rst = rst;
  // Bindings to selector_fused_level_0_rd0_select

  // selector_bright_weights_normed_gauss_blur_1_rd3_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd3_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd3_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd3_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd3_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd3_select_out;
  bright_weights_normed_gauss_blur_1_rd3_select selector_bright_weights_normed_gauss_blur_1_rd3_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd3_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd3_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd3_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd3_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd3_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd3_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd3_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd3_select

  // selector_bright_weights_normed_gauss_blur_1_rd2_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd2_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd2_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd2_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd2_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd2_select_out;
  bright_weights_normed_gauss_blur_1_rd2_select selector_bright_weights_normed_gauss_blur_1_rd2_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd2_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd2_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd2_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd2_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd2_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd2_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd2_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd2_select

  // selector_bright_weights_normed_gauss_blur_1_rd1_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd1_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_1_rd1_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd1_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd1_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_1_rd1_select_out;
  bright_weights_normed_gauss_blur_1_rd1_select selector_bright_weights_normed_gauss_blur_1_rd1_select(.clk(selector_bright_weights_normed_gauss_blur_1_rd1_select_clk), .rst(selector_bright_weights_normed_gauss_blur_1_rd1_select_rst), .d0(selector_bright_weights_normed_gauss_blur_1_rd1_select_d0), .d1(selector_bright_weights_normed_gauss_blur_1_rd1_select_d1), .out(selector_bright_weights_normed_gauss_blur_1_rd1_select_out));
  assign selector_bright_weights_normed_gauss_blur_1_rd1_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_1_rd1_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_1_rd1_select

  // bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_clk;
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_rst;
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_start;
  logic [0:0] bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_done;
  bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0 bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0(.clk(bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_clk), .rst(bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_rst), .start(bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_start), .done(bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_done));
  assign bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_clk = clk;
  assign bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0_rst = rst;
  // Bindings to bright_weights_normed_bright_weights_normed_update_0_write0_to_fused_level_0_rd0

  // Bindings to bright_weights_normed_gauss_blur_1_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_gauss_blur_1_update_0_read_dummy;

  // Bindings to fused_level_0_update_0_read_rdata
    // wr_5
  assign fused_level_0_update_0_read_rdata = rd_4;



endmodule


module in_wire_bright_weights_normed_update_0_write_wdata(output [31:0] bright_weights_normed_update_0_write_wdata);

endmodule


module in_wire_bright_weights_normed_gauss_blur_1_update_0_read_dummy(output [287:0] bright_weights_normed_gauss_blur_1_update_0_read_dummy);

endmodule


module bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module bright_weights_normed_gauss_ds_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_weights_normed_gauss_blur_1_update_0_write_wen(output [0:0] bright_weights_normed_gauss_blur_1_update_0_write_wen);

endmodule


module in_wire_bright_weights_normed_gauss_blur_1_update_0_write_wdata(output [31:0] bright_weights_normed_gauss_blur_1_update_0_write_wdata);

endmodule


module bright_weights_normed_gauss_blur_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] bright_weights_normed_gauss_ds_1_update_0_read_rdata, input [31:0] bright_weights_normed_gauss_ds_1_update_0_read_dummy, input [31:0] bright_weights_normed_gauss_blur_1_update_0_write_wdata, input [0:0] bright_weights_normed_gauss_blur_1_update_0_write_wen);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to bright_weights_normed_gauss_ds_1_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_gauss_ds_1_update_0_read_rdata = rd_2;

  // bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1
  logic [0:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_done;
  bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1 bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1(.clk(bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_clk), .rst(bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_rst), .start(bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_start), .done(bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_done));
  assign bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_clk = clk;
  assign bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1

  // Bindings to bright_weights_normed_gauss_ds_1_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_gauss_ds_1_update_0_read_dummy;

  // Bindings to bright_weights_normed_gauss_blur_1_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_normed_gauss_blur_1_update_0_write_wdata;

  // selector_bright_weights_normed_gauss_ds_1_rd0_select
  logic [0:0] selector_bright_weights_normed_gauss_ds_1_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_ds_1_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_ds_1_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_ds_1_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_ds_1_rd0_select_out;
  bright_weights_normed_gauss_ds_1_rd0_select selector_bright_weights_normed_gauss_ds_1_rd0_select(.clk(selector_bright_weights_normed_gauss_ds_1_rd0_select_clk), .rst(selector_bright_weights_normed_gauss_ds_1_rd0_select_rst), .d0(selector_bright_weights_normed_gauss_ds_1_rd0_select_d0), .d1(selector_bright_weights_normed_gauss_ds_1_rd0_select_d1), .out(selector_bright_weights_normed_gauss_ds_1_rd0_select_out));
  assign selector_bright_weights_normed_gauss_ds_1_rd0_select_clk = clk;
  assign selector_bright_weights_normed_gauss_ds_1_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_ds_1_rd0_select

  // Bindings to bright_weights_normed_gauss_blur_1_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_normed_gauss_blur_1_update_0_write_wen;



endmodule


module in_wire_bright_weights_normed_gauss_ds_1_update_0_read_dummy(output [31:0] bright_weights_normed_gauss_ds_1_update_0_read_dummy);

endmodule


module out_wire_bright_weights_normed_gauss_ds_1_update_0_read_rdata(input [31:0] bright_weights_normed_gauss_ds_1_update_0_read_rdata);

endmodule


module in_wire_bright_weights_normed_gauss_blur_2_update_0_write_wen(output [0:0] bright_weights_normed_gauss_blur_2_update_0_write_wen);

endmodule


module bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module bright_weights_normed_gauss_ds_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_weights_normed_gauss_blur_2_update_0_write_wdata(output [31:0] bright_weights_normed_gauss_blur_2_update_0_write_wdata);

endmodule


module bright_weights_normed_gauss_blur_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_weights_normed_gauss_blur_3_update_0_write_wen, input [31:0] bright_weights_normed_gauss_ds_3_update_0_read_dummy, output [31:0] bright_weights_normed_gauss_ds_3_update_0_read_rdata, input [31:0] bright_weights_normed_gauss_blur_3_update_0_write_wdata);

  logic [31:0] rd_1;
  logic [31:0] rd_2;
  logic [0:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;
  reg [0:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1
  logic [0:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_done;
  bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1 bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1(.clk(bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_clk), .rst(bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_rst), .start(bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_start), .done(bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_done));
  assign bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_clk = clk;
  assign bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1

  // Bindings to bright_weights_normed_gauss_blur_3_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_normed_gauss_blur_3_update_0_write_wen;

  // selector_bright_weights_normed_gauss_ds_3_rd0_select
  logic [0:0] selector_bright_weights_normed_gauss_ds_3_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_ds_3_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_ds_3_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_ds_3_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_ds_3_rd0_select_out;
  bright_weights_normed_gauss_ds_3_rd0_select selector_bright_weights_normed_gauss_ds_3_rd0_select(.clk(selector_bright_weights_normed_gauss_ds_3_rd0_select_clk), .rst(selector_bright_weights_normed_gauss_ds_3_rd0_select_rst), .d0(selector_bright_weights_normed_gauss_ds_3_rd0_select_d0), .d1(selector_bright_weights_normed_gauss_ds_3_rd0_select_d1), .out(selector_bright_weights_normed_gauss_ds_3_rd0_select_out));
  assign selector_bright_weights_normed_gauss_ds_3_rd0_select_clk = clk;
  assign selector_bright_weights_normed_gauss_ds_3_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_ds_3_rd0_select

  // Bindings to bright_weights_normed_gauss_ds_3_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_gauss_ds_3_update_0_read_dummy;

  // Bindings to bright_weights_normed_gauss_ds_3_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_gauss_ds_3_update_0_read_rdata = rd_2;

  // Bindings to bright_weights_normed_gauss_blur_3_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_normed_gauss_blur_3_update_0_write_wdata;



endmodule


module in_wire_bright_weights_normed_gauss_ds_2_update_0_read_dummy(output [31:0] bright_weights_normed_gauss_ds_2_update_0_read_dummy);

endmodule


module out_wire_bright_weights_normed_gauss_ds_2_update_0_read_rdata(input [31:0] bright_weights_normed_gauss_ds_2_update_0_read_rdata);

endmodule


module bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_312 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_312 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16



endmodule


module bright_weights_normed_gauss_blur_3_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (311 - d0 >= 0) ? (630) : (-312 + d0 == 0) ? (630) : 0;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 632;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_3_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 317;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_3_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_3_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 631;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_3_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 316;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_3_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_3_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module in_wire_bright_weights_normed_gauss_ds_2_update_0_write_wen(output [0:0] bright_weights_normed_gauss_ds_2_update_0_write_wen);

endmodule


module bright_weights_normed_gauss_blur_3_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (311 - d0 >= 0) ? (315) : (-312 + d0 == 0) ? (315) : 0;
    end
  end

endmodule


module in_wire_bright_weights_normed_gauss_ds_2_update_0_write_wdata(output [31:0] bright_weights_normed_gauss_ds_2_update_0_write_wdata);

endmodule


module in_wire_bright_weights_normed_gauss_blur_3_update_0_read_dummy(output [287:0] bright_weights_normed_gauss_blur_3_update_0_read_dummy);

endmodule


module out_wire_bright_weights_normed_gauss_blur_3_update_0_read_rdata(input [287:0] bright_weights_normed_gauss_blur_3_update_0_read_rdata);

endmodule


module dark_dark_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_1260 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_1260 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16



endmodule


module dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_3790 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f314
  logic [0:0] f314_wen;
  logic [31:0] f314_wdata;
  logic [0:0] f314_clk;
  logic [0:0] f314_rst;
  logic [31:0] f314_rdata;
  sr_buffer_32_1 f314(.wen(f314_wen), .wdata(f314_wdata), .clk(f314_clk), .rst(f314_rst), .rdata(f314_rdata));
  assign f314_clk = clk;
  assign f314_rst = rst;
  // Bindings to f314

  // f316
  logic [0:0] f316_wen;
  logic [31:0] f316_wdata;
  logic [0:0] f316_clk;
  logic [0:0] f316_rst;
  logic [31:0] f316_rdata;
  sr_buffer_32_1 f316(.wen(f316_wen), .wdata(f316_wdata), .clk(f316_clk), .rst(f316_rst), .rdata(f316_rdata));
  assign f316_clk = clk;
  assign f316_rst = rst;
  // Bindings to f316

  // f318
  logic [0:0] f318_wen;
  logic [31:0] f318_wdata;
  logic [0:0] f318_clk;
  logic [0:0] f318_rst;
  logic [31:0] f318_rdata;
  sr_buffer_32_1 f318(.wen(f318_wen), .wdata(f318_wdata), .clk(f318_clk), .rst(f318_rst), .rdata(f318_rdata));
  assign f318_clk = clk;
  assign f318_rst = rst;
  // Bindings to f318

  // f320
  logic [0:0] f320_wen;
  logic [31:0] f320_wdata;
  logic [0:0] f320_clk;
  logic [0:0] f320_rst;
  logic [31:0] f320_rdata;
  sr_buffer_32_1 f320(.wen(f320_wen), .wdata(f320_wdata), .clk(f320_clk), .rst(f320_rst), .rdata(f320_rdata));
  assign f320_clk = clk;
  assign f320_rst = rst;
  // Bindings to f320

  // f322
  logic [0:0] f322_wen;
  logic [31:0] f322_wdata;
  logic [0:0] f322_clk;
  logic [0:0] f322_rst;
  logic [31:0] f322_rdata;
  sr_buffer_32_1 f322(.wen(f322_wen), .wdata(f322_wdata), .clk(f322_clk), .rst(f322_rst), .rdata(f322_rdata));
  assign f322_clk = clk;
  assign f322_rst = rst;
  // Bindings to f322

  // f324
  logic [0:0] f324_wen;
  logic [31:0] f324_wdata;
  logic [0:0] f324_clk;
  logic [0:0] f324_rst;
  logic [31:0] f324_rdata;
  sr_buffer_32_1 f324(.wen(f324_wen), .wdata(f324_wdata), .clk(f324_clk), .rst(f324_rst), .rdata(f324_rdata));
  assign f324_clk = clk;
  assign f324_rst = rst;
  // Bindings to f324

  // f326
  logic [0:0] f326_wen;
  logic [31:0] f326_wdata;
  logic [0:0] f326_clk;
  logic [0:0] f326_rst;
  logic [31:0] f326_rdata;
  sr_buffer_32_1 f326(.wen(f326_wen), .wdata(f326_wdata), .clk(f326_clk), .rst(f326_rst), .rdata(f326_rdata));
  assign f326_clk = clk;
  assign f326_rst = rst;
  // Bindings to f326

  // f328
  logic [0:0] f328_wen;
  logic [31:0] f328_wdata;
  logic [0:0] f328_clk;
  logic [0:0] f328_rst;
  logic [31:0] f328_rdata;
  sr_buffer_32_1 f328(.wen(f328_wen), .wdata(f328_wdata), .clk(f328_clk), .rst(f328_rst), .rdata(f328_rdata));
  assign f328_clk = clk;
  assign f328_rst = rst;
  // Bindings to f328

  // f330
  logic [0:0] f330_wen;
  logic [31:0] f330_wdata;
  logic [0:0] f330_clk;
  logic [0:0] f330_rst;
  logic [31:0] f330_rdata;
  sr_buffer_32_1 f330(.wen(f330_wen), .wdata(f330_wdata), .clk(f330_clk), .rst(f330_rst), .rdata(f330_rdata));
  assign f330_clk = clk;
  assign f330_rst = rst;
  // Bindings to f330

  // f332
  logic [0:0] f332_wen;
  logic [31:0] f332_wdata;
  logic [0:0] f332_clk;
  logic [0:0] f332_rst;
  logic [31:0] f332_rdata;
  sr_buffer_32_1 f332(.wen(f332_wen), .wdata(f332_wdata), .clk(f332_clk), .rst(f332_rst), .rdata(f332_rdata));
  assign f332_clk = clk;
  assign f332_rst = rst;
  // Bindings to f332

  // f334
  logic [0:0] f334_wen;
  logic [31:0] f334_wdata;
  logic [0:0] f334_clk;
  logic [0:0] f334_rst;
  logic [31:0] f334_rdata;
  sr_buffer_32_1 f334(.wen(f334_wen), .wdata(f334_wdata), .clk(f334_clk), .rst(f334_rst), .rdata(f334_rdata));
  assign f334_clk = clk;
  assign f334_rst = rst;
  // Bindings to f334

  // f336
  logic [0:0] f336_wen;
  logic [31:0] f336_wdata;
  logic [0:0] f336_clk;
  logic [0:0] f336_rst;
  logic [31:0] f336_rdata;
  sr_buffer_32_1 f336(.wen(f336_wen), .wdata(f336_wdata), .clk(f336_clk), .rst(f336_rst), .rdata(f336_rdata));
  assign f336_clk = clk;
  assign f336_rst = rst;
  // Bindings to f336

  // f338
  logic [0:0] f338_wen;
  logic [31:0] f338_wdata;
  logic [0:0] f338_clk;
  logic [0:0] f338_rst;
  logic [31:0] f338_rdata;
  sr_buffer_32_1 f338(.wen(f338_wen), .wdata(f338_wdata), .clk(f338_clk), .rst(f338_rst), .rdata(f338_rdata));
  assign f338_clk = clk;
  assign f338_rst = rst;
  // Bindings to f338

  // f340
  logic [0:0] f340_wen;
  logic [31:0] f340_wdata;
  logic [0:0] f340_clk;
  logic [0:0] f340_rst;
  logic [31:0] f340_rdata;
  sr_buffer_32_1 f340(.wen(f340_wen), .wdata(f340_wdata), .clk(f340_clk), .rst(f340_rst), .rdata(f340_rdata));
  assign f340_clk = clk;
  assign f340_rst = rst;
  // Bindings to f340

  // f342
  logic [0:0] f342_wen;
  logic [31:0] f342_wdata;
  logic [0:0] f342_clk;
  logic [0:0] f342_rst;
  logic [31:0] f342_rdata;
  sr_buffer_32_1 f342(.wen(f342_wen), .wdata(f342_wdata), .clk(f342_clk), .rst(f342_rst), .rdata(f342_rdata));
  assign f342_clk = clk;
  assign f342_rst = rst;
  // Bindings to f342

  // f344
  logic [0:0] f344_wen;
  logic [31:0] f344_wdata;
  logic [0:0] f344_clk;
  logic [0:0] f344_rst;
  logic [31:0] f344_rdata;
  sr_buffer_32_1 f344(.wen(f344_wen), .wdata(f344_wdata), .clk(f344_clk), .rst(f344_rst), .rdata(f344_rdata));
  assign f344_clk = clk;
  assign f344_rst = rst;
  // Bindings to f344

  // f346
  logic [0:0] f346_wen;
  logic [31:0] f346_wdata;
  logic [0:0] f346_clk;
  logic [0:0] f346_rst;
  logic [31:0] f346_rdata;
  sr_buffer_32_1 f346(.wen(f346_wen), .wdata(f346_wdata), .clk(f346_clk), .rst(f346_rst), .rdata(f346_rdata));
  assign f346_clk = clk;
  assign f346_rst = rst;
  // Bindings to f346

  // f348
  logic [0:0] f348_wen;
  logic [31:0] f348_wdata;
  logic [0:0] f348_clk;
  logic [0:0] f348_rst;
  logic [31:0] f348_rdata;
  sr_buffer_32_1 f348(.wen(f348_wen), .wdata(f348_wdata), .clk(f348_clk), .rst(f348_rst), .rdata(f348_rdata));
  assign f348_clk = clk;
  assign f348_rst = rst;
  // Bindings to f348

  // f350
  logic [0:0] f350_wen;
  logic [31:0] f350_wdata;
  logic [0:0] f350_clk;
  logic [0:0] f350_rst;
  logic [31:0] f350_rdata;
  sr_buffer_32_1 f350(.wen(f350_wen), .wdata(f350_wdata), .clk(f350_clk), .rst(f350_rst), .rdata(f350_rdata));
  assign f350_clk = clk;
  assign f350_rst = rst;
  // Bindings to f350

  // f352
  logic [0:0] f352_wen;
  logic [31:0] f352_wdata;
  logic [0:0] f352_clk;
  logic [0:0] f352_rst;
  logic [31:0] f352_rdata;
  sr_buffer_32_1 f352(.wen(f352_wen), .wdata(f352_wdata), .clk(f352_clk), .rst(f352_rst), .rdata(f352_rdata));
  assign f352_clk = clk;
  assign f352_rst = rst;
  // Bindings to f352

  // f354
  logic [0:0] f354_wen;
  logic [31:0] f354_wdata;
  logic [0:0] f354_clk;
  logic [0:0] f354_rst;
  logic [31:0] f354_rdata;
  sr_buffer_32_1 f354(.wen(f354_wen), .wdata(f354_wdata), .clk(f354_clk), .rst(f354_rst), .rdata(f354_rdata));
  assign f354_clk = clk;
  assign f354_rst = rst;
  // Bindings to f354

  // f356
  logic [0:0] f356_wen;
  logic [31:0] f356_wdata;
  logic [0:0] f356_clk;
  logic [0:0] f356_rst;
  logic [31:0] f356_rdata;
  sr_buffer_32_1 f356(.wen(f356_wen), .wdata(f356_wdata), .clk(f356_clk), .rst(f356_rst), .rdata(f356_rdata));
  assign f356_clk = clk;
  assign f356_rst = rst;
  // Bindings to f356

  // f358
  logic [0:0] f358_wen;
  logic [31:0] f358_wdata;
  logic [0:0] f358_clk;
  logic [0:0] f358_rst;
  logic [31:0] f358_rdata;
  sr_buffer_32_1 f358(.wen(f358_wen), .wdata(f358_wdata), .clk(f358_clk), .rst(f358_rst), .rdata(f358_rdata));
  assign f358_clk = clk;
  assign f358_rst = rst;
  // Bindings to f358

  // f360
  logic [0:0] f360_wen;
  logic [31:0] f360_wdata;
  logic [0:0] f360_clk;
  logic [0:0] f360_rst;
  logic [31:0] f360_rdata;
  sr_buffer_32_1 f360(.wen(f360_wen), .wdata(f360_wdata), .clk(f360_clk), .rst(f360_rst), .rdata(f360_rdata));
  assign f360_clk = clk;
  assign f360_rst = rst;
  // Bindings to f360

  // f362
  logic [0:0] f362_wen;
  logic [31:0] f362_wdata;
  logic [0:0] f362_clk;
  logic [0:0] f362_rst;
  logic [31:0] f362_rdata;
  sr_buffer_32_1 f362(.wen(f362_wen), .wdata(f362_wdata), .clk(f362_clk), .rst(f362_rst), .rdata(f362_rdata));
  assign f362_clk = clk;
  assign f362_rst = rst;
  // Bindings to f362

  // f364
  logic [0:0] f364_wen;
  logic [31:0] f364_wdata;
  logic [0:0] f364_clk;
  logic [0:0] f364_rst;
  logic [31:0] f364_rdata;
  sr_buffer_32_1 f364(.wen(f364_wen), .wdata(f364_wdata), .clk(f364_clk), .rst(f364_rst), .rdata(f364_rdata));
  assign f364_clk = clk;
  assign f364_rst = rst;
  // Bindings to f364

  // f366
  logic [0:0] f366_wen;
  logic [31:0] f366_wdata;
  logic [0:0] f366_clk;
  logic [0:0] f366_rst;
  logic [31:0] f366_rdata;
  sr_buffer_32_1 f366(.wen(f366_wen), .wdata(f366_wdata), .clk(f366_clk), .rst(f366_rst), .rdata(f366_rdata));
  assign f366_clk = clk;
  assign f366_rst = rst;
  // Bindings to f366

  // f368
  logic [0:0] f368_wen;
  logic [31:0] f368_wdata;
  logic [0:0] f368_clk;
  logic [0:0] f368_rst;
  logic [31:0] f368_rdata;
  sr_buffer_32_1 f368(.wen(f368_wen), .wdata(f368_wdata), .clk(f368_clk), .rst(f368_rst), .rdata(f368_rdata));
  assign f368_clk = clk;
  assign f368_rst = rst;
  // Bindings to f368

  // f370
  logic [0:0] f370_wen;
  logic [31:0] f370_wdata;
  logic [0:0] f370_clk;
  logic [0:0] f370_rst;
  logic [31:0] f370_rdata;
  sr_buffer_32_1 f370(.wen(f370_wen), .wdata(f370_wdata), .clk(f370_clk), .rst(f370_rst), .rdata(f370_rdata));
  assign f370_clk = clk;
  assign f370_rst = rst;
  // Bindings to f370

  // f372
  logic [0:0] f372_wen;
  logic [31:0] f372_wdata;
  logic [0:0] f372_clk;
  logic [0:0] f372_rst;
  logic [31:0] f372_rdata;
  sr_buffer_32_1 f372(.wen(f372_wen), .wdata(f372_wdata), .clk(f372_clk), .rst(f372_rst), .rdata(f372_rdata));
  assign f372_clk = clk;
  assign f372_rst = rst;
  // Bindings to f372

  // f374
  logic [0:0] f374_wen;
  logic [31:0] f374_wdata;
  logic [0:0] f374_clk;
  logic [0:0] f374_rst;
  logic [31:0] f374_rdata;
  sr_buffer_32_1 f374(.wen(f374_wen), .wdata(f374_wdata), .clk(f374_clk), .rst(f374_rst), .rdata(f374_rdata));
  assign f374_clk = clk;
  assign f374_rst = rst;
  // Bindings to f374

  // f376
  logic [0:0] f376_wen;
  logic [31:0] f376_wdata;
  logic [0:0] f376_clk;
  logic [0:0] f376_rst;
  logic [31:0] f376_rdata;
  sr_buffer_32_1 f376(.wen(f376_wen), .wdata(f376_wdata), .clk(f376_clk), .rst(f376_rst), .rdata(f376_rdata));
  assign f376_clk = clk;
  assign f376_rst = rst;
  // Bindings to f376

  // f378
  logic [0:0] f378_wen;
  logic [31:0] f378_wdata;
  logic [0:0] f378_clk;
  logic [0:0] f378_rst;
  logic [31:0] f378_rdata;
  sr_buffer_32_1 f378(.wen(f378_wen), .wdata(f378_wdata), .clk(f378_clk), .rst(f378_rst), .rdata(f378_rdata));
  assign f378_clk = clk;
  assign f378_rst = rst;
  // Bindings to f378

  // f380
  logic [0:0] f380_wen;
  logic [31:0] f380_wdata;
  logic [0:0] f380_clk;
  logic [0:0] f380_rst;
  logic [31:0] f380_rdata;
  sr_buffer_32_1 f380(.wen(f380_wen), .wdata(f380_wdata), .clk(f380_clk), .rst(f380_rst), .rdata(f380_rdata));
  assign f380_clk = clk;
  assign f380_rst = rst;
  // Bindings to f380

  // f382
  logic [0:0] f382_wen;
  logic [31:0] f382_wdata;
  logic [0:0] f382_clk;
  logic [0:0] f382_rst;
  logic [31:0] f382_rdata;
  sr_buffer_32_1 f382(.wen(f382_wen), .wdata(f382_wdata), .clk(f382_clk), .rst(f382_rst), .rdata(f382_rdata));
  assign f382_clk = clk;
  assign f382_rst = rst;
  // Bindings to f382

  // f384
  logic [0:0] f384_wen;
  logic [31:0] f384_wdata;
  logic [0:0] f384_clk;
  logic [0:0] f384_rst;
  logic [31:0] f384_rdata;
  sr_buffer_32_1 f384(.wen(f384_wen), .wdata(f384_wdata), .clk(f384_clk), .rst(f384_rst), .rdata(f384_rdata));
  assign f384_clk = clk;
  assign f384_rst = rst;
  // Bindings to f384

  // f386
  logic [0:0] f386_wen;
  logic [31:0] f386_wdata;
  logic [0:0] f386_clk;
  logic [0:0] f386_rst;
  logic [31:0] f386_rdata;
  sr_buffer_32_1 f386(.wen(f386_wen), .wdata(f386_wdata), .clk(f386_clk), .rst(f386_rst), .rdata(f386_rdata));
  assign f386_clk = clk;
  assign f386_rst = rst;
  // Bindings to f386

  // f388
  logic [0:0] f388_wen;
  logic [31:0] f388_wdata;
  logic [0:0] f388_clk;
  logic [0:0] f388_rst;
  logic [31:0] f388_rdata;
  sr_buffer_32_1 f388(.wen(f388_wen), .wdata(f388_wdata), .clk(f388_clk), .rst(f388_rst), .rdata(f388_rdata));
  assign f388_clk = clk;
  assign f388_rst = rst;
  // Bindings to f388

  // f390
  logic [0:0] f390_wen;
  logic [31:0] f390_wdata;
  logic [0:0] f390_clk;
  logic [0:0] f390_rst;
  logic [31:0] f390_rdata;
  sr_buffer_32_1 f390(.wen(f390_wen), .wdata(f390_wdata), .clk(f390_clk), .rst(f390_rst), .rdata(f390_rdata));
  assign f390_clk = clk;
  assign f390_rst = rst;
  // Bindings to f390

  // f392
  logic [0:0] f392_wen;
  logic [31:0] f392_wdata;
  logic [0:0] f392_clk;
  logic [0:0] f392_rst;
  logic [31:0] f392_rdata;
  sr_buffer_32_1 f392(.wen(f392_wen), .wdata(f392_wdata), .clk(f392_clk), .rst(f392_rst), .rdata(f392_rdata));
  assign f392_clk = clk;
  assign f392_rst = rst;
  // Bindings to f392

  // f394
  logic [0:0] f394_wen;
  logic [31:0] f394_wdata;
  logic [0:0] f394_clk;
  logic [0:0] f394_rst;
  logic [31:0] f394_rdata;
  sr_buffer_32_1 f394(.wen(f394_wen), .wdata(f394_wdata), .clk(f394_clk), .rst(f394_rst), .rdata(f394_rdata));
  assign f394_clk = clk;
  assign f394_rst = rst;
  // Bindings to f394

  // f396
  logic [0:0] f396_wen;
  logic [31:0] f396_wdata;
  logic [0:0] f396_clk;
  logic [0:0] f396_rst;
  logic [31:0] f396_rdata;
  sr_buffer_32_1 f396(.wen(f396_wen), .wdata(f396_wdata), .clk(f396_clk), .rst(f396_rst), .rdata(f396_rdata));
  assign f396_clk = clk;
  assign f396_rst = rst;
  // Bindings to f396

  // f398
  logic [0:0] f398_wen;
  logic [31:0] f398_wdata;
  logic [0:0] f398_clk;
  logic [0:0] f398_rst;
  logic [31:0] f398_rdata;
  sr_buffer_32_1 f398(.wen(f398_wen), .wdata(f398_wdata), .clk(f398_clk), .rst(f398_rst), .rdata(f398_rdata));
  assign f398_clk = clk;
  assign f398_rst = rst;
  // Bindings to f398

  // f400
  logic [0:0] f400_wen;
  logic [31:0] f400_wdata;
  logic [0:0] f400_clk;
  logic [0:0] f400_rst;
  logic [31:0] f400_rdata;
  sr_buffer_32_1 f400(.wen(f400_wen), .wdata(f400_wdata), .clk(f400_clk), .rst(f400_rst), .rdata(f400_rdata));
  assign f400_clk = clk;
  assign f400_rst = rst;
  // Bindings to f400

  // f402
  logic [0:0] f402_wen;
  logic [31:0] f402_wdata;
  logic [0:0] f402_clk;
  logic [0:0] f402_rst;
  logic [31:0] f402_rdata;
  sr_buffer_32_1 f402(.wen(f402_wen), .wdata(f402_wdata), .clk(f402_clk), .rst(f402_rst), .rdata(f402_rdata));
  assign f402_clk = clk;
  assign f402_rst = rst;
  // Bindings to f402

  // f404
  logic [0:0] f404_wen;
  logic [31:0] f404_wdata;
  logic [0:0] f404_clk;
  logic [0:0] f404_rst;
  logic [31:0] f404_rdata;
  sr_buffer_32_1 f404(.wen(f404_wen), .wdata(f404_wdata), .clk(f404_clk), .rst(f404_rst), .rdata(f404_rdata));
  assign f404_clk = clk;
  assign f404_rst = rst;
  // Bindings to f404

  // f406
  logic [0:0] f406_wen;
  logic [31:0] f406_wdata;
  logic [0:0] f406_clk;
  logic [0:0] f406_rst;
  logic [31:0] f406_rdata;
  sr_buffer_32_1 f406(.wen(f406_wen), .wdata(f406_wdata), .clk(f406_clk), .rst(f406_rst), .rdata(f406_rdata));
  assign f406_clk = clk;
  assign f406_rst = rst;
  // Bindings to f406

  // f408
  logic [0:0] f408_wen;
  logic [31:0] f408_wdata;
  logic [0:0] f408_clk;
  logic [0:0] f408_rst;
  logic [31:0] f408_rdata;
  sr_buffer_32_1 f408(.wen(f408_wen), .wdata(f408_wdata), .clk(f408_clk), .rst(f408_rst), .rdata(f408_rdata));
  assign f408_clk = clk;
  assign f408_rst = rst;
  // Bindings to f408

  // f410
  logic [0:0] f410_wen;
  logic [31:0] f410_wdata;
  logic [0:0] f410_clk;
  logic [0:0] f410_rst;
  logic [31:0] f410_rdata;
  sr_buffer_32_1 f410(.wen(f410_wen), .wdata(f410_wdata), .clk(f410_clk), .rst(f410_rst), .rdata(f410_rdata));
  assign f410_clk = clk;
  assign f410_rst = rst;
  // Bindings to f410

  // f412
  logic [0:0] f412_wen;
  logic [31:0] f412_wdata;
  logic [0:0] f412_clk;
  logic [0:0] f412_rst;
  logic [31:0] f412_rdata;
  sr_buffer_32_1 f412(.wen(f412_wen), .wdata(f412_wdata), .clk(f412_clk), .rst(f412_rst), .rdata(f412_rdata));
  assign f412_clk = clk;
  assign f412_rst = rst;
  // Bindings to f412

  // f414
  logic [0:0] f414_wen;
  logic [31:0] f414_wdata;
  logic [0:0] f414_clk;
  logic [0:0] f414_rst;
  logic [31:0] f414_rdata;
  sr_buffer_32_1 f414(.wen(f414_wen), .wdata(f414_wdata), .clk(f414_clk), .rst(f414_rst), .rdata(f414_rdata));
  assign f414_clk = clk;
  assign f414_rst = rst;
  // Bindings to f414

  // f416
  logic [0:0] f416_wen;
  logic [31:0] f416_wdata;
  logic [0:0] f416_clk;
  logic [0:0] f416_rst;
  logic [31:0] f416_rdata;
  sr_buffer_32_1 f416(.wen(f416_wen), .wdata(f416_wdata), .clk(f416_clk), .rst(f416_rst), .rdata(f416_rdata));
  assign f416_clk = clk;
  assign f416_rst = rst;
  // Bindings to f416

  // f418
  logic [0:0] f418_wen;
  logic [31:0] f418_wdata;
  logic [0:0] f418_clk;
  logic [0:0] f418_rst;
  logic [31:0] f418_rdata;
  sr_buffer_32_1 f418(.wen(f418_wen), .wdata(f418_wdata), .clk(f418_clk), .rst(f418_rst), .rdata(f418_rdata));
  assign f418_clk = clk;
  assign f418_rst = rst;
  // Bindings to f418

  // f420
  logic [0:0] f420_wen;
  logic [31:0] f420_wdata;
  logic [0:0] f420_clk;
  logic [0:0] f420_rst;
  logic [31:0] f420_rdata;
  sr_buffer_32_1 f420(.wen(f420_wen), .wdata(f420_wdata), .clk(f420_clk), .rst(f420_rst), .rdata(f420_rdata));
  assign f420_clk = clk;
  assign f420_rst = rst;
  // Bindings to f420

  // f422
  logic [0:0] f422_wen;
  logic [31:0] f422_wdata;
  logic [0:0] f422_clk;
  logic [0:0] f422_rst;
  logic [31:0] f422_rdata;
  sr_buffer_32_1 f422(.wen(f422_wen), .wdata(f422_wdata), .clk(f422_clk), .rst(f422_rst), .rdata(f422_rdata));
  assign f422_clk = clk;
  assign f422_rst = rst;
  // Bindings to f422

  // f424
  logic [0:0] f424_wen;
  logic [31:0] f424_wdata;
  logic [0:0] f424_clk;
  logic [0:0] f424_rst;
  logic [31:0] f424_rdata;
  sr_buffer_32_1 f424(.wen(f424_wen), .wdata(f424_wdata), .clk(f424_clk), .rst(f424_rst), .rdata(f424_rdata));
  assign f424_clk = clk;
  assign f424_rst = rst;
  // Bindings to f424

  // f426
  logic [0:0] f426_wen;
  logic [31:0] f426_wdata;
  logic [0:0] f426_clk;
  logic [0:0] f426_rst;
  logic [31:0] f426_rdata;
  sr_buffer_32_1 f426(.wen(f426_wen), .wdata(f426_wdata), .clk(f426_clk), .rst(f426_rst), .rdata(f426_rdata));
  assign f426_clk = clk;
  assign f426_rst = rst;
  // Bindings to f426

  // f428
  logic [0:0] f428_wen;
  logic [31:0] f428_wdata;
  logic [0:0] f428_clk;
  logic [0:0] f428_rst;
  logic [31:0] f428_rdata;
  sr_buffer_32_1 f428(.wen(f428_wen), .wdata(f428_wdata), .clk(f428_clk), .rst(f428_rst), .rdata(f428_rdata));
  assign f428_clk = clk;
  assign f428_rst = rst;
  // Bindings to f428

  // f430
  logic [0:0] f430_wen;
  logic [31:0] f430_wdata;
  logic [0:0] f430_clk;
  logic [0:0] f430_rst;
  logic [31:0] f430_rdata;
  sr_buffer_32_1 f430(.wen(f430_wen), .wdata(f430_wdata), .clk(f430_clk), .rst(f430_rst), .rdata(f430_rdata));
  assign f430_clk = clk;
  assign f430_rst = rst;
  // Bindings to f430

  // f432
  logic [0:0] f432_wen;
  logic [31:0] f432_wdata;
  logic [0:0] f432_clk;
  logic [0:0] f432_rst;
  logic [31:0] f432_rdata;
  sr_buffer_32_1 f432(.wen(f432_wen), .wdata(f432_wdata), .clk(f432_clk), .rst(f432_rst), .rdata(f432_rdata));
  assign f432_clk = clk;
  assign f432_rst = rst;
  // Bindings to f432

  // f434
  logic [0:0] f434_wen;
  logic [31:0] f434_wdata;
  logic [0:0] f434_clk;
  logic [0:0] f434_rst;
  logic [31:0] f434_rdata;
  sr_buffer_32_1 f434(.wen(f434_wen), .wdata(f434_wdata), .clk(f434_clk), .rst(f434_rst), .rdata(f434_rdata));
  assign f434_clk = clk;
  assign f434_rst = rst;
  // Bindings to f434

  // f436
  logic [0:0] f436_wen;
  logic [31:0] f436_wdata;
  logic [0:0] f436_clk;
  logic [0:0] f436_rst;
  logic [31:0] f436_rdata;
  sr_buffer_32_1 f436(.wen(f436_wen), .wdata(f436_wdata), .clk(f436_clk), .rst(f436_rst), .rdata(f436_rdata));
  assign f436_clk = clk;
  assign f436_rst = rst;
  // Bindings to f436

  // f438
  logic [0:0] f438_wen;
  logic [31:0] f438_wdata;
  logic [0:0] f438_clk;
  logic [0:0] f438_rst;
  logic [31:0] f438_rdata;
  sr_buffer_32_1 f438(.wen(f438_wen), .wdata(f438_wdata), .clk(f438_clk), .rst(f438_rst), .rdata(f438_rdata));
  assign f438_clk = clk;
  assign f438_rst = rst;
  // Bindings to f438

  // f440
  logic [0:0] f440_wen;
  logic [31:0] f440_wdata;
  logic [0:0] f440_clk;
  logic [0:0] f440_rst;
  logic [31:0] f440_rdata;
  sr_buffer_32_1 f440(.wen(f440_wen), .wdata(f440_wdata), .clk(f440_clk), .rst(f440_rst), .rdata(f440_rdata));
  assign f440_clk = clk;
  assign f440_rst = rst;
  // Bindings to f440

  // f442
  logic [0:0] f442_wen;
  logic [31:0] f442_wdata;
  logic [0:0] f442_clk;
  logic [0:0] f442_rst;
  logic [31:0] f442_rdata;
  sr_buffer_32_1 f442(.wen(f442_wen), .wdata(f442_wdata), .clk(f442_clk), .rst(f442_rst), .rdata(f442_rdata));
  assign f442_clk = clk;
  assign f442_rst = rst;
  // Bindings to f442

  // f444
  logic [0:0] f444_wen;
  logic [31:0] f444_wdata;
  logic [0:0] f444_clk;
  logic [0:0] f444_rst;
  logic [31:0] f444_rdata;
  sr_buffer_32_1 f444(.wen(f444_wen), .wdata(f444_wdata), .clk(f444_clk), .rst(f444_rst), .rdata(f444_rdata));
  assign f444_clk = clk;
  assign f444_rst = rst;
  // Bindings to f444

  // f446
  logic [0:0] f446_wen;
  logic [31:0] f446_wdata;
  logic [0:0] f446_clk;
  logic [0:0] f446_rst;
  logic [31:0] f446_rdata;
  sr_buffer_32_1 f446(.wen(f446_wen), .wdata(f446_wdata), .clk(f446_clk), .rst(f446_rst), .rdata(f446_rdata));
  assign f446_clk = clk;
  assign f446_rst = rst;
  // Bindings to f446

  // f448
  logic [0:0] f448_wen;
  logic [31:0] f448_wdata;
  logic [0:0] f448_clk;
  logic [0:0] f448_rst;
  logic [31:0] f448_rdata;
  sr_buffer_32_1 f448(.wen(f448_wen), .wdata(f448_wdata), .clk(f448_clk), .rst(f448_rst), .rdata(f448_rdata));
  assign f448_clk = clk;
  assign f448_rst = rst;
  // Bindings to f448

  // f450
  logic [0:0] f450_wen;
  logic [31:0] f450_wdata;
  logic [0:0] f450_clk;
  logic [0:0] f450_rst;
  logic [31:0] f450_rdata;
  sr_buffer_32_1 f450(.wen(f450_wen), .wdata(f450_wdata), .clk(f450_clk), .rst(f450_rst), .rdata(f450_rdata));
  assign f450_clk = clk;
  assign f450_rst = rst;
  // Bindings to f450

  // f452
  logic [0:0] f452_wen;
  logic [31:0] f452_wdata;
  logic [0:0] f452_clk;
  logic [0:0] f452_rst;
  logic [31:0] f452_rdata;
  sr_buffer_32_1 f452(.wen(f452_wen), .wdata(f452_wdata), .clk(f452_clk), .rst(f452_rst), .rdata(f452_rdata));
  assign f452_clk = clk;
  assign f452_rst = rst;
  // Bindings to f452

  // f454
  logic [0:0] f454_wen;
  logic [31:0] f454_wdata;
  logic [0:0] f454_clk;
  logic [0:0] f454_rst;
  logic [31:0] f454_rdata;
  sr_buffer_32_1 f454(.wen(f454_wen), .wdata(f454_wdata), .clk(f454_clk), .rst(f454_rst), .rdata(f454_rdata));
  assign f454_clk = clk;
  assign f454_rst = rst;
  // Bindings to f454

  // f456
  logic [0:0] f456_wen;
  logic [31:0] f456_wdata;
  logic [0:0] f456_clk;
  logic [0:0] f456_rst;
  logic [31:0] f456_rdata;
  sr_buffer_32_1 f456(.wen(f456_wen), .wdata(f456_wdata), .clk(f456_clk), .rst(f456_rst), .rdata(f456_rdata));
  assign f456_clk = clk;
  assign f456_rst = rst;
  // Bindings to f456

  // f458
  logic [0:0] f458_wen;
  logic [31:0] f458_wdata;
  logic [0:0] f458_clk;
  logic [0:0] f458_rst;
  logic [31:0] f458_rdata;
  sr_buffer_32_1 f458(.wen(f458_wen), .wdata(f458_wdata), .clk(f458_clk), .rst(f458_rst), .rdata(f458_rdata));
  assign f458_clk = clk;
  assign f458_rst = rst;
  // Bindings to f458

  // f460
  logic [0:0] f460_wen;
  logic [31:0] f460_wdata;
  logic [0:0] f460_clk;
  logic [0:0] f460_rst;
  logic [31:0] f460_rdata;
  sr_buffer_32_1 f460(.wen(f460_wen), .wdata(f460_wdata), .clk(f460_clk), .rst(f460_rst), .rdata(f460_rdata));
  assign f460_clk = clk;
  assign f460_rst = rst;
  // Bindings to f460

  // f462
  logic [0:0] f462_wen;
  logic [31:0] f462_wdata;
  logic [0:0] f462_clk;
  logic [0:0] f462_rst;
  logic [31:0] f462_rdata;
  sr_buffer_32_1 f462(.wen(f462_wen), .wdata(f462_wdata), .clk(f462_clk), .rst(f462_rst), .rdata(f462_rdata));
  assign f462_clk = clk;
  assign f462_rst = rst;
  // Bindings to f462

  // f464
  logic [0:0] f464_wen;
  logic [31:0] f464_wdata;
  logic [0:0] f464_clk;
  logic [0:0] f464_rst;
  logic [31:0] f464_rdata;
  sr_buffer_32_1 f464(.wen(f464_wen), .wdata(f464_wdata), .clk(f464_clk), .rst(f464_rst), .rdata(f464_rdata));
  assign f464_clk = clk;
  assign f464_rst = rst;
  // Bindings to f464

  // f466
  logic [0:0] f466_wen;
  logic [31:0] f466_wdata;
  logic [0:0] f466_clk;
  logic [0:0] f466_rst;
  logic [31:0] f466_rdata;
  sr_buffer_32_1 f466(.wen(f466_wen), .wdata(f466_wdata), .clk(f466_clk), .rst(f466_rst), .rdata(f466_rdata));
  assign f466_clk = clk;
  assign f466_rst = rst;
  // Bindings to f466

  // f468
  logic [0:0] f468_wen;
  logic [31:0] f468_wdata;
  logic [0:0] f468_clk;
  logic [0:0] f468_rst;
  logic [31:0] f468_rdata;
  sr_buffer_32_1 f468(.wen(f468_wen), .wdata(f468_wdata), .clk(f468_clk), .rst(f468_rst), .rdata(f468_rdata));
  assign f468_clk = clk;
  assign f468_rst = rst;
  // Bindings to f468

  // f470
  logic [0:0] f470_wen;
  logic [31:0] f470_wdata;
  logic [0:0] f470_clk;
  logic [0:0] f470_rst;
  logic [31:0] f470_rdata;
  sr_buffer_32_1 f470(.wen(f470_wen), .wdata(f470_wdata), .clk(f470_clk), .rst(f470_rst), .rdata(f470_rdata));
  assign f470_clk = clk;
  assign f470_rst = rst;
  // Bindings to f470

  // f472
  logic [0:0] f472_wen;
  logic [31:0] f472_wdata;
  logic [0:0] f472_clk;
  logic [0:0] f472_rst;
  logic [31:0] f472_rdata;
  sr_buffer_32_1 f472(.wen(f472_wen), .wdata(f472_wdata), .clk(f472_clk), .rst(f472_rst), .rdata(f472_rdata));
  assign f472_clk = clk;
  assign f472_rst = rst;
  // Bindings to f472

  // f474
  logic [0:0] f474_wen;
  logic [31:0] f474_wdata;
  logic [0:0] f474_clk;
  logic [0:0] f474_rst;
  logic [31:0] f474_rdata;
  sr_buffer_32_1 f474(.wen(f474_wen), .wdata(f474_wdata), .clk(f474_clk), .rst(f474_rst), .rdata(f474_rdata));
  assign f474_clk = clk;
  assign f474_rst = rst;
  // Bindings to f474

  // f476
  logic [0:0] f476_wen;
  logic [31:0] f476_wdata;
  logic [0:0] f476_clk;
  logic [0:0] f476_rst;
  logic [31:0] f476_rdata;
  sr_buffer_32_1 f476(.wen(f476_wen), .wdata(f476_wdata), .clk(f476_clk), .rst(f476_rst), .rdata(f476_rdata));
  assign f476_clk = clk;
  assign f476_rst = rst;
  // Bindings to f476

  // f478
  logic [0:0] f478_wen;
  logic [31:0] f478_wdata;
  logic [0:0] f478_clk;
  logic [0:0] f478_rst;
  logic [31:0] f478_rdata;
  sr_buffer_32_1 f478(.wen(f478_wen), .wdata(f478_wdata), .clk(f478_clk), .rst(f478_rst), .rdata(f478_rdata));
  assign f478_clk = clk;
  assign f478_rst = rst;
  // Bindings to f478

  // f480
  logic [0:0] f480_wen;
  logic [31:0] f480_wdata;
  logic [0:0] f480_clk;
  logic [0:0] f480_rst;
  logic [31:0] f480_rdata;
  sr_buffer_32_1 f480(.wen(f480_wen), .wdata(f480_wdata), .clk(f480_clk), .rst(f480_rst), .rdata(f480_rdata));
  assign f480_clk = clk;
  assign f480_rst = rst;
  // Bindings to f480

  // f482
  logic [0:0] f482_wen;
  logic [31:0] f482_wdata;
  logic [0:0] f482_clk;
  logic [0:0] f482_rst;
  logic [31:0] f482_rdata;
  sr_buffer_32_1 f482(.wen(f482_wen), .wdata(f482_wdata), .clk(f482_clk), .rst(f482_rst), .rdata(f482_rdata));
  assign f482_clk = clk;
  assign f482_rst = rst;
  // Bindings to f482

  // f484
  logic [0:0] f484_wen;
  logic [31:0] f484_wdata;
  logic [0:0] f484_clk;
  logic [0:0] f484_rst;
  logic [31:0] f484_rdata;
  sr_buffer_32_1 f484(.wen(f484_wen), .wdata(f484_wdata), .clk(f484_clk), .rst(f484_rst), .rdata(f484_rdata));
  assign f484_clk = clk;
  assign f484_rst = rst;
  // Bindings to f484

  // f486
  logic [0:0] f486_wen;
  logic [31:0] f486_wdata;
  logic [0:0] f486_clk;
  logic [0:0] f486_rst;
  logic [31:0] f486_rdata;
  sr_buffer_32_1 f486(.wen(f486_wen), .wdata(f486_wdata), .clk(f486_clk), .rst(f486_rst), .rdata(f486_rdata));
  assign f486_clk = clk;
  assign f486_rst = rst;
  // Bindings to f486

  // f488
  logic [0:0] f488_wen;
  logic [31:0] f488_wdata;
  logic [0:0] f488_clk;
  logic [0:0] f488_rst;
  logic [31:0] f488_rdata;
  sr_buffer_32_1 f488(.wen(f488_wen), .wdata(f488_wdata), .clk(f488_clk), .rst(f488_rst), .rdata(f488_rdata));
  assign f488_clk = clk;
  assign f488_rst = rst;
  // Bindings to f488

  // f490
  logic [0:0] f490_wen;
  logic [31:0] f490_wdata;
  logic [0:0] f490_clk;
  logic [0:0] f490_rst;
  logic [31:0] f490_rdata;
  sr_buffer_32_1 f490(.wen(f490_wen), .wdata(f490_wdata), .clk(f490_clk), .rst(f490_rst), .rdata(f490_rdata));
  assign f490_clk = clk;
  assign f490_rst = rst;
  // Bindings to f490

  // f492
  logic [0:0] f492_wen;
  logic [31:0] f492_wdata;
  logic [0:0] f492_clk;
  logic [0:0] f492_rst;
  logic [31:0] f492_rdata;
  sr_buffer_32_1 f492(.wen(f492_wen), .wdata(f492_wdata), .clk(f492_clk), .rst(f492_rst), .rdata(f492_rdata));
  assign f492_clk = clk;
  assign f492_rst = rst;
  // Bindings to f492

  // f494
  logic [0:0] f494_wen;
  logic [31:0] f494_wdata;
  logic [0:0] f494_clk;
  logic [0:0] f494_rst;
  logic [31:0] f494_rdata;
  sr_buffer_32_1 f494(.wen(f494_wen), .wdata(f494_wdata), .clk(f494_clk), .rst(f494_rst), .rdata(f494_rdata));
  assign f494_clk = clk;
  assign f494_rst = rst;
  // Bindings to f494

  // f496
  logic [0:0] f496_wen;
  logic [31:0] f496_wdata;
  logic [0:0] f496_clk;
  logic [0:0] f496_rst;
  logic [31:0] f496_rdata;
  sr_buffer_32_1 f496(.wen(f496_wen), .wdata(f496_wdata), .clk(f496_clk), .rst(f496_rst), .rdata(f496_rdata));
  assign f496_clk = clk;
  assign f496_rst = rst;
  // Bindings to f496

  // f498
  logic [0:0] f498_wen;
  logic [31:0] f498_wdata;
  logic [0:0] f498_clk;
  logic [0:0] f498_rst;
  logic [31:0] f498_rdata;
  sr_buffer_32_1 f498(.wen(f498_wen), .wdata(f498_wdata), .clk(f498_clk), .rst(f498_rst), .rdata(f498_rdata));
  assign f498_clk = clk;
  assign f498_rst = rst;
  // Bindings to f498

  // f500
  logic [0:0] f500_wen;
  logic [31:0] f500_wdata;
  logic [0:0] f500_clk;
  logic [0:0] f500_rst;
  logic [31:0] f500_rdata;
  sr_buffer_32_1 f500(.wen(f500_wen), .wdata(f500_wdata), .clk(f500_clk), .rst(f500_rst), .rdata(f500_rdata));
  assign f500_clk = clk;
  assign f500_rst = rst;
  // Bindings to f500

  // f502
  logic [0:0] f502_wen;
  logic [31:0] f502_wdata;
  logic [0:0] f502_clk;
  logic [0:0] f502_rst;
  logic [31:0] f502_rdata;
  sr_buffer_32_1 f502(.wen(f502_wen), .wdata(f502_wdata), .clk(f502_clk), .rst(f502_rst), .rdata(f502_rdata));
  assign f502_clk = clk;
  assign f502_rst = rst;
  // Bindings to f502

  // f504
  logic [0:0] f504_wen;
  logic [31:0] f504_wdata;
  logic [0:0] f504_clk;
  logic [0:0] f504_rst;
  logic [31:0] f504_rdata;
  sr_buffer_32_1 f504(.wen(f504_wen), .wdata(f504_wdata), .clk(f504_clk), .rst(f504_rst), .rdata(f504_rdata));
  assign f504_clk = clk;
  assign f504_rst = rst;
  // Bindings to f504

  // f506
  logic [0:0] f506_wen;
  logic [31:0] f506_wdata;
  logic [0:0] f506_clk;
  logic [0:0] f506_rst;
  logic [31:0] f506_rdata;
  sr_buffer_32_1 f506(.wen(f506_wen), .wdata(f506_wdata), .clk(f506_clk), .rst(f506_rst), .rdata(f506_rdata));
  assign f506_clk = clk;
  assign f506_rst = rst;
  // Bindings to f506

  // f508
  logic [0:0] f508_wen;
  logic [31:0] f508_wdata;
  logic [0:0] f508_clk;
  logic [0:0] f508_rst;
  logic [31:0] f508_rdata;
  sr_buffer_32_1 f508(.wen(f508_wen), .wdata(f508_wdata), .clk(f508_clk), .rst(f508_rst), .rdata(f508_rdata));
  assign f508_clk = clk;
  assign f508_rst = rst;
  // Bindings to f508

  // f510
  logic [0:0] f510_wen;
  logic [31:0] f510_wdata;
  logic [0:0] f510_clk;
  logic [0:0] f510_rst;
  logic [31:0] f510_rdata;
  sr_buffer_32_1 f510(.wen(f510_wen), .wdata(f510_wdata), .clk(f510_clk), .rst(f510_rst), .rdata(f510_rdata));
  assign f510_clk = clk;
  assign f510_rst = rst;
  // Bindings to f510

  // f512
  logic [0:0] f512_wen;
  logic [31:0] f512_wdata;
  logic [0:0] f512_clk;
  logic [0:0] f512_rst;
  logic [31:0] f512_rdata;
  sr_buffer_32_1 f512(.wen(f512_wen), .wdata(f512_wdata), .clk(f512_clk), .rst(f512_rst), .rdata(f512_rdata));
  assign f512_clk = clk;
  assign f512_rst = rst;
  // Bindings to f512

  // f514
  logic [0:0] f514_wen;
  logic [31:0] f514_wdata;
  logic [0:0] f514_clk;
  logic [0:0] f514_rst;
  logic [31:0] f514_rdata;
  sr_buffer_32_1 f514(.wen(f514_wen), .wdata(f514_wdata), .clk(f514_clk), .rst(f514_rst), .rdata(f514_rdata));
  assign f514_clk = clk;
  assign f514_rst = rst;
  // Bindings to f514

  // f516
  logic [0:0] f516_wen;
  logic [31:0] f516_wdata;
  logic [0:0] f516_clk;
  logic [0:0] f516_rst;
  logic [31:0] f516_rdata;
  sr_buffer_32_1 f516(.wen(f516_wen), .wdata(f516_wdata), .clk(f516_clk), .rst(f516_rst), .rdata(f516_rdata));
  assign f516_clk = clk;
  assign f516_rst = rst;
  // Bindings to f516

  // f518
  logic [0:0] f518_wen;
  logic [31:0] f518_wdata;
  logic [0:0] f518_clk;
  logic [0:0] f518_rst;
  logic [31:0] f518_rdata;
  sr_buffer_32_1 f518(.wen(f518_wen), .wdata(f518_wdata), .clk(f518_clk), .rst(f518_rst), .rdata(f518_rdata));
  assign f518_clk = clk;
  assign f518_rst = rst;
  // Bindings to f518

  // f520
  logic [0:0] f520_wen;
  logic [31:0] f520_wdata;
  logic [0:0] f520_clk;
  logic [0:0] f520_rst;
  logic [31:0] f520_rdata;
  sr_buffer_32_1 f520(.wen(f520_wen), .wdata(f520_wdata), .clk(f520_clk), .rst(f520_rst), .rdata(f520_rdata));
  assign f520_clk = clk;
  assign f520_rst = rst;
  // Bindings to f520

  // f522
  logic [0:0] f522_wen;
  logic [31:0] f522_wdata;
  logic [0:0] f522_clk;
  logic [0:0] f522_rst;
  logic [31:0] f522_rdata;
  sr_buffer_32_1 f522(.wen(f522_wen), .wdata(f522_wdata), .clk(f522_clk), .rst(f522_rst), .rdata(f522_rdata));
  assign f522_clk = clk;
  assign f522_rst = rst;
  // Bindings to f522

  // f524
  logic [0:0] f524_wen;
  logic [31:0] f524_wdata;
  logic [0:0] f524_clk;
  logic [0:0] f524_rst;
  logic [31:0] f524_rdata;
  sr_buffer_32_1 f524(.wen(f524_wen), .wdata(f524_wdata), .clk(f524_clk), .rst(f524_rst), .rdata(f524_rdata));
  assign f524_clk = clk;
  assign f524_rst = rst;
  // Bindings to f524

  // f526
  logic [0:0] f526_wen;
  logic [31:0] f526_wdata;
  logic [0:0] f526_clk;
  logic [0:0] f526_rst;
  logic [31:0] f526_rdata;
  sr_buffer_32_1 f526(.wen(f526_wen), .wdata(f526_wdata), .clk(f526_clk), .rst(f526_rst), .rdata(f526_rdata));
  assign f526_clk = clk;
  assign f526_rst = rst;
  // Bindings to f526

  // f528
  logic [0:0] f528_wen;
  logic [31:0] f528_wdata;
  logic [0:0] f528_clk;
  logic [0:0] f528_rst;
  logic [31:0] f528_rdata;
  sr_buffer_32_1 f528(.wen(f528_wen), .wdata(f528_wdata), .clk(f528_clk), .rst(f528_rst), .rdata(f528_rdata));
  assign f528_clk = clk;
  assign f528_rst = rst;
  // Bindings to f528

  // f530
  logic [0:0] f530_wen;
  logic [31:0] f530_wdata;
  logic [0:0] f530_clk;
  logic [0:0] f530_rst;
  logic [31:0] f530_rdata;
  sr_buffer_32_1 f530(.wen(f530_wen), .wdata(f530_wdata), .clk(f530_clk), .rst(f530_rst), .rdata(f530_rdata));
  assign f530_clk = clk;
  assign f530_rst = rst;
  // Bindings to f530

  // f532
  logic [0:0] f532_wen;
  logic [31:0] f532_wdata;
  logic [0:0] f532_clk;
  logic [0:0] f532_rst;
  logic [31:0] f532_rdata;
  sr_buffer_32_1 f532(.wen(f532_wen), .wdata(f532_wdata), .clk(f532_clk), .rst(f532_rst), .rdata(f532_rdata));
  assign f532_clk = clk;
  assign f532_rst = rst;
  // Bindings to f532

  // f534
  logic [0:0] f534_wen;
  logic [31:0] f534_wdata;
  logic [0:0] f534_clk;
  logic [0:0] f534_rst;
  logic [31:0] f534_rdata;
  sr_buffer_32_1 f534(.wen(f534_wen), .wdata(f534_wdata), .clk(f534_clk), .rst(f534_rst), .rdata(f534_rdata));
  assign f534_clk = clk;
  assign f534_rst = rst;
  // Bindings to f534

  // f536
  logic [0:0] f536_wen;
  logic [31:0] f536_wdata;
  logic [0:0] f536_clk;
  logic [0:0] f536_rst;
  logic [31:0] f536_rdata;
  sr_buffer_32_1 f536(.wen(f536_wen), .wdata(f536_wdata), .clk(f536_clk), .rst(f536_rst), .rdata(f536_rdata));
  assign f536_clk = clk;
  assign f536_rst = rst;
  // Bindings to f536

  // f538
  logic [0:0] f538_wen;
  logic [31:0] f538_wdata;
  logic [0:0] f538_clk;
  logic [0:0] f538_rst;
  logic [31:0] f538_rdata;
  sr_buffer_32_1 f538(.wen(f538_wen), .wdata(f538_wdata), .clk(f538_clk), .rst(f538_rst), .rdata(f538_rdata));
  assign f538_clk = clk;
  assign f538_rst = rst;
  // Bindings to f538

  // f540
  logic [0:0] f540_wen;
  logic [31:0] f540_wdata;
  logic [0:0] f540_clk;
  logic [0:0] f540_rst;
  logic [31:0] f540_rdata;
  sr_buffer_32_1 f540(.wen(f540_wen), .wdata(f540_wdata), .clk(f540_clk), .rst(f540_rst), .rdata(f540_rdata));
  assign f540_clk = clk;
  assign f540_rst = rst;
  // Bindings to f540

  // f542
  logic [0:0] f542_wen;
  logic [31:0] f542_wdata;
  logic [0:0] f542_clk;
  logic [0:0] f542_rst;
  logic [31:0] f542_rdata;
  sr_buffer_32_1 f542(.wen(f542_wen), .wdata(f542_wdata), .clk(f542_clk), .rst(f542_rst), .rdata(f542_rdata));
  assign f542_clk = clk;
  assign f542_rst = rst;
  // Bindings to f542

  // f544
  logic [0:0] f544_wen;
  logic [31:0] f544_wdata;
  logic [0:0] f544_clk;
  logic [0:0] f544_rst;
  logic [31:0] f544_rdata;
  sr_buffer_32_1 f544(.wen(f544_wen), .wdata(f544_wdata), .clk(f544_clk), .rst(f544_rst), .rdata(f544_rdata));
  assign f544_clk = clk;
  assign f544_rst = rst;
  // Bindings to f544

  // f546
  logic [0:0] f546_wen;
  logic [31:0] f546_wdata;
  logic [0:0] f546_clk;
  logic [0:0] f546_rst;
  logic [31:0] f546_rdata;
  sr_buffer_32_1 f546(.wen(f546_wen), .wdata(f546_wdata), .clk(f546_clk), .rst(f546_rst), .rdata(f546_rdata));
  assign f546_clk = clk;
  assign f546_rst = rst;
  // Bindings to f546

  // f548
  logic [0:0] f548_wen;
  logic [31:0] f548_wdata;
  logic [0:0] f548_clk;
  logic [0:0] f548_rst;
  logic [31:0] f548_rdata;
  sr_buffer_32_1 f548(.wen(f548_wen), .wdata(f548_wdata), .clk(f548_clk), .rst(f548_rst), .rdata(f548_rdata));
  assign f548_clk = clk;
  assign f548_rst = rst;
  // Bindings to f548

  // f550
  logic [0:0] f550_wen;
  logic [31:0] f550_wdata;
  logic [0:0] f550_clk;
  logic [0:0] f550_rst;
  logic [31:0] f550_rdata;
  sr_buffer_32_1 f550(.wen(f550_wen), .wdata(f550_wdata), .clk(f550_clk), .rst(f550_rst), .rdata(f550_rdata));
  assign f550_clk = clk;
  assign f550_rst = rst;
  // Bindings to f550

  // f552
  logic [0:0] f552_wen;
  logic [31:0] f552_wdata;
  logic [0:0] f552_clk;
  logic [0:0] f552_rst;
  logic [31:0] f552_rdata;
  sr_buffer_32_1 f552(.wen(f552_wen), .wdata(f552_wdata), .clk(f552_clk), .rst(f552_rst), .rdata(f552_rdata));
  assign f552_clk = clk;
  assign f552_rst = rst;
  // Bindings to f552

  // f554
  logic [0:0] f554_wen;
  logic [31:0] f554_wdata;
  logic [0:0] f554_clk;
  logic [0:0] f554_rst;
  logic [31:0] f554_rdata;
  sr_buffer_32_1 f554(.wen(f554_wen), .wdata(f554_wdata), .clk(f554_clk), .rst(f554_rst), .rdata(f554_rdata));
  assign f554_clk = clk;
  assign f554_rst = rst;
  // Bindings to f554

  // f556
  logic [0:0] f556_wen;
  logic [31:0] f556_wdata;
  logic [0:0] f556_clk;
  logic [0:0] f556_rst;
  logic [31:0] f556_rdata;
  sr_buffer_32_1 f556(.wen(f556_wen), .wdata(f556_wdata), .clk(f556_clk), .rst(f556_rst), .rdata(f556_rdata));
  assign f556_clk = clk;
  assign f556_rst = rst;
  // Bindings to f556

  // f558
  logic [0:0] f558_wen;
  logic [31:0] f558_wdata;
  logic [0:0] f558_clk;
  logic [0:0] f558_rst;
  logic [31:0] f558_rdata;
  sr_buffer_32_1 f558(.wen(f558_wen), .wdata(f558_wdata), .clk(f558_clk), .rst(f558_rst), .rdata(f558_rdata));
  assign f558_clk = clk;
  assign f558_rst = rst;
  // Bindings to f558

  // f560
  logic [0:0] f560_wen;
  logic [31:0] f560_wdata;
  logic [0:0] f560_clk;
  logic [0:0] f560_rst;
  logic [31:0] f560_rdata;
  sr_buffer_32_1 f560(.wen(f560_wen), .wdata(f560_wdata), .clk(f560_clk), .rst(f560_rst), .rdata(f560_rdata));
  assign f560_clk = clk;
  assign f560_rst = rst;
  // Bindings to f560

  // f562
  logic [0:0] f562_wen;
  logic [31:0] f562_wdata;
  logic [0:0] f562_clk;
  logic [0:0] f562_rst;
  logic [31:0] f562_rdata;
  sr_buffer_32_1 f562(.wen(f562_wen), .wdata(f562_wdata), .clk(f562_clk), .rst(f562_rst), .rdata(f562_rdata));
  assign f562_clk = clk;
  assign f562_rst = rst;
  // Bindings to f562

  // f564
  logic [0:0] f564_wen;
  logic [31:0] f564_wdata;
  logic [0:0] f564_clk;
  logic [0:0] f564_rst;
  logic [31:0] f564_rdata;
  sr_buffer_32_1 f564(.wen(f564_wen), .wdata(f564_wdata), .clk(f564_clk), .rst(f564_rst), .rdata(f564_rdata));
  assign f564_clk = clk;
  assign f564_rst = rst;
  // Bindings to f564

  // f566
  logic [0:0] f566_wen;
  logic [31:0] f566_wdata;
  logic [0:0] f566_clk;
  logic [0:0] f566_rst;
  logic [31:0] f566_rdata;
  sr_buffer_32_1 f566(.wen(f566_wen), .wdata(f566_wdata), .clk(f566_clk), .rst(f566_rst), .rdata(f566_rdata));
  assign f566_clk = clk;
  assign f566_rst = rst;
  // Bindings to f566

  // f568
  logic [0:0] f568_wen;
  logic [31:0] f568_wdata;
  logic [0:0] f568_clk;
  logic [0:0] f568_rst;
  logic [31:0] f568_rdata;
  sr_buffer_32_1 f568(.wen(f568_wen), .wdata(f568_wdata), .clk(f568_clk), .rst(f568_rst), .rdata(f568_rdata));
  assign f568_clk = clk;
  assign f568_rst = rst;
  // Bindings to f568

  // f570
  logic [0:0] f570_wen;
  logic [31:0] f570_wdata;
  logic [0:0] f570_clk;
  logic [0:0] f570_rst;
  logic [31:0] f570_rdata;
  sr_buffer_32_1 f570(.wen(f570_wen), .wdata(f570_wdata), .clk(f570_clk), .rst(f570_rst), .rdata(f570_rdata));
  assign f570_clk = clk;
  assign f570_rst = rst;
  // Bindings to f570

  // f572
  logic [0:0] f572_wen;
  logic [31:0] f572_wdata;
  logic [0:0] f572_clk;
  logic [0:0] f572_rst;
  logic [31:0] f572_rdata;
  sr_buffer_32_1 f572(.wen(f572_wen), .wdata(f572_wdata), .clk(f572_clk), .rst(f572_rst), .rdata(f572_rdata));
  assign f572_clk = clk;
  assign f572_rst = rst;
  // Bindings to f572

  // f574
  logic [0:0] f574_wen;
  logic [31:0] f574_wdata;
  logic [0:0] f574_clk;
  logic [0:0] f574_rst;
  logic [31:0] f574_rdata;
  sr_buffer_32_1 f574(.wen(f574_wen), .wdata(f574_wdata), .clk(f574_clk), .rst(f574_rst), .rdata(f574_rdata));
  assign f574_clk = clk;
  assign f574_rst = rst;
  // Bindings to f574

  // f576
  logic [0:0] f576_wen;
  logic [31:0] f576_wdata;
  logic [0:0] f576_clk;
  logic [0:0] f576_rst;
  logic [31:0] f576_rdata;
  sr_buffer_32_1 f576(.wen(f576_wen), .wdata(f576_wdata), .clk(f576_clk), .rst(f576_rst), .rdata(f576_rdata));
  assign f576_clk = clk;
  assign f576_rst = rst;
  // Bindings to f576

  // f578
  logic [0:0] f578_wen;
  logic [31:0] f578_wdata;
  logic [0:0] f578_clk;
  logic [0:0] f578_rst;
  logic [31:0] f578_rdata;
  sr_buffer_32_1 f578(.wen(f578_wen), .wdata(f578_wdata), .clk(f578_clk), .rst(f578_rst), .rdata(f578_rdata));
  assign f578_clk = clk;
  assign f578_rst = rst;
  // Bindings to f578

  // f580
  logic [0:0] f580_wen;
  logic [31:0] f580_wdata;
  logic [0:0] f580_clk;
  logic [0:0] f580_rst;
  logic [31:0] f580_rdata;
  sr_buffer_32_1 f580(.wen(f580_wen), .wdata(f580_wdata), .clk(f580_clk), .rst(f580_rst), .rdata(f580_rdata));
  assign f580_clk = clk;
  assign f580_rst = rst;
  // Bindings to f580

  // f582
  logic [0:0] f582_wen;
  logic [31:0] f582_wdata;
  logic [0:0] f582_clk;
  logic [0:0] f582_rst;
  logic [31:0] f582_rdata;
  sr_buffer_32_1 f582(.wen(f582_wen), .wdata(f582_wdata), .clk(f582_clk), .rst(f582_rst), .rdata(f582_rdata));
  assign f582_clk = clk;
  assign f582_rst = rst;
  // Bindings to f582

  // f584
  logic [0:0] f584_wen;
  logic [31:0] f584_wdata;
  logic [0:0] f584_clk;
  logic [0:0] f584_rst;
  logic [31:0] f584_rdata;
  sr_buffer_32_1 f584(.wen(f584_wen), .wdata(f584_wdata), .clk(f584_clk), .rst(f584_rst), .rdata(f584_rdata));
  assign f584_clk = clk;
  assign f584_rst = rst;
  // Bindings to f584

  // f586
  logic [0:0] f586_wen;
  logic [31:0] f586_wdata;
  logic [0:0] f586_clk;
  logic [0:0] f586_rst;
  logic [31:0] f586_rdata;
  sr_buffer_32_1 f586(.wen(f586_wen), .wdata(f586_wdata), .clk(f586_clk), .rst(f586_rst), .rdata(f586_rdata));
  assign f586_clk = clk;
  assign f586_rst = rst;
  // Bindings to f586

  // f588
  logic [0:0] f588_wen;
  logic [31:0] f588_wdata;
  logic [0:0] f588_clk;
  logic [0:0] f588_rst;
  logic [31:0] f588_rdata;
  sr_buffer_32_1 f588(.wen(f588_wen), .wdata(f588_wdata), .clk(f588_clk), .rst(f588_rst), .rdata(f588_rdata));
  assign f588_clk = clk;
  assign f588_rst = rst;
  // Bindings to f588

  // f590
  logic [0:0] f590_wen;
  logic [31:0] f590_wdata;
  logic [0:0] f590_clk;
  logic [0:0] f590_rst;
  logic [31:0] f590_rdata;
  sr_buffer_32_1 f590(.wen(f590_wen), .wdata(f590_wdata), .clk(f590_clk), .rst(f590_rst), .rdata(f590_rdata));
  assign f590_clk = clk;
  assign f590_rst = rst;
  // Bindings to f590

  // f592
  logic [0:0] f592_wen;
  logic [31:0] f592_wdata;
  logic [0:0] f592_clk;
  logic [0:0] f592_rst;
  logic [31:0] f592_rdata;
  sr_buffer_32_1 f592(.wen(f592_wen), .wdata(f592_wdata), .clk(f592_clk), .rst(f592_rst), .rdata(f592_rdata));
  assign f592_clk = clk;
  assign f592_rst = rst;
  // Bindings to f592

  // f594
  logic [0:0] f594_wen;
  logic [31:0] f594_wdata;
  logic [0:0] f594_clk;
  logic [0:0] f594_rst;
  logic [31:0] f594_rdata;
  sr_buffer_32_1 f594(.wen(f594_wen), .wdata(f594_wdata), .clk(f594_clk), .rst(f594_rst), .rdata(f594_rdata));
  assign f594_clk = clk;
  assign f594_rst = rst;
  // Bindings to f594

  // f596
  logic [0:0] f596_wen;
  logic [31:0] f596_wdata;
  logic [0:0] f596_clk;
  logic [0:0] f596_rst;
  logic [31:0] f596_rdata;
  sr_buffer_32_1 f596(.wen(f596_wen), .wdata(f596_wdata), .clk(f596_clk), .rst(f596_rst), .rdata(f596_rdata));
  assign f596_clk = clk;
  assign f596_rst = rst;
  // Bindings to f596

  // f598
  logic [0:0] f598_wen;
  logic [31:0] f598_wdata;
  logic [0:0] f598_clk;
  logic [0:0] f598_rst;
  logic [31:0] f598_rdata;
  sr_buffer_32_1 f598(.wen(f598_wen), .wdata(f598_wdata), .clk(f598_clk), .rst(f598_rst), .rdata(f598_rdata));
  assign f598_clk = clk;
  assign f598_rst = rst;
  // Bindings to f598

  // f600
  logic [0:0] f600_wen;
  logic [31:0] f600_wdata;
  logic [0:0] f600_clk;
  logic [0:0] f600_rst;
  logic [31:0] f600_rdata;
  sr_buffer_32_1 f600(.wen(f600_wen), .wdata(f600_wdata), .clk(f600_clk), .rst(f600_rst), .rdata(f600_rdata));
  assign f600_clk = clk;
  assign f600_rst = rst;
  // Bindings to f600

  // f602
  logic [0:0] f602_wen;
  logic [31:0] f602_wdata;
  logic [0:0] f602_clk;
  logic [0:0] f602_rst;
  logic [31:0] f602_rdata;
  sr_buffer_32_1 f602(.wen(f602_wen), .wdata(f602_wdata), .clk(f602_clk), .rst(f602_rst), .rdata(f602_rdata));
  assign f602_clk = clk;
  assign f602_rst = rst;
  // Bindings to f602

  // f604
  logic [0:0] f604_wen;
  logic [31:0] f604_wdata;
  logic [0:0] f604_clk;
  logic [0:0] f604_rst;
  logic [31:0] f604_rdata;
  sr_buffer_32_1 f604(.wen(f604_wen), .wdata(f604_wdata), .clk(f604_clk), .rst(f604_rst), .rdata(f604_rdata));
  assign f604_clk = clk;
  assign f604_rst = rst;
  // Bindings to f604

  // f606
  logic [0:0] f606_wen;
  logic [31:0] f606_wdata;
  logic [0:0] f606_clk;
  logic [0:0] f606_rst;
  logic [31:0] f606_rdata;
  sr_buffer_32_1 f606(.wen(f606_wen), .wdata(f606_wdata), .clk(f606_clk), .rst(f606_rst), .rdata(f606_rdata));
  assign f606_clk = clk;
  assign f606_rst = rst;
  // Bindings to f606

  // f608
  logic [0:0] f608_wen;
  logic [31:0] f608_wdata;
  logic [0:0] f608_clk;
  logic [0:0] f608_rst;
  logic [31:0] f608_rdata;
  sr_buffer_32_1 f608(.wen(f608_wen), .wdata(f608_wdata), .clk(f608_clk), .rst(f608_rst), .rdata(f608_rdata));
  assign f608_clk = clk;
  assign f608_rst = rst;
  // Bindings to f608

  // f610
  logic [0:0] f610_wen;
  logic [31:0] f610_wdata;
  logic [0:0] f610_clk;
  logic [0:0] f610_rst;
  logic [31:0] f610_rdata;
  sr_buffer_32_1 f610(.wen(f610_wen), .wdata(f610_wdata), .clk(f610_clk), .rst(f610_rst), .rdata(f610_rdata));
  assign f610_clk = clk;
  assign f610_rst = rst;
  // Bindings to f610

  // f612
  logic [0:0] f612_wen;
  logic [31:0] f612_wdata;
  logic [0:0] f612_clk;
  logic [0:0] f612_rst;
  logic [31:0] f612_rdata;
  sr_buffer_32_1 f612(.wen(f612_wen), .wdata(f612_wdata), .clk(f612_clk), .rst(f612_rst), .rdata(f612_rdata));
  assign f612_clk = clk;
  assign f612_rst = rst;
  // Bindings to f612

  // f614
  logic [0:0] f614_wen;
  logic [31:0] f614_wdata;
  logic [0:0] f614_clk;
  logic [0:0] f614_rst;
  logic [31:0] f614_rdata;
  sr_buffer_32_1 f614(.wen(f614_wen), .wdata(f614_wdata), .clk(f614_clk), .rst(f614_rst), .rdata(f614_rdata));
  assign f614_clk = clk;
  assign f614_rst = rst;
  // Bindings to f614

  // f616
  logic [0:0] f616_wen;
  logic [31:0] f616_wdata;
  logic [0:0] f616_clk;
  logic [0:0] f616_rst;
  logic [31:0] f616_rdata;
  sr_buffer_32_1 f616(.wen(f616_wen), .wdata(f616_wdata), .clk(f616_clk), .rst(f616_rst), .rdata(f616_rdata));
  assign f616_clk = clk;
  assign f616_rst = rst;
  // Bindings to f616

  // f618
  logic [0:0] f618_wen;
  logic [31:0] f618_wdata;
  logic [0:0] f618_clk;
  logic [0:0] f618_rst;
  logic [31:0] f618_rdata;
  sr_buffer_32_1 f618(.wen(f618_wen), .wdata(f618_wdata), .clk(f618_clk), .rst(f618_rst), .rdata(f618_rdata));
  assign f618_clk = clk;
  assign f618_rst = rst;
  // Bindings to f618

  // f620
  logic [0:0] f620_wen;
  logic [31:0] f620_wdata;
  logic [0:0] f620_clk;
  logic [0:0] f620_rst;
  logic [31:0] f620_rdata;
  sr_buffer_32_1 f620(.wen(f620_wen), .wdata(f620_wdata), .clk(f620_clk), .rst(f620_rst), .rdata(f620_rdata));
  assign f620_clk = clk;
  assign f620_rst = rst;
  // Bindings to f620

  // f622
  logic [0:0] f622_wen;
  logic [31:0] f622_wdata;
  logic [0:0] f622_clk;
  logic [0:0] f622_rst;
  logic [31:0] f622_rdata;
  sr_buffer_32_1 f622(.wen(f622_wen), .wdata(f622_wdata), .clk(f622_clk), .rst(f622_rst), .rdata(f622_rdata));
  assign f622_clk = clk;
  assign f622_rst = rst;
  // Bindings to f622

  // f624
  logic [0:0] f624_wen;
  logic [31:0] f624_wdata;
  logic [0:0] f624_clk;
  logic [0:0] f624_rst;
  logic [31:0] f624_rdata;
  sr_buffer_32_1 f624(.wen(f624_wen), .wdata(f624_wdata), .clk(f624_clk), .rst(f624_rst), .rdata(f624_rdata));
  assign f624_clk = clk;
  assign f624_rst = rst;
  // Bindings to f624

  // f626
  logic [0:0] f626_wen;
  logic [31:0] f626_wdata;
  logic [0:0] f626_clk;
  logic [0:0] f626_rst;
  logic [31:0] f626_rdata;
  sr_buffer_32_1 f626(.wen(f626_wen), .wdata(f626_wdata), .clk(f626_clk), .rst(f626_rst), .rdata(f626_rdata));
  assign f626_clk = clk;
  assign f626_rst = rst;
  // Bindings to f626

  // f628
  logic [0:0] f628_wen;
  logic [31:0] f628_wdata;
  logic [0:0] f628_clk;
  logic [0:0] f628_rst;
  logic [31:0] f628_rdata;
  sr_buffer_32_1 f628(.wen(f628_wen), .wdata(f628_wdata), .clk(f628_clk), .rst(f628_rst), .rdata(f628_rdata));
  assign f628_clk = clk;
  assign f628_rst = rst;
  // Bindings to f628

  // f630
  logic [0:0] f630_wen;
  logic [31:0] f630_wdata;
  logic [0:0] f630_clk;
  logic [0:0] f630_rst;
  logic [31:0] f630_rdata;
  sr_buffer_32_1 f630(.wen(f630_wen), .wdata(f630_wdata), .clk(f630_clk), .rst(f630_rst), .rdata(f630_rdata));
  assign f630_clk = clk;
  assign f630_rst = rst;
  // Bindings to f630

  // f632
  logic [0:0] f632_wen;
  logic [31:0] f632_wdata;
  logic [0:0] f632_clk;
  logic [0:0] f632_rst;
  logic [31:0] f632_rdata;
  sr_buffer_32_1 f632(.wen(f632_wen), .wdata(f632_wdata), .clk(f632_clk), .rst(f632_rst), .rdata(f632_rdata));
  assign f632_clk = clk;
  assign f632_rst = rst;
  // Bindings to f632

  // f634
  logic [0:0] f634_wen;
  logic [31:0] f634_wdata;
  logic [0:0] f634_clk;
  logic [0:0] f634_rst;
  logic [31:0] f634_rdata;
  sr_buffer_32_1 f634(.wen(f634_wen), .wdata(f634_wdata), .clk(f634_clk), .rst(f634_rst), .rdata(f634_rdata));
  assign f634_clk = clk;
  assign f634_rst = rst;
  // Bindings to f634

  // f636
  logic [0:0] f636_wen;
  logic [31:0] f636_wdata;
  logic [0:0] f636_clk;
  logic [0:0] f636_rst;
  logic [31:0] f636_rdata;
  sr_buffer_32_1 f636(.wen(f636_wen), .wdata(f636_wdata), .clk(f636_clk), .rst(f636_rst), .rdata(f636_rdata));
  assign f636_clk = clk;
  assign f636_rst = rst;
  // Bindings to f636

  // f638
  logic [0:0] f638_wen;
  logic [31:0] f638_wdata;
  logic [0:0] f638_clk;
  logic [0:0] f638_rst;
  logic [31:0] f638_rdata;
  sr_buffer_32_1 f638(.wen(f638_wen), .wdata(f638_wdata), .clk(f638_clk), .rst(f638_rst), .rdata(f638_rdata));
  assign f638_clk = clk;
  assign f638_rst = rst;
  // Bindings to f638

  // f640
  logic [0:0] f640_wen;
  logic [31:0] f640_wdata;
  logic [0:0] f640_clk;
  logic [0:0] f640_rst;
  logic [31:0] f640_rdata;
  sr_buffer_32_1 f640(.wen(f640_wen), .wdata(f640_wdata), .clk(f640_clk), .rst(f640_rst), .rdata(f640_rdata));
  assign f640_clk = clk;
  assign f640_rst = rst;
  // Bindings to f640

  // f642
  logic [0:0] f642_wen;
  logic [31:0] f642_wdata;
  logic [0:0] f642_clk;
  logic [0:0] f642_rst;
  logic [31:0] f642_rdata;
  sr_buffer_32_1 f642(.wen(f642_wen), .wdata(f642_wdata), .clk(f642_clk), .rst(f642_rst), .rdata(f642_rdata));
  assign f642_clk = clk;
  assign f642_rst = rst;
  // Bindings to f642

  // f644
  logic [0:0] f644_wen;
  logic [31:0] f644_wdata;
  logic [0:0] f644_clk;
  logic [0:0] f644_rst;
  logic [31:0] f644_rdata;
  sr_buffer_32_1 f644(.wen(f644_wen), .wdata(f644_wdata), .clk(f644_clk), .rst(f644_rst), .rdata(f644_rdata));
  assign f644_clk = clk;
  assign f644_rst = rst;
  // Bindings to f644

  // f646
  logic [0:0] f646_wen;
  logic [31:0] f646_wdata;
  logic [0:0] f646_clk;
  logic [0:0] f646_rst;
  logic [31:0] f646_rdata;
  sr_buffer_32_1 f646(.wen(f646_wen), .wdata(f646_wdata), .clk(f646_clk), .rst(f646_rst), .rdata(f646_rdata));
  assign f646_clk = clk;
  assign f646_rst = rst;
  // Bindings to f646

  // f648
  logic [0:0] f648_wen;
  logic [31:0] f648_wdata;
  logic [0:0] f648_clk;
  logic [0:0] f648_rst;
  logic [31:0] f648_rdata;
  sr_buffer_32_1 f648(.wen(f648_wen), .wdata(f648_wdata), .clk(f648_clk), .rst(f648_rst), .rdata(f648_rdata));
  assign f648_clk = clk;
  assign f648_rst = rst;
  // Bindings to f648

  // f650
  logic [0:0] f650_wen;
  logic [31:0] f650_wdata;
  logic [0:0] f650_clk;
  logic [0:0] f650_rst;
  logic [31:0] f650_rdata;
  sr_buffer_32_1 f650(.wen(f650_wen), .wdata(f650_wdata), .clk(f650_clk), .rst(f650_rst), .rdata(f650_rdata));
  assign f650_clk = clk;
  assign f650_rst = rst;
  // Bindings to f650

  // f652
  logic [0:0] f652_wen;
  logic [31:0] f652_wdata;
  logic [0:0] f652_clk;
  logic [0:0] f652_rst;
  logic [31:0] f652_rdata;
  sr_buffer_32_1 f652(.wen(f652_wen), .wdata(f652_wdata), .clk(f652_clk), .rst(f652_rst), .rdata(f652_rdata));
  assign f652_clk = clk;
  assign f652_rst = rst;
  // Bindings to f652

  // f654
  logic [0:0] f654_wen;
  logic [31:0] f654_wdata;
  logic [0:0] f654_clk;
  logic [0:0] f654_rst;
  logic [31:0] f654_rdata;
  sr_buffer_32_1 f654(.wen(f654_wen), .wdata(f654_wdata), .clk(f654_clk), .rst(f654_rst), .rdata(f654_rdata));
  assign f654_clk = clk;
  assign f654_rst = rst;
  // Bindings to f654

  // f656
  logic [0:0] f656_wen;
  logic [31:0] f656_wdata;
  logic [0:0] f656_clk;
  logic [0:0] f656_rst;
  logic [31:0] f656_rdata;
  sr_buffer_32_1 f656(.wen(f656_wen), .wdata(f656_wdata), .clk(f656_clk), .rst(f656_rst), .rdata(f656_rdata));
  assign f656_clk = clk;
  assign f656_rst = rst;
  // Bindings to f656

  // f658
  logic [0:0] f658_wen;
  logic [31:0] f658_wdata;
  logic [0:0] f658_clk;
  logic [0:0] f658_rst;
  logic [31:0] f658_rdata;
  sr_buffer_32_1 f658(.wen(f658_wen), .wdata(f658_wdata), .clk(f658_clk), .rst(f658_rst), .rdata(f658_rdata));
  assign f658_clk = clk;
  assign f658_rst = rst;
  // Bindings to f658

  // f660
  logic [0:0] f660_wen;
  logic [31:0] f660_wdata;
  logic [0:0] f660_clk;
  logic [0:0] f660_rst;
  logic [31:0] f660_rdata;
  sr_buffer_32_1 f660(.wen(f660_wen), .wdata(f660_wdata), .clk(f660_clk), .rst(f660_rst), .rdata(f660_rdata));
  assign f660_clk = clk;
  assign f660_rst = rst;
  // Bindings to f660

  // f662
  logic [0:0] f662_wen;
  logic [31:0] f662_wdata;
  logic [0:0] f662_clk;
  logic [0:0] f662_rst;
  logic [31:0] f662_rdata;
  sr_buffer_32_1 f662(.wen(f662_wen), .wdata(f662_wdata), .clk(f662_clk), .rst(f662_rst), .rdata(f662_rdata));
  assign f662_clk = clk;
  assign f662_rst = rst;
  // Bindings to f662

  // f664
  logic [0:0] f664_wen;
  logic [31:0] f664_wdata;
  logic [0:0] f664_clk;
  logic [0:0] f664_rst;
  logic [31:0] f664_rdata;
  sr_buffer_32_1 f664(.wen(f664_wen), .wdata(f664_wdata), .clk(f664_clk), .rst(f664_rst), .rdata(f664_rdata));
  assign f664_clk = clk;
  assign f664_rst = rst;
  // Bindings to f664

  // f666
  logic [0:0] f666_wen;
  logic [31:0] f666_wdata;
  logic [0:0] f666_clk;
  logic [0:0] f666_rst;
  logic [31:0] f666_rdata;
  sr_buffer_32_1 f666(.wen(f666_wen), .wdata(f666_wdata), .clk(f666_clk), .rst(f666_rst), .rdata(f666_rdata));
  assign f666_clk = clk;
  assign f666_rst = rst;
  // Bindings to f666

  // f668
  logic [0:0] f668_wen;
  logic [31:0] f668_wdata;
  logic [0:0] f668_clk;
  logic [0:0] f668_rst;
  logic [31:0] f668_rdata;
  sr_buffer_32_1 f668(.wen(f668_wen), .wdata(f668_wdata), .clk(f668_clk), .rst(f668_rst), .rdata(f668_rdata));
  assign f668_clk = clk;
  assign f668_rst = rst;
  // Bindings to f668

  // f670
  logic [0:0] f670_wen;
  logic [31:0] f670_wdata;
  logic [0:0] f670_clk;
  logic [0:0] f670_rst;
  logic [31:0] f670_rdata;
  sr_buffer_32_1 f670(.wen(f670_wen), .wdata(f670_wdata), .clk(f670_clk), .rst(f670_rst), .rdata(f670_rdata));
  assign f670_clk = clk;
  assign f670_rst = rst;
  // Bindings to f670

  // f672
  logic [0:0] f672_wen;
  logic [31:0] f672_wdata;
  logic [0:0] f672_clk;
  logic [0:0] f672_rst;
  logic [31:0] f672_rdata;
  sr_buffer_32_1 f672(.wen(f672_wen), .wdata(f672_wdata), .clk(f672_clk), .rst(f672_rst), .rdata(f672_rdata));
  assign f672_clk = clk;
  assign f672_rst = rst;
  // Bindings to f672

  // f674
  logic [0:0] f674_wen;
  logic [31:0] f674_wdata;
  logic [0:0] f674_clk;
  logic [0:0] f674_rst;
  logic [31:0] f674_rdata;
  sr_buffer_32_1 f674(.wen(f674_wen), .wdata(f674_wdata), .clk(f674_clk), .rst(f674_rst), .rdata(f674_rdata));
  assign f674_clk = clk;
  assign f674_rst = rst;
  // Bindings to f674

  // f676
  logic [0:0] f676_wen;
  logic [31:0] f676_wdata;
  logic [0:0] f676_clk;
  logic [0:0] f676_rst;
  logic [31:0] f676_rdata;
  sr_buffer_32_1 f676(.wen(f676_wen), .wdata(f676_wdata), .clk(f676_clk), .rst(f676_rst), .rdata(f676_rdata));
  assign f676_clk = clk;
  assign f676_rst = rst;
  // Bindings to f676

  // f678
  logic [0:0] f678_wen;
  logic [31:0] f678_wdata;
  logic [0:0] f678_clk;
  logic [0:0] f678_rst;
  logic [31:0] f678_rdata;
  sr_buffer_32_1 f678(.wen(f678_wen), .wdata(f678_wdata), .clk(f678_clk), .rst(f678_rst), .rdata(f678_rdata));
  assign f678_clk = clk;
  assign f678_rst = rst;
  // Bindings to f678

  // f680
  logic [0:0] f680_wen;
  logic [31:0] f680_wdata;
  logic [0:0] f680_clk;
  logic [0:0] f680_rst;
  logic [31:0] f680_rdata;
  sr_buffer_32_1 f680(.wen(f680_wen), .wdata(f680_wdata), .clk(f680_clk), .rst(f680_rst), .rdata(f680_rdata));
  assign f680_clk = clk;
  assign f680_rst = rst;
  // Bindings to f680

  // f682
  logic [0:0] f682_wen;
  logic [31:0] f682_wdata;
  logic [0:0] f682_clk;
  logic [0:0] f682_rst;
  logic [31:0] f682_rdata;
  sr_buffer_32_1 f682(.wen(f682_wen), .wdata(f682_wdata), .clk(f682_clk), .rst(f682_rst), .rdata(f682_rdata));
  assign f682_clk = clk;
  assign f682_rst = rst;
  // Bindings to f682

  // f684
  logic [0:0] f684_wen;
  logic [31:0] f684_wdata;
  logic [0:0] f684_clk;
  logic [0:0] f684_rst;
  logic [31:0] f684_rdata;
  sr_buffer_32_1 f684(.wen(f684_wen), .wdata(f684_wdata), .clk(f684_clk), .rst(f684_rst), .rdata(f684_rdata));
  assign f684_clk = clk;
  assign f684_rst = rst;
  // Bindings to f684

  // f686
  logic [0:0] f686_wen;
  logic [31:0] f686_wdata;
  logic [0:0] f686_clk;
  logic [0:0] f686_rst;
  logic [31:0] f686_rdata;
  sr_buffer_32_1 f686(.wen(f686_wen), .wdata(f686_wdata), .clk(f686_clk), .rst(f686_rst), .rdata(f686_rdata));
  assign f686_clk = clk;
  assign f686_rst = rst;
  // Bindings to f686

  // f688
  logic [0:0] f688_wen;
  logic [31:0] f688_wdata;
  logic [0:0] f688_clk;
  logic [0:0] f688_rst;
  logic [31:0] f688_rdata;
  sr_buffer_32_1 f688(.wen(f688_wen), .wdata(f688_wdata), .clk(f688_clk), .rst(f688_rst), .rdata(f688_rdata));
  assign f688_clk = clk;
  assign f688_rst = rst;
  // Bindings to f688

  // f690
  logic [0:0] f690_wen;
  logic [31:0] f690_wdata;
  logic [0:0] f690_clk;
  logic [0:0] f690_rst;
  logic [31:0] f690_rdata;
  sr_buffer_32_1 f690(.wen(f690_wen), .wdata(f690_wdata), .clk(f690_clk), .rst(f690_rst), .rdata(f690_rdata));
  assign f690_clk = clk;
  assign f690_rst = rst;
  // Bindings to f690

  // f692
  logic [0:0] f692_wen;
  logic [31:0] f692_wdata;
  logic [0:0] f692_clk;
  logic [0:0] f692_rst;
  logic [31:0] f692_rdata;
  sr_buffer_32_1 f692(.wen(f692_wen), .wdata(f692_wdata), .clk(f692_clk), .rst(f692_rst), .rdata(f692_rdata));
  assign f692_clk = clk;
  assign f692_rst = rst;
  // Bindings to f692

  // f694
  logic [0:0] f694_wen;
  logic [31:0] f694_wdata;
  logic [0:0] f694_clk;
  logic [0:0] f694_rst;
  logic [31:0] f694_rdata;
  sr_buffer_32_1 f694(.wen(f694_wen), .wdata(f694_wdata), .clk(f694_clk), .rst(f694_rst), .rdata(f694_rdata));
  assign f694_clk = clk;
  assign f694_rst = rst;
  // Bindings to f694

  // f696
  logic [0:0] f696_wen;
  logic [31:0] f696_wdata;
  logic [0:0] f696_clk;
  logic [0:0] f696_rst;
  logic [31:0] f696_rdata;
  sr_buffer_32_1 f696(.wen(f696_wen), .wdata(f696_wdata), .clk(f696_clk), .rst(f696_rst), .rdata(f696_rdata));
  assign f696_clk = clk;
  assign f696_rst = rst;
  // Bindings to f696

  // f698
  logic [0:0] f698_wen;
  logic [31:0] f698_wdata;
  logic [0:0] f698_clk;
  logic [0:0] f698_rst;
  logic [31:0] f698_rdata;
  sr_buffer_32_1 f698(.wen(f698_wen), .wdata(f698_wdata), .clk(f698_clk), .rst(f698_rst), .rdata(f698_rdata));
  assign f698_clk = clk;
  assign f698_rst = rst;
  // Bindings to f698

  // f700
  logic [0:0] f700_wen;
  logic [31:0] f700_wdata;
  logic [0:0] f700_clk;
  logic [0:0] f700_rst;
  logic [31:0] f700_rdata;
  sr_buffer_32_1 f700(.wen(f700_wen), .wdata(f700_wdata), .clk(f700_clk), .rst(f700_rst), .rdata(f700_rdata));
  assign f700_clk = clk;
  assign f700_rst = rst;
  // Bindings to f700

  // f702
  logic [0:0] f702_wen;
  logic [31:0] f702_wdata;
  logic [0:0] f702_clk;
  logic [0:0] f702_rst;
  logic [31:0] f702_rdata;
  sr_buffer_32_1 f702(.wen(f702_wen), .wdata(f702_wdata), .clk(f702_clk), .rst(f702_rst), .rdata(f702_rdata));
  assign f702_clk = clk;
  assign f702_rst = rst;
  // Bindings to f702

  // f704
  logic [0:0] f704_wen;
  logic [31:0] f704_wdata;
  logic [0:0] f704_clk;
  logic [0:0] f704_rst;
  logic [31:0] f704_rdata;
  sr_buffer_32_1 f704(.wen(f704_wen), .wdata(f704_wdata), .clk(f704_clk), .rst(f704_rst), .rdata(f704_rdata));
  assign f704_clk = clk;
  assign f704_rst = rst;
  // Bindings to f704

  // f706
  logic [0:0] f706_wen;
  logic [31:0] f706_wdata;
  logic [0:0] f706_clk;
  logic [0:0] f706_rst;
  logic [31:0] f706_rdata;
  sr_buffer_32_1 f706(.wen(f706_wen), .wdata(f706_wdata), .clk(f706_clk), .rst(f706_rst), .rdata(f706_rdata));
  assign f706_clk = clk;
  assign f706_rst = rst;
  // Bindings to f706

  // f708
  logic [0:0] f708_wen;
  logic [31:0] f708_wdata;
  logic [0:0] f708_clk;
  logic [0:0] f708_rst;
  logic [31:0] f708_rdata;
  sr_buffer_32_1 f708(.wen(f708_wen), .wdata(f708_wdata), .clk(f708_clk), .rst(f708_rst), .rdata(f708_rdata));
  assign f708_clk = clk;
  assign f708_rst = rst;
  // Bindings to f708

  // f710
  logic [0:0] f710_wen;
  logic [31:0] f710_wdata;
  logic [0:0] f710_clk;
  logic [0:0] f710_rst;
  logic [31:0] f710_rdata;
  sr_buffer_32_1 f710(.wen(f710_wen), .wdata(f710_wdata), .clk(f710_clk), .rst(f710_rst), .rdata(f710_rdata));
  assign f710_clk = clk;
  assign f710_rst = rst;
  // Bindings to f710

  // f712
  logic [0:0] f712_wen;
  logic [31:0] f712_wdata;
  logic [0:0] f712_clk;
  logic [0:0] f712_rst;
  logic [31:0] f712_rdata;
  sr_buffer_32_1 f712(.wen(f712_wen), .wdata(f712_wdata), .clk(f712_clk), .rst(f712_rst), .rdata(f712_rdata));
  assign f712_clk = clk;
  assign f712_rst = rst;
  // Bindings to f712

  // f714
  logic [0:0] f714_wen;
  logic [31:0] f714_wdata;
  logic [0:0] f714_clk;
  logic [0:0] f714_rst;
  logic [31:0] f714_rdata;
  sr_buffer_32_1 f714(.wen(f714_wen), .wdata(f714_wdata), .clk(f714_clk), .rst(f714_rst), .rdata(f714_rdata));
  assign f714_clk = clk;
  assign f714_rst = rst;
  // Bindings to f714

  // f716
  logic [0:0] f716_wen;
  logic [31:0] f716_wdata;
  logic [0:0] f716_clk;
  logic [0:0] f716_rst;
  logic [31:0] f716_rdata;
  sr_buffer_32_1 f716(.wen(f716_wen), .wdata(f716_wdata), .clk(f716_clk), .rst(f716_rst), .rdata(f716_rdata));
  assign f716_clk = clk;
  assign f716_rst = rst;
  // Bindings to f716

  // f718
  logic [0:0] f718_wen;
  logic [31:0] f718_wdata;
  logic [0:0] f718_clk;
  logic [0:0] f718_rst;
  logic [31:0] f718_rdata;
  sr_buffer_32_1 f718(.wen(f718_wen), .wdata(f718_wdata), .clk(f718_clk), .rst(f718_rst), .rdata(f718_rdata));
  assign f718_clk = clk;
  assign f718_rst = rst;
  // Bindings to f718

  // f720
  logic [0:0] f720_wen;
  logic [31:0] f720_wdata;
  logic [0:0] f720_clk;
  logic [0:0] f720_rst;
  logic [31:0] f720_rdata;
  sr_buffer_32_1 f720(.wen(f720_wen), .wdata(f720_wdata), .clk(f720_clk), .rst(f720_rst), .rdata(f720_rdata));
  assign f720_clk = clk;
  assign f720_rst = rst;
  // Bindings to f720

  // f722
  logic [0:0] f722_wen;
  logic [31:0] f722_wdata;
  logic [0:0] f722_clk;
  logic [0:0] f722_rst;
  logic [31:0] f722_rdata;
  sr_buffer_32_1 f722(.wen(f722_wen), .wdata(f722_wdata), .clk(f722_clk), .rst(f722_rst), .rdata(f722_rdata));
  assign f722_clk = clk;
  assign f722_rst = rst;
  // Bindings to f722

  // f724
  logic [0:0] f724_wen;
  logic [31:0] f724_wdata;
  logic [0:0] f724_clk;
  logic [0:0] f724_rst;
  logic [31:0] f724_rdata;
  sr_buffer_32_1 f724(.wen(f724_wen), .wdata(f724_wdata), .clk(f724_clk), .rst(f724_rst), .rdata(f724_rdata));
  assign f724_clk = clk;
  assign f724_rst = rst;
  // Bindings to f724

  // f726
  logic [0:0] f726_wen;
  logic [31:0] f726_wdata;
  logic [0:0] f726_clk;
  logic [0:0] f726_rst;
  logic [31:0] f726_rdata;
  sr_buffer_32_1 f726(.wen(f726_wen), .wdata(f726_wdata), .clk(f726_clk), .rst(f726_rst), .rdata(f726_rdata));
  assign f726_clk = clk;
  assign f726_rst = rst;
  // Bindings to f726

  // f728
  logic [0:0] f728_wen;
  logic [31:0] f728_wdata;
  logic [0:0] f728_clk;
  logic [0:0] f728_rst;
  logic [31:0] f728_rdata;
  sr_buffer_32_1 f728(.wen(f728_wen), .wdata(f728_wdata), .clk(f728_clk), .rst(f728_rst), .rdata(f728_rdata));
  assign f728_clk = clk;
  assign f728_rst = rst;
  // Bindings to f728

  // f730
  logic [0:0] f730_wen;
  logic [31:0] f730_wdata;
  logic [0:0] f730_clk;
  logic [0:0] f730_rst;
  logic [31:0] f730_rdata;
  sr_buffer_32_1 f730(.wen(f730_wen), .wdata(f730_wdata), .clk(f730_clk), .rst(f730_rst), .rdata(f730_rdata));
  assign f730_clk = clk;
  assign f730_rst = rst;
  // Bindings to f730

  // f732
  logic [0:0] f732_wen;
  logic [31:0] f732_wdata;
  logic [0:0] f732_clk;
  logic [0:0] f732_rst;
  logic [31:0] f732_rdata;
  sr_buffer_32_1 f732(.wen(f732_wen), .wdata(f732_wdata), .clk(f732_clk), .rst(f732_rst), .rdata(f732_rdata));
  assign f732_clk = clk;
  assign f732_rst = rst;
  // Bindings to f732

  // f734
  logic [0:0] f734_wen;
  logic [31:0] f734_wdata;
  logic [0:0] f734_clk;
  logic [0:0] f734_rst;
  logic [31:0] f734_rdata;
  sr_buffer_32_1 f734(.wen(f734_wen), .wdata(f734_wdata), .clk(f734_clk), .rst(f734_rst), .rdata(f734_rdata));
  assign f734_clk = clk;
  assign f734_rst = rst;
  // Bindings to f734

  // f736
  logic [0:0] f736_wen;
  logic [31:0] f736_wdata;
  logic [0:0] f736_clk;
  logic [0:0] f736_rst;
  logic [31:0] f736_rdata;
  sr_buffer_32_1 f736(.wen(f736_wen), .wdata(f736_wdata), .clk(f736_clk), .rst(f736_rst), .rdata(f736_rdata));
  assign f736_clk = clk;
  assign f736_rst = rst;
  // Bindings to f736

  // f738
  logic [0:0] f738_wen;
  logic [31:0] f738_wdata;
  logic [0:0] f738_clk;
  logic [0:0] f738_rst;
  logic [31:0] f738_rdata;
  sr_buffer_32_1 f738(.wen(f738_wen), .wdata(f738_wdata), .clk(f738_clk), .rst(f738_rst), .rdata(f738_rdata));
  assign f738_clk = clk;
  assign f738_rst = rst;
  // Bindings to f738

  // f740
  logic [0:0] f740_wen;
  logic [31:0] f740_wdata;
  logic [0:0] f740_clk;
  logic [0:0] f740_rst;
  logic [31:0] f740_rdata;
  sr_buffer_32_1 f740(.wen(f740_wen), .wdata(f740_wdata), .clk(f740_clk), .rst(f740_rst), .rdata(f740_rdata));
  assign f740_clk = clk;
  assign f740_rst = rst;
  // Bindings to f740

  // f742
  logic [0:0] f742_wen;
  logic [31:0] f742_wdata;
  logic [0:0] f742_clk;
  logic [0:0] f742_rst;
  logic [31:0] f742_rdata;
  sr_buffer_32_1 f742(.wen(f742_wen), .wdata(f742_wdata), .clk(f742_clk), .rst(f742_rst), .rdata(f742_rdata));
  assign f742_clk = clk;
  assign f742_rst = rst;
  // Bindings to f742

  // f744
  logic [0:0] f744_wen;
  logic [31:0] f744_wdata;
  logic [0:0] f744_clk;
  logic [0:0] f744_rst;
  logic [31:0] f744_rdata;
  sr_buffer_32_1 f744(.wen(f744_wen), .wdata(f744_wdata), .clk(f744_clk), .rst(f744_rst), .rdata(f744_rdata));
  assign f744_clk = clk;
  assign f744_rst = rst;
  // Bindings to f744

  // f746
  logic [0:0] f746_wen;
  logic [31:0] f746_wdata;
  logic [0:0] f746_clk;
  logic [0:0] f746_rst;
  logic [31:0] f746_rdata;
  sr_buffer_32_1 f746(.wen(f746_wen), .wdata(f746_wdata), .clk(f746_clk), .rst(f746_rst), .rdata(f746_rdata));
  assign f746_clk = clk;
  assign f746_rst = rst;
  // Bindings to f746

  // f748
  logic [0:0] f748_wen;
  logic [31:0] f748_wdata;
  logic [0:0] f748_clk;
  logic [0:0] f748_rst;
  logic [31:0] f748_rdata;
  sr_buffer_32_1 f748(.wen(f748_wen), .wdata(f748_wdata), .clk(f748_clk), .rst(f748_rst), .rdata(f748_rdata));
  assign f748_clk = clk;
  assign f748_rst = rst;
  // Bindings to f748

  // f750
  logic [0:0] f750_wen;
  logic [31:0] f750_wdata;
  logic [0:0] f750_clk;
  logic [0:0] f750_rst;
  logic [31:0] f750_rdata;
  sr_buffer_32_1 f750(.wen(f750_wen), .wdata(f750_wdata), .clk(f750_clk), .rst(f750_rst), .rdata(f750_rdata));
  assign f750_clk = clk;
  assign f750_rst = rst;
  // Bindings to f750

  // f752
  logic [0:0] f752_wen;
  logic [31:0] f752_wdata;
  logic [0:0] f752_clk;
  logic [0:0] f752_rst;
  logic [31:0] f752_rdata;
  sr_buffer_32_1 f752(.wen(f752_wen), .wdata(f752_wdata), .clk(f752_clk), .rst(f752_rst), .rdata(f752_rdata));
  assign f752_clk = clk;
  assign f752_rst = rst;
  // Bindings to f752

  // f754
  logic [0:0] f754_wen;
  logic [31:0] f754_wdata;
  logic [0:0] f754_clk;
  logic [0:0] f754_rst;
  logic [31:0] f754_rdata;
  sr_buffer_32_1 f754(.wen(f754_wen), .wdata(f754_wdata), .clk(f754_clk), .rst(f754_rst), .rdata(f754_rdata));
  assign f754_clk = clk;
  assign f754_rst = rst;
  // Bindings to f754

  // f756
  logic [0:0] f756_wen;
  logic [31:0] f756_wdata;
  logic [0:0] f756_clk;
  logic [0:0] f756_rst;
  logic [31:0] f756_rdata;
  sr_buffer_32_1 f756(.wen(f756_wen), .wdata(f756_wdata), .clk(f756_clk), .rst(f756_rst), .rdata(f756_rdata));
  assign f756_clk = clk;
  assign f756_rst = rst;
  // Bindings to f756

  // f758
  logic [0:0] f758_wen;
  logic [31:0] f758_wdata;
  logic [0:0] f758_clk;
  logic [0:0] f758_rst;
  logic [31:0] f758_rdata;
  sr_buffer_32_1 f758(.wen(f758_wen), .wdata(f758_wdata), .clk(f758_clk), .rst(f758_rst), .rdata(f758_rdata));
  assign f758_clk = clk;
  assign f758_rst = rst;
  // Bindings to f758

  // f760
  logic [0:0] f760_wen;
  logic [31:0] f760_wdata;
  logic [0:0] f760_clk;
  logic [0:0] f760_rst;
  logic [31:0] f760_rdata;
  sr_buffer_32_1 f760(.wen(f760_wen), .wdata(f760_wdata), .clk(f760_clk), .rst(f760_rst), .rdata(f760_rdata));
  assign f760_clk = clk;
  assign f760_rst = rst;
  // Bindings to f760

  // f762
  logic [0:0] f762_wen;
  logic [31:0] f762_wdata;
  logic [0:0] f762_clk;
  logic [0:0] f762_rst;
  logic [31:0] f762_rdata;
  sr_buffer_32_1 f762(.wen(f762_wen), .wdata(f762_wdata), .clk(f762_clk), .rst(f762_rst), .rdata(f762_rdata));
  assign f762_clk = clk;
  assign f762_rst = rst;
  // Bindings to f762

  // f764
  logic [0:0] f764_wen;
  logic [31:0] f764_wdata;
  logic [0:0] f764_clk;
  logic [0:0] f764_rst;
  logic [31:0] f764_rdata;
  sr_buffer_32_1 f764(.wen(f764_wen), .wdata(f764_wdata), .clk(f764_clk), .rst(f764_rst), .rdata(f764_rdata));
  assign f764_clk = clk;
  assign f764_rst = rst;
  // Bindings to f764

  // f766
  logic [0:0] f766_wen;
  logic [31:0] f766_wdata;
  logic [0:0] f766_clk;
  logic [0:0] f766_rst;
  logic [31:0] f766_rdata;
  sr_buffer_32_1 f766(.wen(f766_wen), .wdata(f766_wdata), .clk(f766_clk), .rst(f766_rst), .rdata(f766_rdata));
  assign f766_clk = clk;
  assign f766_rst = rst;
  // Bindings to f766

  // f768
  logic [0:0] f768_wen;
  logic [31:0] f768_wdata;
  logic [0:0] f768_clk;
  logic [0:0] f768_rst;
  logic [31:0] f768_rdata;
  sr_buffer_32_1 f768(.wen(f768_wen), .wdata(f768_wdata), .clk(f768_clk), .rst(f768_rst), .rdata(f768_rdata));
  assign f768_clk = clk;
  assign f768_rst = rst;
  // Bindings to f768

  // f770
  logic [0:0] f770_wen;
  logic [31:0] f770_wdata;
  logic [0:0] f770_clk;
  logic [0:0] f770_rst;
  logic [31:0] f770_rdata;
  sr_buffer_32_1 f770(.wen(f770_wen), .wdata(f770_wdata), .clk(f770_clk), .rst(f770_rst), .rdata(f770_rdata));
  assign f770_clk = clk;
  assign f770_rst = rst;
  // Bindings to f770

  // f772
  logic [0:0] f772_wen;
  logic [31:0] f772_wdata;
  logic [0:0] f772_clk;
  logic [0:0] f772_rst;
  logic [31:0] f772_rdata;
  sr_buffer_32_1 f772(.wen(f772_wen), .wdata(f772_wdata), .clk(f772_clk), .rst(f772_rst), .rdata(f772_rdata));
  assign f772_clk = clk;
  assign f772_rst = rst;
  // Bindings to f772

  // f774
  logic [0:0] f774_wen;
  logic [31:0] f774_wdata;
  logic [0:0] f774_clk;
  logic [0:0] f774_rst;
  logic [31:0] f774_rdata;
  sr_buffer_32_1 f774(.wen(f774_wen), .wdata(f774_wdata), .clk(f774_clk), .rst(f774_rst), .rdata(f774_rdata));
  assign f774_clk = clk;
  assign f774_rst = rst;
  // Bindings to f774

  // f776
  logic [0:0] f776_wen;
  logic [31:0] f776_wdata;
  logic [0:0] f776_clk;
  logic [0:0] f776_rst;
  logic [31:0] f776_rdata;
  sr_buffer_32_1 f776(.wen(f776_wen), .wdata(f776_wdata), .clk(f776_clk), .rst(f776_rst), .rdata(f776_rdata));
  assign f776_clk = clk;
  assign f776_rst = rst;
  // Bindings to f776

  // f778
  logic [0:0] f778_wen;
  logic [31:0] f778_wdata;
  logic [0:0] f778_clk;
  logic [0:0] f778_rst;
  logic [31:0] f778_rdata;
  sr_buffer_32_1 f778(.wen(f778_wen), .wdata(f778_wdata), .clk(f778_clk), .rst(f778_rst), .rdata(f778_rdata));
  assign f778_clk = clk;
  assign f778_rst = rst;
  // Bindings to f778

  // f780
  logic [0:0] f780_wen;
  logic [31:0] f780_wdata;
  logic [0:0] f780_clk;
  logic [0:0] f780_rst;
  logic [31:0] f780_rdata;
  sr_buffer_32_1 f780(.wen(f780_wen), .wdata(f780_wdata), .clk(f780_clk), .rst(f780_rst), .rdata(f780_rdata));
  assign f780_clk = clk;
  assign f780_rst = rst;
  // Bindings to f780

  // f782
  logic [0:0] f782_wen;
  logic [31:0] f782_wdata;
  logic [0:0] f782_clk;
  logic [0:0] f782_rst;
  logic [31:0] f782_rdata;
  sr_buffer_32_1 f782(.wen(f782_wen), .wdata(f782_wdata), .clk(f782_clk), .rst(f782_rst), .rdata(f782_rdata));
  assign f782_clk = clk;
  assign f782_rst = rst;
  // Bindings to f782

  // f784
  logic [0:0] f784_wen;
  logic [31:0] f784_wdata;
  logic [0:0] f784_clk;
  logic [0:0] f784_rst;
  logic [31:0] f784_rdata;
  sr_buffer_32_1 f784(.wen(f784_wen), .wdata(f784_wdata), .clk(f784_clk), .rst(f784_rst), .rdata(f784_rdata));
  assign f784_clk = clk;
  assign f784_rst = rst;
  // Bindings to f784

  // f786
  logic [0:0] f786_wen;
  logic [31:0] f786_wdata;
  logic [0:0] f786_clk;
  logic [0:0] f786_rst;
  logic [31:0] f786_rdata;
  sr_buffer_32_1 f786(.wen(f786_wen), .wdata(f786_wdata), .clk(f786_clk), .rst(f786_rst), .rdata(f786_rdata));
  assign f786_clk = clk;
  assign f786_rst = rst;
  // Bindings to f786

  // f788
  logic [0:0] f788_wen;
  logic [31:0] f788_wdata;
  logic [0:0] f788_clk;
  logic [0:0] f788_rst;
  logic [31:0] f788_rdata;
  sr_buffer_32_1 f788(.wen(f788_wen), .wdata(f788_wdata), .clk(f788_clk), .rst(f788_rst), .rdata(f788_rdata));
  assign f788_clk = clk;
  assign f788_rst = rst;
  // Bindings to f788

  // f790
  logic [0:0] f790_wen;
  logic [31:0] f790_wdata;
  logic [0:0] f790_clk;
  logic [0:0] f790_rst;
  logic [31:0] f790_rdata;
  sr_buffer_32_1 f790(.wen(f790_wen), .wdata(f790_wdata), .clk(f790_clk), .rst(f790_rst), .rdata(f790_rdata));
  assign f790_clk = clk;
  assign f790_rst = rst;
  // Bindings to f790

  // f792
  logic [0:0] f792_wen;
  logic [31:0] f792_wdata;
  logic [0:0] f792_clk;
  logic [0:0] f792_rst;
  logic [31:0] f792_rdata;
  sr_buffer_32_1 f792(.wen(f792_wen), .wdata(f792_wdata), .clk(f792_clk), .rst(f792_rst), .rdata(f792_rdata));
  assign f792_clk = clk;
  assign f792_rst = rst;
  // Bindings to f792

  // f794
  logic [0:0] f794_wen;
  logic [31:0] f794_wdata;
  logic [0:0] f794_clk;
  logic [0:0] f794_rst;
  logic [31:0] f794_rdata;
  sr_buffer_32_1 f794(.wen(f794_wen), .wdata(f794_wdata), .clk(f794_clk), .rst(f794_rst), .rdata(f794_rdata));
  assign f794_clk = clk;
  assign f794_rst = rst;
  // Bindings to f794

  // f796
  logic [0:0] f796_wen;
  logic [31:0] f796_wdata;
  logic [0:0] f796_clk;
  logic [0:0] f796_rst;
  logic [31:0] f796_rdata;
  sr_buffer_32_1 f796(.wen(f796_wen), .wdata(f796_wdata), .clk(f796_clk), .rst(f796_rst), .rdata(f796_rdata));
  assign f796_clk = clk;
  assign f796_rst = rst;
  // Bindings to f796

  // f798
  logic [0:0] f798_wen;
  logic [31:0] f798_wdata;
  logic [0:0] f798_clk;
  logic [0:0] f798_rst;
  logic [31:0] f798_rdata;
  sr_buffer_32_1 f798(.wen(f798_wen), .wdata(f798_wdata), .clk(f798_clk), .rst(f798_rst), .rdata(f798_rdata));
  assign f798_clk = clk;
  assign f798_rst = rst;
  // Bindings to f798

  // f800
  logic [0:0] f800_wen;
  logic [31:0] f800_wdata;
  logic [0:0] f800_clk;
  logic [0:0] f800_rst;
  logic [31:0] f800_rdata;
  sr_buffer_32_1 f800(.wen(f800_wen), .wdata(f800_wdata), .clk(f800_clk), .rst(f800_rst), .rdata(f800_rdata));
  assign f800_clk = clk;
  assign f800_rst = rst;
  // Bindings to f800

  // f802
  logic [0:0] f802_wen;
  logic [31:0] f802_wdata;
  logic [0:0] f802_clk;
  logic [0:0] f802_rst;
  logic [31:0] f802_rdata;
  sr_buffer_32_1 f802(.wen(f802_wen), .wdata(f802_wdata), .clk(f802_clk), .rst(f802_rst), .rdata(f802_rdata));
  assign f802_clk = clk;
  assign f802_rst = rst;
  // Bindings to f802

  // f804
  logic [0:0] f804_wen;
  logic [31:0] f804_wdata;
  logic [0:0] f804_clk;
  logic [0:0] f804_rst;
  logic [31:0] f804_rdata;
  sr_buffer_32_1 f804(.wen(f804_wen), .wdata(f804_wdata), .clk(f804_clk), .rst(f804_rst), .rdata(f804_rdata));
  assign f804_clk = clk;
  assign f804_rst = rst;
  // Bindings to f804

  // f806
  logic [0:0] f806_wen;
  logic [31:0] f806_wdata;
  logic [0:0] f806_clk;
  logic [0:0] f806_rst;
  logic [31:0] f806_rdata;
  sr_buffer_32_1 f806(.wen(f806_wen), .wdata(f806_wdata), .clk(f806_clk), .rst(f806_rst), .rdata(f806_rdata));
  assign f806_clk = clk;
  assign f806_rst = rst;
  // Bindings to f806

  // f808
  logic [0:0] f808_wen;
  logic [31:0] f808_wdata;
  logic [0:0] f808_clk;
  logic [0:0] f808_rst;
  logic [31:0] f808_rdata;
  sr_buffer_32_1 f808(.wen(f808_wen), .wdata(f808_wdata), .clk(f808_clk), .rst(f808_rst), .rdata(f808_rdata));
  assign f808_clk = clk;
  assign f808_rst = rst;
  // Bindings to f808

  // f810
  logic [0:0] f810_wen;
  logic [31:0] f810_wdata;
  logic [0:0] f810_clk;
  logic [0:0] f810_rst;
  logic [31:0] f810_rdata;
  sr_buffer_32_1 f810(.wen(f810_wen), .wdata(f810_wdata), .clk(f810_clk), .rst(f810_rst), .rdata(f810_rdata));
  assign f810_clk = clk;
  assign f810_rst = rst;
  // Bindings to f810

  // f812
  logic [0:0] f812_wen;
  logic [31:0] f812_wdata;
  logic [0:0] f812_clk;
  logic [0:0] f812_rst;
  logic [31:0] f812_rdata;
  sr_buffer_32_1 f812(.wen(f812_wen), .wdata(f812_wdata), .clk(f812_clk), .rst(f812_rst), .rdata(f812_rdata));
  assign f812_clk = clk;
  assign f812_rst = rst;
  // Bindings to f812

  // f814
  logic [0:0] f814_wen;
  logic [31:0] f814_wdata;
  logic [0:0] f814_clk;
  logic [0:0] f814_rst;
  logic [31:0] f814_rdata;
  sr_buffer_32_1 f814(.wen(f814_wen), .wdata(f814_wdata), .clk(f814_clk), .rst(f814_rst), .rdata(f814_rdata));
  assign f814_clk = clk;
  assign f814_rst = rst;
  // Bindings to f814

  // f816
  logic [0:0] f816_wen;
  logic [31:0] f816_wdata;
  logic [0:0] f816_clk;
  logic [0:0] f816_rst;
  logic [31:0] f816_rdata;
  sr_buffer_32_1 f816(.wen(f816_wen), .wdata(f816_wdata), .clk(f816_clk), .rst(f816_rst), .rdata(f816_rdata));
  assign f816_clk = clk;
  assign f816_rst = rst;
  // Bindings to f816

  // f818
  logic [0:0] f818_wen;
  logic [31:0] f818_wdata;
  logic [0:0] f818_clk;
  logic [0:0] f818_rst;
  logic [31:0] f818_rdata;
  sr_buffer_32_1 f818(.wen(f818_wen), .wdata(f818_wdata), .clk(f818_clk), .rst(f818_rst), .rdata(f818_rdata));
  assign f818_clk = clk;
  assign f818_rst = rst;
  // Bindings to f818

  // f820
  logic [0:0] f820_wen;
  logic [31:0] f820_wdata;
  logic [0:0] f820_clk;
  logic [0:0] f820_rst;
  logic [31:0] f820_rdata;
  sr_buffer_32_1 f820(.wen(f820_wen), .wdata(f820_wdata), .clk(f820_clk), .rst(f820_rst), .rdata(f820_rdata));
  assign f820_clk = clk;
  assign f820_rst = rst;
  // Bindings to f820

  // f822
  logic [0:0] f822_wen;
  logic [31:0] f822_wdata;
  logic [0:0] f822_clk;
  logic [0:0] f822_rst;
  logic [31:0] f822_rdata;
  sr_buffer_32_1 f822(.wen(f822_wen), .wdata(f822_wdata), .clk(f822_clk), .rst(f822_rst), .rdata(f822_rdata));
  assign f822_clk = clk;
  assign f822_rst = rst;
  // Bindings to f822

  // f824
  logic [0:0] f824_wen;
  logic [31:0] f824_wdata;
  logic [0:0] f824_clk;
  logic [0:0] f824_rst;
  logic [31:0] f824_rdata;
  sr_buffer_32_1 f824(.wen(f824_wen), .wdata(f824_wdata), .clk(f824_clk), .rst(f824_rst), .rdata(f824_rdata));
  assign f824_clk = clk;
  assign f824_rst = rst;
  // Bindings to f824

  // f826
  logic [0:0] f826_wen;
  logic [31:0] f826_wdata;
  logic [0:0] f826_clk;
  logic [0:0] f826_rst;
  logic [31:0] f826_rdata;
  sr_buffer_32_1 f826(.wen(f826_wen), .wdata(f826_wdata), .clk(f826_clk), .rst(f826_rst), .rdata(f826_rdata));
  assign f826_clk = clk;
  assign f826_rst = rst;
  // Bindings to f826

  // f828
  logic [0:0] f828_wen;
  logic [31:0] f828_wdata;
  logic [0:0] f828_clk;
  logic [0:0] f828_rst;
  logic [31:0] f828_rdata;
  sr_buffer_32_1 f828(.wen(f828_wen), .wdata(f828_wdata), .clk(f828_clk), .rst(f828_rst), .rdata(f828_rdata));
  assign f828_clk = clk;
  assign f828_rst = rst;
  // Bindings to f828

  // f830
  logic [0:0] f830_wen;
  logic [31:0] f830_wdata;
  logic [0:0] f830_clk;
  logic [0:0] f830_rst;
  logic [31:0] f830_rdata;
  sr_buffer_32_1 f830(.wen(f830_wen), .wdata(f830_wdata), .clk(f830_clk), .rst(f830_rst), .rdata(f830_rdata));
  assign f830_clk = clk;
  assign f830_rst = rst;
  // Bindings to f830

  // f832
  logic [0:0] f832_wen;
  logic [31:0] f832_wdata;
  logic [0:0] f832_clk;
  logic [0:0] f832_rst;
  logic [31:0] f832_rdata;
  sr_buffer_32_1 f832(.wen(f832_wen), .wdata(f832_wdata), .clk(f832_clk), .rst(f832_rst), .rdata(f832_rdata));
  assign f832_clk = clk;
  assign f832_rst = rst;
  // Bindings to f832

  // f834
  logic [0:0] f834_wen;
  logic [31:0] f834_wdata;
  logic [0:0] f834_clk;
  logic [0:0] f834_rst;
  logic [31:0] f834_rdata;
  sr_buffer_32_1 f834(.wen(f834_wen), .wdata(f834_wdata), .clk(f834_clk), .rst(f834_rst), .rdata(f834_rdata));
  assign f834_clk = clk;
  assign f834_rst = rst;
  // Bindings to f834

  // f836
  logic [0:0] f836_wen;
  logic [31:0] f836_wdata;
  logic [0:0] f836_clk;
  logic [0:0] f836_rst;
  logic [31:0] f836_rdata;
  sr_buffer_32_1 f836(.wen(f836_wen), .wdata(f836_wdata), .clk(f836_clk), .rst(f836_rst), .rdata(f836_rdata));
  assign f836_clk = clk;
  assign f836_rst = rst;
  // Bindings to f836

  // f838
  logic [0:0] f838_wen;
  logic [31:0] f838_wdata;
  logic [0:0] f838_clk;
  logic [0:0] f838_rst;
  logic [31:0] f838_rdata;
  sr_buffer_32_1 f838(.wen(f838_wen), .wdata(f838_wdata), .clk(f838_clk), .rst(f838_rst), .rdata(f838_rdata));
  assign f838_clk = clk;
  assign f838_rst = rst;
  // Bindings to f838

  // f840
  logic [0:0] f840_wen;
  logic [31:0] f840_wdata;
  logic [0:0] f840_clk;
  logic [0:0] f840_rst;
  logic [31:0] f840_rdata;
  sr_buffer_32_1 f840(.wen(f840_wen), .wdata(f840_wdata), .clk(f840_clk), .rst(f840_rst), .rdata(f840_rdata));
  assign f840_clk = clk;
  assign f840_rst = rst;
  // Bindings to f840

  // f842
  logic [0:0] f842_wen;
  logic [31:0] f842_wdata;
  logic [0:0] f842_clk;
  logic [0:0] f842_rst;
  logic [31:0] f842_rdata;
  sr_buffer_32_1 f842(.wen(f842_wen), .wdata(f842_wdata), .clk(f842_clk), .rst(f842_rst), .rdata(f842_rdata));
  assign f842_clk = clk;
  assign f842_rst = rst;
  // Bindings to f842

  // f844
  logic [0:0] f844_wen;
  logic [31:0] f844_wdata;
  logic [0:0] f844_clk;
  logic [0:0] f844_rst;
  logic [31:0] f844_rdata;
  sr_buffer_32_1 f844(.wen(f844_wen), .wdata(f844_wdata), .clk(f844_clk), .rst(f844_rst), .rdata(f844_rdata));
  assign f844_clk = clk;
  assign f844_rst = rst;
  // Bindings to f844

  // f846
  logic [0:0] f846_wen;
  logic [31:0] f846_wdata;
  logic [0:0] f846_clk;
  logic [0:0] f846_rst;
  logic [31:0] f846_rdata;
  sr_buffer_32_1 f846(.wen(f846_wen), .wdata(f846_wdata), .clk(f846_clk), .rst(f846_rst), .rdata(f846_rdata));
  assign f846_clk = clk;
  assign f846_rst = rst;
  // Bindings to f846

  // f848
  logic [0:0] f848_wen;
  logic [31:0] f848_wdata;
  logic [0:0] f848_clk;
  logic [0:0] f848_rst;
  logic [31:0] f848_rdata;
  sr_buffer_32_1 f848(.wen(f848_wen), .wdata(f848_wdata), .clk(f848_clk), .rst(f848_rst), .rdata(f848_rdata));
  assign f848_clk = clk;
  assign f848_rst = rst;
  // Bindings to f848

  // f850
  logic [0:0] f850_wen;
  logic [31:0] f850_wdata;
  logic [0:0] f850_clk;
  logic [0:0] f850_rst;
  logic [31:0] f850_rdata;
  sr_buffer_32_1 f850(.wen(f850_wen), .wdata(f850_wdata), .clk(f850_clk), .rst(f850_rst), .rdata(f850_rdata));
  assign f850_clk = clk;
  assign f850_rst = rst;
  // Bindings to f850

  // f852
  logic [0:0] f852_wen;
  logic [31:0] f852_wdata;
  logic [0:0] f852_clk;
  logic [0:0] f852_rst;
  logic [31:0] f852_rdata;
  sr_buffer_32_1 f852(.wen(f852_wen), .wdata(f852_wdata), .clk(f852_clk), .rst(f852_rst), .rdata(f852_rdata));
  assign f852_clk = clk;
  assign f852_rst = rst;
  // Bindings to f852

  // f854
  logic [0:0] f854_wen;
  logic [31:0] f854_wdata;
  logic [0:0] f854_clk;
  logic [0:0] f854_rst;
  logic [31:0] f854_rdata;
  sr_buffer_32_1 f854(.wen(f854_wen), .wdata(f854_wdata), .clk(f854_clk), .rst(f854_rst), .rdata(f854_rdata));
  assign f854_clk = clk;
  assign f854_rst = rst;
  // Bindings to f854

  // f856
  logic [0:0] f856_wen;
  logic [31:0] f856_wdata;
  logic [0:0] f856_clk;
  logic [0:0] f856_rst;
  logic [31:0] f856_rdata;
  sr_buffer_32_1 f856(.wen(f856_wen), .wdata(f856_wdata), .clk(f856_clk), .rst(f856_rst), .rdata(f856_rdata));
  assign f856_clk = clk;
  assign f856_rst = rst;
  // Bindings to f856

  // f858
  logic [0:0] f858_wen;
  logic [31:0] f858_wdata;
  logic [0:0] f858_clk;
  logic [0:0] f858_rst;
  logic [31:0] f858_rdata;
  sr_buffer_32_1 f858(.wen(f858_wen), .wdata(f858_wdata), .clk(f858_clk), .rst(f858_rst), .rdata(f858_rdata));
  assign f858_clk = clk;
  assign f858_rst = rst;
  // Bindings to f858

  // f860
  logic [0:0] f860_wen;
  logic [31:0] f860_wdata;
  logic [0:0] f860_clk;
  logic [0:0] f860_rst;
  logic [31:0] f860_rdata;
  sr_buffer_32_1 f860(.wen(f860_wen), .wdata(f860_wdata), .clk(f860_clk), .rst(f860_rst), .rdata(f860_rdata));
  assign f860_clk = clk;
  assign f860_rst = rst;
  // Bindings to f860

  // f862
  logic [0:0] f862_wen;
  logic [31:0] f862_wdata;
  logic [0:0] f862_clk;
  logic [0:0] f862_rst;
  logic [31:0] f862_rdata;
  sr_buffer_32_1 f862(.wen(f862_wen), .wdata(f862_wdata), .clk(f862_clk), .rst(f862_rst), .rdata(f862_rdata));
  assign f862_clk = clk;
  assign f862_rst = rst;
  // Bindings to f862

  // f864
  logic [0:0] f864_wen;
  logic [31:0] f864_wdata;
  logic [0:0] f864_clk;
  logic [0:0] f864_rst;
  logic [31:0] f864_rdata;
  sr_buffer_32_1 f864(.wen(f864_wen), .wdata(f864_wdata), .clk(f864_clk), .rst(f864_rst), .rdata(f864_rdata));
  assign f864_clk = clk;
  assign f864_rst = rst;
  // Bindings to f864

  // f866
  logic [0:0] f866_wen;
  logic [31:0] f866_wdata;
  logic [0:0] f866_clk;
  logic [0:0] f866_rst;
  logic [31:0] f866_rdata;
  sr_buffer_32_1 f866(.wen(f866_wen), .wdata(f866_wdata), .clk(f866_clk), .rst(f866_rst), .rdata(f866_rdata));
  assign f866_clk = clk;
  assign f866_rst = rst;
  // Bindings to f866

  // f868
  logic [0:0] f868_wen;
  logic [31:0] f868_wdata;
  logic [0:0] f868_clk;
  logic [0:0] f868_rst;
  logic [31:0] f868_rdata;
  sr_buffer_32_1 f868(.wen(f868_wen), .wdata(f868_wdata), .clk(f868_clk), .rst(f868_rst), .rdata(f868_rdata));
  assign f868_clk = clk;
  assign f868_rst = rst;
  // Bindings to f868

  // f870
  logic [0:0] f870_wen;
  logic [31:0] f870_wdata;
  logic [0:0] f870_clk;
  logic [0:0] f870_rst;
  logic [31:0] f870_rdata;
  sr_buffer_32_1 f870(.wen(f870_wen), .wdata(f870_wdata), .clk(f870_clk), .rst(f870_rst), .rdata(f870_rdata));
  assign f870_clk = clk;
  assign f870_rst = rst;
  // Bindings to f870

  // f872
  logic [0:0] f872_wen;
  logic [31:0] f872_wdata;
  logic [0:0] f872_clk;
  logic [0:0] f872_rst;
  logic [31:0] f872_rdata;
  sr_buffer_32_1 f872(.wen(f872_wen), .wdata(f872_wdata), .clk(f872_clk), .rst(f872_rst), .rdata(f872_rdata));
  assign f872_clk = clk;
  assign f872_rst = rst;
  // Bindings to f872

  // f874
  logic [0:0] f874_wen;
  logic [31:0] f874_wdata;
  logic [0:0] f874_clk;
  logic [0:0] f874_rst;
  logic [31:0] f874_rdata;
  sr_buffer_32_1 f874(.wen(f874_wen), .wdata(f874_wdata), .clk(f874_clk), .rst(f874_rst), .rdata(f874_rdata));
  assign f874_clk = clk;
  assign f874_rst = rst;
  // Bindings to f874

  // f876
  logic [0:0] f876_wen;
  logic [31:0] f876_wdata;
  logic [0:0] f876_clk;
  logic [0:0] f876_rst;
  logic [31:0] f876_rdata;
  sr_buffer_32_1 f876(.wen(f876_wen), .wdata(f876_wdata), .clk(f876_clk), .rst(f876_rst), .rdata(f876_rdata));
  assign f876_clk = clk;
  assign f876_rst = rst;
  // Bindings to f876

  // f878
  logic [0:0] f878_wen;
  logic [31:0] f878_wdata;
  logic [0:0] f878_clk;
  logic [0:0] f878_rst;
  logic [31:0] f878_rdata;
  sr_buffer_32_1 f878(.wen(f878_wen), .wdata(f878_wdata), .clk(f878_clk), .rst(f878_rst), .rdata(f878_rdata));
  assign f878_clk = clk;
  assign f878_rst = rst;
  // Bindings to f878

  // f880
  logic [0:0] f880_wen;
  logic [31:0] f880_wdata;
  logic [0:0] f880_clk;
  logic [0:0] f880_rst;
  logic [31:0] f880_rdata;
  sr_buffer_32_1 f880(.wen(f880_wen), .wdata(f880_wdata), .clk(f880_clk), .rst(f880_rst), .rdata(f880_rdata));
  assign f880_clk = clk;
  assign f880_rst = rst;
  // Bindings to f880

  // f882
  logic [0:0] f882_wen;
  logic [31:0] f882_wdata;
  logic [0:0] f882_clk;
  logic [0:0] f882_rst;
  logic [31:0] f882_rdata;
  sr_buffer_32_1 f882(.wen(f882_wen), .wdata(f882_wdata), .clk(f882_clk), .rst(f882_rst), .rdata(f882_rdata));
  assign f882_clk = clk;
  assign f882_rst = rst;
  // Bindings to f882

  // f884
  logic [0:0] f884_wen;
  logic [31:0] f884_wdata;
  logic [0:0] f884_clk;
  logic [0:0] f884_rst;
  logic [31:0] f884_rdata;
  sr_buffer_32_1 f884(.wen(f884_wen), .wdata(f884_wdata), .clk(f884_clk), .rst(f884_rst), .rdata(f884_rdata));
  assign f884_clk = clk;
  assign f884_rst = rst;
  // Bindings to f884

  // f886
  logic [0:0] f886_wen;
  logic [31:0] f886_wdata;
  logic [0:0] f886_clk;
  logic [0:0] f886_rst;
  logic [31:0] f886_rdata;
  sr_buffer_32_1 f886(.wen(f886_wen), .wdata(f886_wdata), .clk(f886_clk), .rst(f886_rst), .rdata(f886_rdata));
  assign f886_clk = clk;
  assign f886_rst = rst;
  // Bindings to f886

  // f888
  logic [0:0] f888_wen;
  logic [31:0] f888_wdata;
  logic [0:0] f888_clk;
  logic [0:0] f888_rst;
  logic [31:0] f888_rdata;
  sr_buffer_32_1 f888(.wen(f888_wen), .wdata(f888_wdata), .clk(f888_clk), .rst(f888_rst), .rdata(f888_rdata));
  assign f888_clk = clk;
  assign f888_rst = rst;
  // Bindings to f888

  // f890
  logic [0:0] f890_wen;
  logic [31:0] f890_wdata;
  logic [0:0] f890_clk;
  logic [0:0] f890_rst;
  logic [31:0] f890_rdata;
  sr_buffer_32_1 f890(.wen(f890_wen), .wdata(f890_wdata), .clk(f890_clk), .rst(f890_rst), .rdata(f890_rdata));
  assign f890_clk = clk;
  assign f890_rst = rst;
  // Bindings to f890

  // f892
  logic [0:0] f892_wen;
  logic [31:0] f892_wdata;
  logic [0:0] f892_clk;
  logic [0:0] f892_rst;
  logic [31:0] f892_rdata;
  sr_buffer_32_1 f892(.wen(f892_wen), .wdata(f892_wdata), .clk(f892_clk), .rst(f892_rst), .rdata(f892_rdata));
  assign f892_clk = clk;
  assign f892_rst = rst;
  // Bindings to f892

  // f894
  logic [0:0] f894_wen;
  logic [31:0] f894_wdata;
  logic [0:0] f894_clk;
  logic [0:0] f894_rst;
  logic [31:0] f894_rdata;
  sr_buffer_32_1 f894(.wen(f894_wen), .wdata(f894_wdata), .clk(f894_clk), .rst(f894_rst), .rdata(f894_rdata));
  assign f894_clk = clk;
  assign f894_rst = rst;
  // Bindings to f894

  // f896
  logic [0:0] f896_wen;
  logic [31:0] f896_wdata;
  logic [0:0] f896_clk;
  logic [0:0] f896_rst;
  logic [31:0] f896_rdata;
  sr_buffer_32_1 f896(.wen(f896_wen), .wdata(f896_wdata), .clk(f896_clk), .rst(f896_rst), .rdata(f896_rdata));
  assign f896_clk = clk;
  assign f896_rst = rst;
  // Bindings to f896

  // f898
  logic [0:0] f898_wen;
  logic [31:0] f898_wdata;
  logic [0:0] f898_clk;
  logic [0:0] f898_rst;
  logic [31:0] f898_rdata;
  sr_buffer_32_1 f898(.wen(f898_wen), .wdata(f898_wdata), .clk(f898_clk), .rst(f898_rst), .rdata(f898_rdata));
  assign f898_clk = clk;
  assign f898_rst = rst;
  // Bindings to f898

  // f900
  logic [0:0] f900_wen;
  logic [31:0] f900_wdata;
  logic [0:0] f900_clk;
  logic [0:0] f900_rst;
  logic [31:0] f900_rdata;
  sr_buffer_32_1 f900(.wen(f900_wen), .wdata(f900_wdata), .clk(f900_clk), .rst(f900_rst), .rdata(f900_rdata));
  assign f900_clk = clk;
  assign f900_rst = rst;
  // Bindings to f900

  // f902
  logic [0:0] f902_wen;
  logic [31:0] f902_wdata;
  logic [0:0] f902_clk;
  logic [0:0] f902_rst;
  logic [31:0] f902_rdata;
  sr_buffer_32_1 f902(.wen(f902_wen), .wdata(f902_wdata), .clk(f902_clk), .rst(f902_rst), .rdata(f902_rdata));
  assign f902_clk = clk;
  assign f902_rst = rst;
  // Bindings to f902

  // f904
  logic [0:0] f904_wen;
  logic [31:0] f904_wdata;
  logic [0:0] f904_clk;
  logic [0:0] f904_rst;
  logic [31:0] f904_rdata;
  sr_buffer_32_1 f904(.wen(f904_wen), .wdata(f904_wdata), .clk(f904_clk), .rst(f904_rst), .rdata(f904_rdata));
  assign f904_clk = clk;
  assign f904_rst = rst;
  // Bindings to f904

  // f906
  logic [0:0] f906_wen;
  logic [31:0] f906_wdata;
  logic [0:0] f906_clk;
  logic [0:0] f906_rst;
  logic [31:0] f906_rdata;
  sr_buffer_32_1 f906(.wen(f906_wen), .wdata(f906_wdata), .clk(f906_clk), .rst(f906_rst), .rdata(f906_rdata));
  assign f906_clk = clk;
  assign f906_rst = rst;
  // Bindings to f906

  // f908
  logic [0:0] f908_wen;
  logic [31:0] f908_wdata;
  logic [0:0] f908_clk;
  logic [0:0] f908_rst;
  logic [31:0] f908_rdata;
  sr_buffer_32_1 f908(.wen(f908_wen), .wdata(f908_wdata), .clk(f908_clk), .rst(f908_rst), .rdata(f908_rdata));
  assign f908_clk = clk;
  assign f908_rst = rst;
  // Bindings to f908

  // f910
  logic [0:0] f910_wen;
  logic [31:0] f910_wdata;
  logic [0:0] f910_clk;
  logic [0:0] f910_rst;
  logic [31:0] f910_rdata;
  sr_buffer_32_1 f910(.wen(f910_wen), .wdata(f910_wdata), .clk(f910_clk), .rst(f910_rst), .rdata(f910_rdata));
  assign f910_clk = clk;
  assign f910_rst = rst;
  // Bindings to f910

  // f912
  logic [0:0] f912_wen;
  logic [31:0] f912_wdata;
  logic [0:0] f912_clk;
  logic [0:0] f912_rst;
  logic [31:0] f912_rdata;
  sr_buffer_32_1 f912(.wen(f912_wen), .wdata(f912_wdata), .clk(f912_clk), .rst(f912_rst), .rdata(f912_rdata));
  assign f912_clk = clk;
  assign f912_rst = rst;
  // Bindings to f912

  // f914
  logic [0:0] f914_wen;
  logic [31:0] f914_wdata;
  logic [0:0] f914_clk;
  logic [0:0] f914_rst;
  logic [31:0] f914_rdata;
  sr_buffer_32_1 f914(.wen(f914_wen), .wdata(f914_wdata), .clk(f914_clk), .rst(f914_rst), .rdata(f914_rdata));
  assign f914_clk = clk;
  assign f914_rst = rst;
  // Bindings to f914

  // f916
  logic [0:0] f916_wen;
  logic [31:0] f916_wdata;
  logic [0:0] f916_clk;
  logic [0:0] f916_rst;
  logic [31:0] f916_rdata;
  sr_buffer_32_1 f916(.wen(f916_wen), .wdata(f916_wdata), .clk(f916_clk), .rst(f916_rst), .rdata(f916_rdata));
  assign f916_clk = clk;
  assign f916_rst = rst;
  // Bindings to f916

  // f918
  logic [0:0] f918_wen;
  logic [31:0] f918_wdata;
  logic [0:0] f918_clk;
  logic [0:0] f918_rst;
  logic [31:0] f918_rdata;
  sr_buffer_32_1 f918(.wen(f918_wen), .wdata(f918_wdata), .clk(f918_clk), .rst(f918_rst), .rdata(f918_rdata));
  assign f918_clk = clk;
  assign f918_rst = rst;
  // Bindings to f918

  // f920
  logic [0:0] f920_wen;
  logic [31:0] f920_wdata;
  logic [0:0] f920_clk;
  logic [0:0] f920_rst;
  logic [31:0] f920_rdata;
  sr_buffer_32_1 f920(.wen(f920_wen), .wdata(f920_wdata), .clk(f920_clk), .rst(f920_rst), .rdata(f920_rdata));
  assign f920_clk = clk;
  assign f920_rst = rst;
  // Bindings to f920

  // f922
  logic [0:0] f922_wen;
  logic [31:0] f922_wdata;
  logic [0:0] f922_clk;
  logic [0:0] f922_rst;
  logic [31:0] f922_rdata;
  sr_buffer_32_1 f922(.wen(f922_wen), .wdata(f922_wdata), .clk(f922_clk), .rst(f922_rst), .rdata(f922_rdata));
  assign f922_clk = clk;
  assign f922_rst = rst;
  // Bindings to f922

  // f924
  logic [0:0] f924_wen;
  logic [31:0] f924_wdata;
  logic [0:0] f924_clk;
  logic [0:0] f924_rst;
  logic [31:0] f924_rdata;
  sr_buffer_32_1 f924(.wen(f924_wen), .wdata(f924_wdata), .clk(f924_clk), .rst(f924_rst), .rdata(f924_rdata));
  assign f924_clk = clk;
  assign f924_rst = rst;
  // Bindings to f924

  // f926
  logic [0:0] f926_wen;
  logic [31:0] f926_wdata;
  logic [0:0] f926_clk;
  logic [0:0] f926_rst;
  logic [31:0] f926_rdata;
  sr_buffer_32_1 f926(.wen(f926_wen), .wdata(f926_wdata), .clk(f926_clk), .rst(f926_rst), .rdata(f926_rdata));
  assign f926_clk = clk;
  assign f926_rst = rst;
  // Bindings to f926

  // f928
  logic [0:0] f928_wen;
  logic [31:0] f928_wdata;
  logic [0:0] f928_clk;
  logic [0:0] f928_rst;
  logic [31:0] f928_rdata;
  sr_buffer_32_1 f928(.wen(f928_wen), .wdata(f928_wdata), .clk(f928_clk), .rst(f928_rst), .rdata(f928_rdata));
  assign f928_clk = clk;
  assign f928_rst = rst;
  // Bindings to f928

  // f930
  logic [0:0] f930_wen;
  logic [31:0] f930_wdata;
  logic [0:0] f930_clk;
  logic [0:0] f930_rst;
  logic [31:0] f930_rdata;
  sr_buffer_32_1 f930(.wen(f930_wen), .wdata(f930_wdata), .clk(f930_clk), .rst(f930_rst), .rdata(f930_rdata));
  assign f930_clk = clk;
  assign f930_rst = rst;
  // Bindings to f930

  // f932
  logic [0:0] f932_wen;
  logic [31:0] f932_wdata;
  logic [0:0] f932_clk;
  logic [0:0] f932_rst;
  logic [31:0] f932_rdata;
  sr_buffer_32_1 f932(.wen(f932_wen), .wdata(f932_wdata), .clk(f932_clk), .rst(f932_rst), .rdata(f932_rdata));
  assign f932_clk = clk;
  assign f932_rst = rst;
  // Bindings to f932

  // f934
  logic [0:0] f934_wen;
  logic [31:0] f934_wdata;
  logic [0:0] f934_clk;
  logic [0:0] f934_rst;
  logic [31:0] f934_rdata;
  sr_buffer_32_1 f934(.wen(f934_wen), .wdata(f934_wdata), .clk(f934_clk), .rst(f934_rst), .rdata(f934_rdata));
  assign f934_clk = clk;
  assign f934_rst = rst;
  // Bindings to f934

  // f936
  logic [0:0] f936_wen;
  logic [31:0] f936_wdata;
  logic [0:0] f936_clk;
  logic [0:0] f936_rst;
  logic [31:0] f936_rdata;
  sr_buffer_32_1 f936(.wen(f936_wen), .wdata(f936_wdata), .clk(f936_clk), .rst(f936_rst), .rdata(f936_rdata));
  assign f936_clk = clk;
  assign f936_rst = rst;
  // Bindings to f936

  // f938
  logic [0:0] f938_wen;
  logic [31:0] f938_wdata;
  logic [0:0] f938_clk;
  logic [0:0] f938_rst;
  logic [31:0] f938_rdata;
  sr_buffer_32_1 f938(.wen(f938_wen), .wdata(f938_wdata), .clk(f938_clk), .rst(f938_rst), .rdata(f938_rdata));
  assign f938_clk = clk;
  assign f938_rst = rst;
  // Bindings to f938

  // f940
  logic [0:0] f940_wen;
  logic [31:0] f940_wdata;
  logic [0:0] f940_clk;
  logic [0:0] f940_rst;
  logic [31:0] f940_rdata;
  sr_buffer_32_1 f940(.wen(f940_wen), .wdata(f940_wdata), .clk(f940_clk), .rst(f940_rst), .rdata(f940_rdata));
  assign f940_clk = clk;
  assign f940_rst = rst;
  // Bindings to f940

  // f942
  logic [0:0] f942_wen;
  logic [31:0] f942_wdata;
  logic [0:0] f942_clk;
  logic [0:0] f942_rst;
  logic [31:0] f942_rdata;
  sr_buffer_32_1 f942(.wen(f942_wen), .wdata(f942_wdata), .clk(f942_clk), .rst(f942_rst), .rdata(f942_rdata));
  assign f942_clk = clk;
  assign f942_rst = rst;
  // Bindings to f942

  // f944
  logic [0:0] f944_wen;
  logic [31:0] f944_wdata;
  logic [0:0] f944_clk;
  logic [0:0] f944_rst;
  logic [31:0] f944_rdata;
  sr_buffer_32_1 f944(.wen(f944_wen), .wdata(f944_wdata), .clk(f944_clk), .rst(f944_rst), .rdata(f944_rdata));
  assign f944_clk = clk;
  assign f944_rst = rst;
  // Bindings to f944

  // f946
  logic [0:0] f946_wen;
  logic [31:0] f946_wdata;
  logic [0:0] f946_clk;
  logic [0:0] f946_rst;
  logic [31:0] f946_rdata;
  sr_buffer_32_1 f946(.wen(f946_wen), .wdata(f946_wdata), .clk(f946_clk), .rst(f946_rst), .rdata(f946_rdata));
  assign f946_clk = clk;
  assign f946_rst = rst;
  // Bindings to f946

  // f948
  logic [0:0] f948_wen;
  logic [31:0] f948_wdata;
  logic [0:0] f948_clk;
  logic [0:0] f948_rst;
  logic [31:0] f948_rdata;
  sr_buffer_32_1 f948(.wen(f948_wen), .wdata(f948_wdata), .clk(f948_clk), .rst(f948_rst), .rdata(f948_rdata));
  assign f948_clk = clk;
  assign f948_rst = rst;
  // Bindings to f948

  // f950
  logic [0:0] f950_wen;
  logic [31:0] f950_wdata;
  logic [0:0] f950_clk;
  logic [0:0] f950_rst;
  logic [31:0] f950_rdata;
  sr_buffer_32_1 f950(.wen(f950_wen), .wdata(f950_wdata), .clk(f950_clk), .rst(f950_rst), .rdata(f950_rdata));
  assign f950_clk = clk;
  assign f950_rst = rst;
  // Bindings to f950

  // f952
  logic [0:0] f952_wen;
  logic [31:0] f952_wdata;
  logic [0:0] f952_clk;
  logic [0:0] f952_rst;
  logic [31:0] f952_rdata;
  sr_buffer_32_1 f952(.wen(f952_wen), .wdata(f952_wdata), .clk(f952_clk), .rst(f952_rst), .rdata(f952_rdata));
  assign f952_clk = clk;
  assign f952_rst = rst;
  // Bindings to f952

  // f954
  logic [0:0] f954_wen;
  logic [31:0] f954_wdata;
  logic [0:0] f954_clk;
  logic [0:0] f954_rst;
  logic [31:0] f954_rdata;
  sr_buffer_32_1 f954(.wen(f954_wen), .wdata(f954_wdata), .clk(f954_clk), .rst(f954_rst), .rdata(f954_rdata));
  assign f954_clk = clk;
  assign f954_rst = rst;
  // Bindings to f954

  // f956
  logic [0:0] f956_wen;
  logic [31:0] f956_wdata;
  logic [0:0] f956_clk;
  logic [0:0] f956_rst;
  logic [31:0] f956_rdata;
  sr_buffer_32_1 f956(.wen(f956_wen), .wdata(f956_wdata), .clk(f956_clk), .rst(f956_rst), .rdata(f956_rdata));
  assign f956_clk = clk;
  assign f956_rst = rst;
  // Bindings to f956

  // f958
  logic [0:0] f958_wen;
  logic [31:0] f958_wdata;
  logic [0:0] f958_clk;
  logic [0:0] f958_rst;
  logic [31:0] f958_rdata;
  sr_buffer_32_1 f958(.wen(f958_wen), .wdata(f958_wdata), .clk(f958_clk), .rst(f958_rst), .rdata(f958_rdata));
  assign f958_clk = clk;
  assign f958_rst = rst;
  // Bindings to f958

  // f960
  logic [0:0] f960_wen;
  logic [31:0] f960_wdata;
  logic [0:0] f960_clk;
  logic [0:0] f960_rst;
  logic [31:0] f960_rdata;
  sr_buffer_32_1 f960(.wen(f960_wen), .wdata(f960_wdata), .clk(f960_clk), .rst(f960_rst), .rdata(f960_rdata));
  assign f960_clk = clk;
  assign f960_rst = rst;
  // Bindings to f960

  // f962
  logic [0:0] f962_wen;
  logic [31:0] f962_wdata;
  logic [0:0] f962_clk;
  logic [0:0] f962_rst;
  logic [31:0] f962_rdata;
  sr_buffer_32_1 f962(.wen(f962_wen), .wdata(f962_wdata), .clk(f962_clk), .rst(f962_rst), .rdata(f962_rdata));
  assign f962_clk = clk;
  assign f962_rst = rst;
  // Bindings to f962

  // f964
  logic [0:0] f964_wen;
  logic [31:0] f964_wdata;
  logic [0:0] f964_clk;
  logic [0:0] f964_rst;
  logic [31:0] f964_rdata;
  sr_buffer_32_1 f964(.wen(f964_wen), .wdata(f964_wdata), .clk(f964_clk), .rst(f964_rst), .rdata(f964_rdata));
  assign f964_clk = clk;
  assign f964_rst = rst;
  // Bindings to f964

  // f966
  logic [0:0] f966_wen;
  logic [31:0] f966_wdata;
  logic [0:0] f966_clk;
  logic [0:0] f966_rst;
  logic [31:0] f966_rdata;
  sr_buffer_32_1 f966(.wen(f966_wen), .wdata(f966_wdata), .clk(f966_clk), .rst(f966_rst), .rdata(f966_rdata));
  assign f966_clk = clk;
  assign f966_rst = rst;
  // Bindings to f966

  // f968
  logic [0:0] f968_wen;
  logic [31:0] f968_wdata;
  logic [0:0] f968_clk;
  logic [0:0] f968_rst;
  logic [31:0] f968_rdata;
  sr_buffer_32_1 f968(.wen(f968_wen), .wdata(f968_wdata), .clk(f968_clk), .rst(f968_rst), .rdata(f968_rdata));
  assign f968_clk = clk;
  assign f968_rst = rst;
  // Bindings to f968

  // f970
  logic [0:0] f970_wen;
  logic [31:0] f970_wdata;
  logic [0:0] f970_clk;
  logic [0:0] f970_rst;
  logic [31:0] f970_rdata;
  sr_buffer_32_1 f970(.wen(f970_wen), .wdata(f970_wdata), .clk(f970_clk), .rst(f970_rst), .rdata(f970_rdata));
  assign f970_clk = clk;
  assign f970_rst = rst;
  // Bindings to f970

  // f972
  logic [0:0] f972_wen;
  logic [31:0] f972_wdata;
  logic [0:0] f972_clk;
  logic [0:0] f972_rst;
  logic [31:0] f972_rdata;
  sr_buffer_32_1 f972(.wen(f972_wen), .wdata(f972_wdata), .clk(f972_clk), .rst(f972_rst), .rdata(f972_rdata));
  assign f972_clk = clk;
  assign f972_rst = rst;
  // Bindings to f972

  // f974
  logic [0:0] f974_wen;
  logic [31:0] f974_wdata;
  logic [0:0] f974_clk;
  logic [0:0] f974_rst;
  logic [31:0] f974_rdata;
  sr_buffer_32_1 f974(.wen(f974_wen), .wdata(f974_wdata), .clk(f974_clk), .rst(f974_rst), .rdata(f974_rdata));
  assign f974_clk = clk;
  assign f974_rst = rst;
  // Bindings to f974

  // f976
  logic [0:0] f976_wen;
  logic [31:0] f976_wdata;
  logic [0:0] f976_clk;
  logic [0:0] f976_rst;
  logic [31:0] f976_rdata;
  sr_buffer_32_1 f976(.wen(f976_wen), .wdata(f976_wdata), .clk(f976_clk), .rst(f976_rst), .rdata(f976_rdata));
  assign f976_clk = clk;
  assign f976_rst = rst;
  // Bindings to f976

  // f978
  logic [0:0] f978_wen;
  logic [31:0] f978_wdata;
  logic [0:0] f978_clk;
  logic [0:0] f978_rst;
  logic [31:0] f978_rdata;
  sr_buffer_32_1 f978(.wen(f978_wen), .wdata(f978_wdata), .clk(f978_clk), .rst(f978_rst), .rdata(f978_rdata));
  assign f978_clk = clk;
  assign f978_rst = rst;
  // Bindings to f978

  // f980
  logic [0:0] f980_wen;
  logic [31:0] f980_wdata;
  logic [0:0] f980_clk;
  logic [0:0] f980_rst;
  logic [31:0] f980_rdata;
  sr_buffer_32_1 f980(.wen(f980_wen), .wdata(f980_wdata), .clk(f980_clk), .rst(f980_rst), .rdata(f980_rdata));
  assign f980_clk = clk;
  assign f980_rst = rst;
  // Bindings to f980

  // f982
  logic [0:0] f982_wen;
  logic [31:0] f982_wdata;
  logic [0:0] f982_clk;
  logic [0:0] f982_rst;
  logic [31:0] f982_rdata;
  sr_buffer_32_1 f982(.wen(f982_wen), .wdata(f982_wdata), .clk(f982_clk), .rst(f982_rst), .rdata(f982_rdata));
  assign f982_clk = clk;
  assign f982_rst = rst;
  // Bindings to f982

  // f984
  logic [0:0] f984_wen;
  logic [31:0] f984_wdata;
  logic [0:0] f984_clk;
  logic [0:0] f984_rst;
  logic [31:0] f984_rdata;
  sr_buffer_32_1 f984(.wen(f984_wen), .wdata(f984_wdata), .clk(f984_clk), .rst(f984_rst), .rdata(f984_rdata));
  assign f984_clk = clk;
  assign f984_rst = rst;
  // Bindings to f984

  // f986
  logic [0:0] f986_wen;
  logic [31:0] f986_wdata;
  logic [0:0] f986_clk;
  logic [0:0] f986_rst;
  logic [31:0] f986_rdata;
  sr_buffer_32_1 f986(.wen(f986_wen), .wdata(f986_wdata), .clk(f986_clk), .rst(f986_rst), .rdata(f986_rdata));
  assign f986_clk = clk;
  assign f986_rst = rst;
  // Bindings to f986

  // f988
  logic [0:0] f988_wen;
  logic [31:0] f988_wdata;
  logic [0:0] f988_clk;
  logic [0:0] f988_rst;
  logic [31:0] f988_rdata;
  sr_buffer_32_1 f988(.wen(f988_wen), .wdata(f988_wdata), .clk(f988_clk), .rst(f988_rst), .rdata(f988_rdata));
  assign f988_clk = clk;
  assign f988_rst = rst;
  // Bindings to f988

  // f990
  logic [0:0] f990_wen;
  logic [31:0] f990_wdata;
  logic [0:0] f990_clk;
  logic [0:0] f990_rst;
  logic [31:0] f990_rdata;
  sr_buffer_32_1 f990(.wen(f990_wen), .wdata(f990_wdata), .clk(f990_clk), .rst(f990_rst), .rdata(f990_rdata));
  assign f990_clk = clk;
  assign f990_rst = rst;
  // Bindings to f990

  // f992
  logic [0:0] f992_wen;
  logic [31:0] f992_wdata;
  logic [0:0] f992_clk;
  logic [0:0] f992_rst;
  logic [31:0] f992_rdata;
  sr_buffer_32_1 f992(.wen(f992_wen), .wdata(f992_wdata), .clk(f992_clk), .rst(f992_rst), .rdata(f992_rdata));
  assign f992_clk = clk;
  assign f992_rst = rst;
  // Bindings to f992

  // f994
  logic [0:0] f994_wen;
  logic [31:0] f994_wdata;
  logic [0:0] f994_clk;
  logic [0:0] f994_rst;
  logic [31:0] f994_rdata;
  sr_buffer_32_1 f994(.wen(f994_wen), .wdata(f994_wdata), .clk(f994_clk), .rst(f994_rst), .rdata(f994_rdata));
  assign f994_clk = clk;
  assign f994_rst = rst;
  // Bindings to f994

  // f996
  logic [0:0] f996_wen;
  logic [31:0] f996_wdata;
  logic [0:0] f996_clk;
  logic [0:0] f996_rst;
  logic [31:0] f996_rdata;
  sr_buffer_32_1 f996(.wen(f996_wen), .wdata(f996_wdata), .clk(f996_clk), .rst(f996_rst), .rdata(f996_rdata));
  assign f996_clk = clk;
  assign f996_rst = rst;
  // Bindings to f996

  // f998
  logic [0:0] f998_wen;
  logic [31:0] f998_wdata;
  logic [0:0] f998_clk;
  logic [0:0] f998_rst;
  logic [31:0] f998_rdata;
  sr_buffer_32_1 f998(.wen(f998_wen), .wdata(f998_wdata), .clk(f998_clk), .rst(f998_rst), .rdata(f998_rdata));
  assign f998_clk = clk;
  assign f998_rst = rst;
  // Bindings to f998

  // f1000
  logic [0:0] f1000_wen;
  logic [31:0] f1000_wdata;
  logic [0:0] f1000_clk;
  logic [0:0] f1000_rst;
  logic [31:0] f1000_rdata;
  sr_buffer_32_1 f1000(.wen(f1000_wen), .wdata(f1000_wdata), .clk(f1000_clk), .rst(f1000_rst), .rdata(f1000_rdata));
  assign f1000_clk = clk;
  assign f1000_rst = rst;
  // Bindings to f1000

  // f1002
  logic [0:0] f1002_wen;
  logic [31:0] f1002_wdata;
  logic [0:0] f1002_clk;
  logic [0:0] f1002_rst;
  logic [31:0] f1002_rdata;
  sr_buffer_32_1 f1002(.wen(f1002_wen), .wdata(f1002_wdata), .clk(f1002_clk), .rst(f1002_rst), .rdata(f1002_rdata));
  assign f1002_clk = clk;
  assign f1002_rst = rst;
  // Bindings to f1002

  // f1004
  logic [0:0] f1004_wen;
  logic [31:0] f1004_wdata;
  logic [0:0] f1004_clk;
  logic [0:0] f1004_rst;
  logic [31:0] f1004_rdata;
  sr_buffer_32_1 f1004(.wen(f1004_wen), .wdata(f1004_wdata), .clk(f1004_clk), .rst(f1004_rst), .rdata(f1004_rdata));
  assign f1004_clk = clk;
  assign f1004_rst = rst;
  // Bindings to f1004

  // f1006
  logic [0:0] f1006_wen;
  logic [31:0] f1006_wdata;
  logic [0:0] f1006_clk;
  logic [0:0] f1006_rst;
  logic [31:0] f1006_rdata;
  sr_buffer_32_1 f1006(.wen(f1006_wen), .wdata(f1006_wdata), .clk(f1006_clk), .rst(f1006_rst), .rdata(f1006_rdata));
  assign f1006_clk = clk;
  assign f1006_rst = rst;
  // Bindings to f1006

  // f1008
  logic [0:0] f1008_wen;
  logic [31:0] f1008_wdata;
  logic [0:0] f1008_clk;
  logic [0:0] f1008_rst;
  logic [31:0] f1008_rdata;
  sr_buffer_32_1 f1008(.wen(f1008_wen), .wdata(f1008_wdata), .clk(f1008_clk), .rst(f1008_rst), .rdata(f1008_rdata));
  assign f1008_clk = clk;
  assign f1008_rst = rst;
  // Bindings to f1008

  // f1010
  logic [0:0] f1010_wen;
  logic [31:0] f1010_wdata;
  logic [0:0] f1010_clk;
  logic [0:0] f1010_rst;
  logic [31:0] f1010_rdata;
  sr_buffer_32_1 f1010(.wen(f1010_wen), .wdata(f1010_wdata), .clk(f1010_clk), .rst(f1010_rst), .rdata(f1010_rdata));
  assign f1010_clk = clk;
  assign f1010_rst = rst;
  // Bindings to f1010

  // f1012
  logic [0:0] f1012_wen;
  logic [31:0] f1012_wdata;
  logic [0:0] f1012_clk;
  logic [0:0] f1012_rst;
  logic [31:0] f1012_rdata;
  sr_buffer_32_1 f1012(.wen(f1012_wen), .wdata(f1012_wdata), .clk(f1012_clk), .rst(f1012_rst), .rdata(f1012_rdata));
  assign f1012_clk = clk;
  assign f1012_rst = rst;
  // Bindings to f1012

  // f1014
  logic [0:0] f1014_wen;
  logic [31:0] f1014_wdata;
  logic [0:0] f1014_clk;
  logic [0:0] f1014_rst;
  logic [31:0] f1014_rdata;
  sr_buffer_32_1 f1014(.wen(f1014_wen), .wdata(f1014_wdata), .clk(f1014_clk), .rst(f1014_rst), .rdata(f1014_rdata));
  assign f1014_clk = clk;
  assign f1014_rst = rst;
  // Bindings to f1014

  // f1016
  logic [0:0] f1016_wen;
  logic [31:0] f1016_wdata;
  logic [0:0] f1016_clk;
  logic [0:0] f1016_rst;
  logic [31:0] f1016_rdata;
  sr_buffer_32_1 f1016(.wen(f1016_wen), .wdata(f1016_wdata), .clk(f1016_clk), .rst(f1016_rst), .rdata(f1016_rdata));
  assign f1016_clk = clk;
  assign f1016_rst = rst;
  // Bindings to f1016

  // f1018
  logic [0:0] f1018_wen;
  logic [31:0] f1018_wdata;
  logic [0:0] f1018_clk;
  logic [0:0] f1018_rst;
  logic [31:0] f1018_rdata;
  sr_buffer_32_1 f1018(.wen(f1018_wen), .wdata(f1018_wdata), .clk(f1018_clk), .rst(f1018_rst), .rdata(f1018_rdata));
  assign f1018_clk = clk;
  assign f1018_rst = rst;
  // Bindings to f1018

  // f1020
  logic [0:0] f1020_wen;
  logic [31:0] f1020_wdata;
  logic [0:0] f1020_clk;
  logic [0:0] f1020_rst;
  logic [31:0] f1020_rdata;
  sr_buffer_32_1 f1020(.wen(f1020_wen), .wdata(f1020_wdata), .clk(f1020_clk), .rst(f1020_rst), .rdata(f1020_rdata));
  assign f1020_clk = clk;
  assign f1020_rst = rst;
  // Bindings to f1020

  // f1022
  logic [0:0] f1022_wen;
  logic [31:0] f1022_wdata;
  logic [0:0] f1022_clk;
  logic [0:0] f1022_rst;
  logic [31:0] f1022_rdata;
  sr_buffer_32_1 f1022(.wen(f1022_wen), .wdata(f1022_wdata), .clk(f1022_clk), .rst(f1022_rst), .rdata(f1022_rdata));
  assign f1022_clk = clk;
  assign f1022_rst = rst;
  // Bindings to f1022

  // f1024
  logic [0:0] f1024_wen;
  logic [31:0] f1024_wdata;
  logic [0:0] f1024_clk;
  logic [0:0] f1024_rst;
  logic [31:0] f1024_rdata;
  sr_buffer_32_1 f1024(.wen(f1024_wen), .wdata(f1024_wdata), .clk(f1024_clk), .rst(f1024_rst), .rdata(f1024_rdata));
  assign f1024_clk = clk;
  assign f1024_rst = rst;
  // Bindings to f1024

  // f1026
  logic [0:0] f1026_wen;
  logic [31:0] f1026_wdata;
  logic [0:0] f1026_clk;
  logic [0:0] f1026_rst;
  logic [31:0] f1026_rdata;
  sr_buffer_32_1 f1026(.wen(f1026_wen), .wdata(f1026_wdata), .clk(f1026_clk), .rst(f1026_rst), .rdata(f1026_rdata));
  assign f1026_clk = clk;
  assign f1026_rst = rst;
  // Bindings to f1026

  // f1028
  logic [0:0] f1028_wen;
  logic [31:0] f1028_wdata;
  logic [0:0] f1028_clk;
  logic [0:0] f1028_rst;
  logic [31:0] f1028_rdata;
  sr_buffer_32_1 f1028(.wen(f1028_wen), .wdata(f1028_wdata), .clk(f1028_clk), .rst(f1028_rst), .rdata(f1028_rdata));
  assign f1028_clk = clk;
  assign f1028_rst = rst;
  // Bindings to f1028

  // f1030
  logic [0:0] f1030_wen;
  logic [31:0] f1030_wdata;
  logic [0:0] f1030_clk;
  logic [0:0] f1030_rst;
  logic [31:0] f1030_rdata;
  sr_buffer_32_1 f1030(.wen(f1030_wen), .wdata(f1030_wdata), .clk(f1030_clk), .rst(f1030_rst), .rdata(f1030_rdata));
  assign f1030_clk = clk;
  assign f1030_rst = rst;
  // Bindings to f1030

  // f1032
  logic [0:0] f1032_wen;
  logic [31:0] f1032_wdata;
  logic [0:0] f1032_clk;
  logic [0:0] f1032_rst;
  logic [31:0] f1032_rdata;
  sr_buffer_32_1 f1032(.wen(f1032_wen), .wdata(f1032_wdata), .clk(f1032_clk), .rst(f1032_rst), .rdata(f1032_rdata));
  assign f1032_clk = clk;
  assign f1032_rst = rst;
  // Bindings to f1032

  // f1034
  logic [0:0] f1034_wen;
  logic [31:0] f1034_wdata;
  logic [0:0] f1034_clk;
  logic [0:0] f1034_rst;
  logic [31:0] f1034_rdata;
  sr_buffer_32_1 f1034(.wen(f1034_wen), .wdata(f1034_wdata), .clk(f1034_clk), .rst(f1034_rst), .rdata(f1034_rdata));
  assign f1034_clk = clk;
  assign f1034_rst = rst;
  // Bindings to f1034

  // f1036
  logic [0:0] f1036_wen;
  logic [31:0] f1036_wdata;
  logic [0:0] f1036_clk;
  logic [0:0] f1036_rst;
  logic [31:0] f1036_rdata;
  sr_buffer_32_1 f1036(.wen(f1036_wen), .wdata(f1036_wdata), .clk(f1036_clk), .rst(f1036_rst), .rdata(f1036_rdata));
  assign f1036_clk = clk;
  assign f1036_rst = rst;
  // Bindings to f1036

  // f1038
  logic [0:0] f1038_wen;
  logic [31:0] f1038_wdata;
  logic [0:0] f1038_clk;
  logic [0:0] f1038_rst;
  logic [31:0] f1038_rdata;
  sr_buffer_32_1 f1038(.wen(f1038_wen), .wdata(f1038_wdata), .clk(f1038_clk), .rst(f1038_rst), .rdata(f1038_rdata));
  assign f1038_clk = clk;
  assign f1038_rst = rst;
  // Bindings to f1038

  // f1040
  logic [0:0] f1040_wen;
  logic [31:0] f1040_wdata;
  logic [0:0] f1040_clk;
  logic [0:0] f1040_rst;
  logic [31:0] f1040_rdata;
  sr_buffer_32_1 f1040(.wen(f1040_wen), .wdata(f1040_wdata), .clk(f1040_clk), .rst(f1040_rst), .rdata(f1040_rdata));
  assign f1040_clk = clk;
  assign f1040_rst = rst;
  // Bindings to f1040

  // f1042
  logic [0:0] f1042_wen;
  logic [31:0] f1042_wdata;
  logic [0:0] f1042_clk;
  logic [0:0] f1042_rst;
  logic [31:0] f1042_rdata;
  sr_buffer_32_1 f1042(.wen(f1042_wen), .wdata(f1042_wdata), .clk(f1042_clk), .rst(f1042_rst), .rdata(f1042_rdata));
  assign f1042_clk = clk;
  assign f1042_rst = rst;
  // Bindings to f1042

  // f1044
  logic [0:0] f1044_wen;
  logic [31:0] f1044_wdata;
  logic [0:0] f1044_clk;
  logic [0:0] f1044_rst;
  logic [31:0] f1044_rdata;
  sr_buffer_32_1 f1044(.wen(f1044_wen), .wdata(f1044_wdata), .clk(f1044_clk), .rst(f1044_rst), .rdata(f1044_rdata));
  assign f1044_clk = clk;
  assign f1044_rst = rst;
  // Bindings to f1044

  // f1046
  logic [0:0] f1046_wen;
  logic [31:0] f1046_wdata;
  logic [0:0] f1046_clk;
  logic [0:0] f1046_rst;
  logic [31:0] f1046_rdata;
  sr_buffer_32_1 f1046(.wen(f1046_wen), .wdata(f1046_wdata), .clk(f1046_clk), .rst(f1046_rst), .rdata(f1046_rdata));
  assign f1046_clk = clk;
  assign f1046_rst = rst;
  // Bindings to f1046

  // f1048
  logic [0:0] f1048_wen;
  logic [31:0] f1048_wdata;
  logic [0:0] f1048_clk;
  logic [0:0] f1048_rst;
  logic [31:0] f1048_rdata;
  sr_buffer_32_1 f1048(.wen(f1048_wen), .wdata(f1048_wdata), .clk(f1048_clk), .rst(f1048_rst), .rdata(f1048_rdata));
  assign f1048_clk = clk;
  assign f1048_rst = rst;
  // Bindings to f1048

  // f1050
  logic [0:0] f1050_wen;
  logic [31:0] f1050_wdata;
  logic [0:0] f1050_clk;
  logic [0:0] f1050_rst;
  logic [31:0] f1050_rdata;
  sr_buffer_32_1 f1050(.wen(f1050_wen), .wdata(f1050_wdata), .clk(f1050_clk), .rst(f1050_rst), .rdata(f1050_rdata));
  assign f1050_clk = clk;
  assign f1050_rst = rst;
  // Bindings to f1050

  // f1052
  logic [0:0] f1052_wen;
  logic [31:0] f1052_wdata;
  logic [0:0] f1052_clk;
  logic [0:0] f1052_rst;
  logic [31:0] f1052_rdata;
  sr_buffer_32_1 f1052(.wen(f1052_wen), .wdata(f1052_wdata), .clk(f1052_clk), .rst(f1052_rst), .rdata(f1052_rdata));
  assign f1052_clk = clk;
  assign f1052_rst = rst;
  // Bindings to f1052

  // f1054
  logic [0:0] f1054_wen;
  logic [31:0] f1054_wdata;
  logic [0:0] f1054_clk;
  logic [0:0] f1054_rst;
  logic [31:0] f1054_rdata;
  sr_buffer_32_1 f1054(.wen(f1054_wen), .wdata(f1054_wdata), .clk(f1054_clk), .rst(f1054_rst), .rdata(f1054_rdata));
  assign f1054_clk = clk;
  assign f1054_rst = rst;
  // Bindings to f1054

  // f1056
  logic [0:0] f1056_wen;
  logic [31:0] f1056_wdata;
  logic [0:0] f1056_clk;
  logic [0:0] f1056_rst;
  logic [31:0] f1056_rdata;
  sr_buffer_32_1 f1056(.wen(f1056_wen), .wdata(f1056_wdata), .clk(f1056_clk), .rst(f1056_rst), .rdata(f1056_rdata));
  assign f1056_clk = clk;
  assign f1056_rst = rst;
  // Bindings to f1056

  // f1058
  logic [0:0] f1058_wen;
  logic [31:0] f1058_wdata;
  logic [0:0] f1058_clk;
  logic [0:0] f1058_rst;
  logic [31:0] f1058_rdata;
  sr_buffer_32_1 f1058(.wen(f1058_wen), .wdata(f1058_wdata), .clk(f1058_clk), .rst(f1058_rst), .rdata(f1058_rdata));
  assign f1058_clk = clk;
  assign f1058_rst = rst;
  // Bindings to f1058

  // f1060
  logic [0:0] f1060_wen;
  logic [31:0] f1060_wdata;
  logic [0:0] f1060_clk;
  logic [0:0] f1060_rst;
  logic [31:0] f1060_rdata;
  sr_buffer_32_1 f1060(.wen(f1060_wen), .wdata(f1060_wdata), .clk(f1060_clk), .rst(f1060_rst), .rdata(f1060_rdata));
  assign f1060_clk = clk;
  assign f1060_rst = rst;
  // Bindings to f1060

  // f1062
  logic [0:0] f1062_wen;
  logic [31:0] f1062_wdata;
  logic [0:0] f1062_clk;
  logic [0:0] f1062_rst;
  logic [31:0] f1062_rdata;
  sr_buffer_32_1 f1062(.wen(f1062_wen), .wdata(f1062_wdata), .clk(f1062_clk), .rst(f1062_rst), .rdata(f1062_rdata));
  assign f1062_clk = clk;
  assign f1062_rst = rst;
  // Bindings to f1062

  // f1064
  logic [0:0] f1064_wen;
  logic [31:0] f1064_wdata;
  logic [0:0] f1064_clk;
  logic [0:0] f1064_rst;
  logic [31:0] f1064_rdata;
  sr_buffer_32_1 f1064(.wen(f1064_wen), .wdata(f1064_wdata), .clk(f1064_clk), .rst(f1064_rst), .rdata(f1064_rdata));
  assign f1064_clk = clk;
  assign f1064_rst = rst;
  // Bindings to f1064

  // f1066
  logic [0:0] f1066_wen;
  logic [31:0] f1066_wdata;
  logic [0:0] f1066_clk;
  logic [0:0] f1066_rst;
  logic [31:0] f1066_rdata;
  sr_buffer_32_1 f1066(.wen(f1066_wen), .wdata(f1066_wdata), .clk(f1066_clk), .rst(f1066_rst), .rdata(f1066_rdata));
  assign f1066_clk = clk;
  assign f1066_rst = rst;
  // Bindings to f1066

  // f1068
  logic [0:0] f1068_wen;
  logic [31:0] f1068_wdata;
  logic [0:0] f1068_clk;
  logic [0:0] f1068_rst;
  logic [31:0] f1068_rdata;
  sr_buffer_32_1 f1068(.wen(f1068_wen), .wdata(f1068_wdata), .clk(f1068_clk), .rst(f1068_rst), .rdata(f1068_rdata));
  assign f1068_clk = clk;
  assign f1068_rst = rst;
  // Bindings to f1068

  // f1070
  logic [0:0] f1070_wen;
  logic [31:0] f1070_wdata;
  logic [0:0] f1070_clk;
  logic [0:0] f1070_rst;
  logic [31:0] f1070_rdata;
  sr_buffer_32_1 f1070(.wen(f1070_wen), .wdata(f1070_wdata), .clk(f1070_clk), .rst(f1070_rst), .rdata(f1070_rdata));
  assign f1070_clk = clk;
  assign f1070_rst = rst;
  // Bindings to f1070

  // f1072
  logic [0:0] f1072_wen;
  logic [31:0] f1072_wdata;
  logic [0:0] f1072_clk;
  logic [0:0] f1072_rst;
  logic [31:0] f1072_rdata;
  sr_buffer_32_1 f1072(.wen(f1072_wen), .wdata(f1072_wdata), .clk(f1072_clk), .rst(f1072_rst), .rdata(f1072_rdata));
  assign f1072_clk = clk;
  assign f1072_rst = rst;
  // Bindings to f1072

  // f1074
  logic [0:0] f1074_wen;
  logic [31:0] f1074_wdata;
  logic [0:0] f1074_clk;
  logic [0:0] f1074_rst;
  logic [31:0] f1074_rdata;
  sr_buffer_32_1 f1074(.wen(f1074_wen), .wdata(f1074_wdata), .clk(f1074_clk), .rst(f1074_rst), .rdata(f1074_rdata));
  assign f1074_clk = clk;
  assign f1074_rst = rst;
  // Bindings to f1074

  // f1076
  logic [0:0] f1076_wen;
  logic [31:0] f1076_wdata;
  logic [0:0] f1076_clk;
  logic [0:0] f1076_rst;
  logic [31:0] f1076_rdata;
  sr_buffer_32_1 f1076(.wen(f1076_wen), .wdata(f1076_wdata), .clk(f1076_clk), .rst(f1076_rst), .rdata(f1076_rdata));
  assign f1076_clk = clk;
  assign f1076_rst = rst;
  // Bindings to f1076

  // f1078
  logic [0:0] f1078_wen;
  logic [31:0] f1078_wdata;
  logic [0:0] f1078_clk;
  logic [0:0] f1078_rst;
  logic [31:0] f1078_rdata;
  sr_buffer_32_1 f1078(.wen(f1078_wen), .wdata(f1078_wdata), .clk(f1078_clk), .rst(f1078_rst), .rdata(f1078_rdata));
  assign f1078_clk = clk;
  assign f1078_rst = rst;
  // Bindings to f1078

  // f1080
  logic [0:0] f1080_wen;
  logic [31:0] f1080_wdata;
  logic [0:0] f1080_clk;
  logic [0:0] f1080_rst;
  logic [31:0] f1080_rdata;
  sr_buffer_32_1 f1080(.wen(f1080_wen), .wdata(f1080_wdata), .clk(f1080_clk), .rst(f1080_rst), .rdata(f1080_rdata));
  assign f1080_clk = clk;
  assign f1080_rst = rst;
  // Bindings to f1080

  // f1082
  logic [0:0] f1082_wen;
  logic [31:0] f1082_wdata;
  logic [0:0] f1082_clk;
  logic [0:0] f1082_rst;
  logic [31:0] f1082_rdata;
  sr_buffer_32_1 f1082(.wen(f1082_wen), .wdata(f1082_wdata), .clk(f1082_clk), .rst(f1082_rst), .rdata(f1082_rdata));
  assign f1082_clk = clk;
  assign f1082_rst = rst;
  // Bindings to f1082

  // f1084
  logic [0:0] f1084_wen;
  logic [31:0] f1084_wdata;
  logic [0:0] f1084_clk;
  logic [0:0] f1084_rst;
  logic [31:0] f1084_rdata;
  sr_buffer_32_1 f1084(.wen(f1084_wen), .wdata(f1084_wdata), .clk(f1084_clk), .rst(f1084_rst), .rdata(f1084_rdata));
  assign f1084_clk = clk;
  assign f1084_rst = rst;
  // Bindings to f1084

  // f1086
  logic [0:0] f1086_wen;
  logic [31:0] f1086_wdata;
  logic [0:0] f1086_clk;
  logic [0:0] f1086_rst;
  logic [31:0] f1086_rdata;
  sr_buffer_32_1 f1086(.wen(f1086_wen), .wdata(f1086_wdata), .clk(f1086_clk), .rst(f1086_rst), .rdata(f1086_rdata));
  assign f1086_clk = clk;
  assign f1086_rst = rst;
  // Bindings to f1086

  // f1088
  logic [0:0] f1088_wen;
  logic [31:0] f1088_wdata;
  logic [0:0] f1088_clk;
  logic [0:0] f1088_rst;
  logic [31:0] f1088_rdata;
  sr_buffer_32_1 f1088(.wen(f1088_wen), .wdata(f1088_wdata), .clk(f1088_clk), .rst(f1088_rst), .rdata(f1088_rdata));
  assign f1088_clk = clk;
  assign f1088_rst = rst;
  // Bindings to f1088

  // f1090
  logic [0:0] f1090_wen;
  logic [31:0] f1090_wdata;
  logic [0:0] f1090_clk;
  logic [0:0] f1090_rst;
  logic [31:0] f1090_rdata;
  sr_buffer_32_1 f1090(.wen(f1090_wen), .wdata(f1090_wdata), .clk(f1090_clk), .rst(f1090_rst), .rdata(f1090_rdata));
  assign f1090_clk = clk;
  assign f1090_rst = rst;
  // Bindings to f1090

  // f1092
  logic [0:0] f1092_wen;
  logic [31:0] f1092_wdata;
  logic [0:0] f1092_clk;
  logic [0:0] f1092_rst;
  logic [31:0] f1092_rdata;
  sr_buffer_32_1 f1092(.wen(f1092_wen), .wdata(f1092_wdata), .clk(f1092_clk), .rst(f1092_rst), .rdata(f1092_rdata));
  assign f1092_clk = clk;
  assign f1092_rst = rst;
  // Bindings to f1092

  // f1094
  logic [0:0] f1094_wen;
  logic [31:0] f1094_wdata;
  logic [0:0] f1094_clk;
  logic [0:0] f1094_rst;
  logic [31:0] f1094_rdata;
  sr_buffer_32_1 f1094(.wen(f1094_wen), .wdata(f1094_wdata), .clk(f1094_clk), .rst(f1094_rst), .rdata(f1094_rdata));
  assign f1094_clk = clk;
  assign f1094_rst = rst;
  // Bindings to f1094

  // f1096
  logic [0:0] f1096_wen;
  logic [31:0] f1096_wdata;
  logic [0:0] f1096_clk;
  logic [0:0] f1096_rst;
  logic [31:0] f1096_rdata;
  sr_buffer_32_1 f1096(.wen(f1096_wen), .wdata(f1096_wdata), .clk(f1096_clk), .rst(f1096_rst), .rdata(f1096_rdata));
  assign f1096_clk = clk;
  assign f1096_rst = rst;
  // Bindings to f1096

  // f1098
  logic [0:0] f1098_wen;
  logic [31:0] f1098_wdata;
  logic [0:0] f1098_clk;
  logic [0:0] f1098_rst;
  logic [31:0] f1098_rdata;
  sr_buffer_32_1 f1098(.wen(f1098_wen), .wdata(f1098_wdata), .clk(f1098_clk), .rst(f1098_rst), .rdata(f1098_rdata));
  assign f1098_clk = clk;
  assign f1098_rst = rst;
  // Bindings to f1098

  // f1100
  logic [0:0] f1100_wen;
  logic [31:0] f1100_wdata;
  logic [0:0] f1100_clk;
  logic [0:0] f1100_rst;
  logic [31:0] f1100_rdata;
  sr_buffer_32_1 f1100(.wen(f1100_wen), .wdata(f1100_wdata), .clk(f1100_clk), .rst(f1100_rst), .rdata(f1100_rdata));
  assign f1100_clk = clk;
  assign f1100_rst = rst;
  // Bindings to f1100

  // f1102
  logic [0:0] f1102_wen;
  logic [31:0] f1102_wdata;
  logic [0:0] f1102_clk;
  logic [0:0] f1102_rst;
  logic [31:0] f1102_rdata;
  sr_buffer_32_1 f1102(.wen(f1102_wen), .wdata(f1102_wdata), .clk(f1102_clk), .rst(f1102_rst), .rdata(f1102_rdata));
  assign f1102_clk = clk;
  assign f1102_rst = rst;
  // Bindings to f1102

  // f1104
  logic [0:0] f1104_wen;
  logic [31:0] f1104_wdata;
  logic [0:0] f1104_clk;
  logic [0:0] f1104_rst;
  logic [31:0] f1104_rdata;
  sr_buffer_32_1 f1104(.wen(f1104_wen), .wdata(f1104_wdata), .clk(f1104_clk), .rst(f1104_rst), .rdata(f1104_rdata));
  assign f1104_clk = clk;
  assign f1104_rst = rst;
  // Bindings to f1104

  // f1106
  logic [0:0] f1106_wen;
  logic [31:0] f1106_wdata;
  logic [0:0] f1106_clk;
  logic [0:0] f1106_rst;
  logic [31:0] f1106_rdata;
  sr_buffer_32_1 f1106(.wen(f1106_wen), .wdata(f1106_wdata), .clk(f1106_clk), .rst(f1106_rst), .rdata(f1106_rdata));
  assign f1106_clk = clk;
  assign f1106_rst = rst;
  // Bindings to f1106

  // f1108
  logic [0:0] f1108_wen;
  logic [31:0] f1108_wdata;
  logic [0:0] f1108_clk;
  logic [0:0] f1108_rst;
  logic [31:0] f1108_rdata;
  sr_buffer_32_1 f1108(.wen(f1108_wen), .wdata(f1108_wdata), .clk(f1108_clk), .rst(f1108_rst), .rdata(f1108_rdata));
  assign f1108_clk = clk;
  assign f1108_rst = rst;
  // Bindings to f1108

  // f1110
  logic [0:0] f1110_wen;
  logic [31:0] f1110_wdata;
  logic [0:0] f1110_clk;
  logic [0:0] f1110_rst;
  logic [31:0] f1110_rdata;
  sr_buffer_32_1 f1110(.wen(f1110_wen), .wdata(f1110_wdata), .clk(f1110_clk), .rst(f1110_rst), .rdata(f1110_rdata));
  assign f1110_clk = clk;
  assign f1110_rst = rst;
  // Bindings to f1110

  // f1112
  logic [0:0] f1112_wen;
  logic [31:0] f1112_wdata;
  logic [0:0] f1112_clk;
  logic [0:0] f1112_rst;
  logic [31:0] f1112_rdata;
  sr_buffer_32_1 f1112(.wen(f1112_wen), .wdata(f1112_wdata), .clk(f1112_clk), .rst(f1112_rst), .rdata(f1112_rdata));
  assign f1112_clk = clk;
  assign f1112_rst = rst;
  // Bindings to f1112

  // f1114
  logic [0:0] f1114_wen;
  logic [31:0] f1114_wdata;
  logic [0:0] f1114_clk;
  logic [0:0] f1114_rst;
  logic [31:0] f1114_rdata;
  sr_buffer_32_1 f1114(.wen(f1114_wen), .wdata(f1114_wdata), .clk(f1114_clk), .rst(f1114_rst), .rdata(f1114_rdata));
  assign f1114_clk = clk;
  assign f1114_rst = rst;
  // Bindings to f1114

  // f1116
  logic [0:0] f1116_wen;
  logic [31:0] f1116_wdata;
  logic [0:0] f1116_clk;
  logic [0:0] f1116_rst;
  logic [31:0] f1116_rdata;
  sr_buffer_32_1 f1116(.wen(f1116_wen), .wdata(f1116_wdata), .clk(f1116_clk), .rst(f1116_rst), .rdata(f1116_rdata));
  assign f1116_clk = clk;
  assign f1116_rst = rst;
  // Bindings to f1116

  // f1118
  logic [0:0] f1118_wen;
  logic [31:0] f1118_wdata;
  logic [0:0] f1118_clk;
  logic [0:0] f1118_rst;
  logic [31:0] f1118_rdata;
  sr_buffer_32_1 f1118(.wen(f1118_wen), .wdata(f1118_wdata), .clk(f1118_clk), .rst(f1118_rst), .rdata(f1118_rdata));
  assign f1118_clk = clk;
  assign f1118_rst = rst;
  // Bindings to f1118

  // f1120
  logic [0:0] f1120_wen;
  logic [31:0] f1120_wdata;
  logic [0:0] f1120_clk;
  logic [0:0] f1120_rst;
  logic [31:0] f1120_rdata;
  sr_buffer_32_1 f1120(.wen(f1120_wen), .wdata(f1120_wdata), .clk(f1120_clk), .rst(f1120_rst), .rdata(f1120_rdata));
  assign f1120_clk = clk;
  assign f1120_rst = rst;
  // Bindings to f1120

  // f1122
  logic [0:0] f1122_wen;
  logic [31:0] f1122_wdata;
  logic [0:0] f1122_clk;
  logic [0:0] f1122_rst;
  logic [31:0] f1122_rdata;
  sr_buffer_32_1 f1122(.wen(f1122_wen), .wdata(f1122_wdata), .clk(f1122_clk), .rst(f1122_rst), .rdata(f1122_rdata));
  assign f1122_clk = clk;
  assign f1122_rst = rst;
  // Bindings to f1122

  // f1124
  logic [0:0] f1124_wen;
  logic [31:0] f1124_wdata;
  logic [0:0] f1124_clk;
  logic [0:0] f1124_rst;
  logic [31:0] f1124_rdata;
  sr_buffer_32_1 f1124(.wen(f1124_wen), .wdata(f1124_wdata), .clk(f1124_clk), .rst(f1124_rst), .rdata(f1124_rdata));
  assign f1124_clk = clk;
  assign f1124_rst = rst;
  // Bindings to f1124

  // f1126
  logic [0:0] f1126_wen;
  logic [31:0] f1126_wdata;
  logic [0:0] f1126_clk;
  logic [0:0] f1126_rst;
  logic [31:0] f1126_rdata;
  sr_buffer_32_1 f1126(.wen(f1126_wen), .wdata(f1126_wdata), .clk(f1126_clk), .rst(f1126_rst), .rdata(f1126_rdata));
  assign f1126_clk = clk;
  assign f1126_rst = rst;
  // Bindings to f1126

  // f1128
  logic [0:0] f1128_wen;
  logic [31:0] f1128_wdata;
  logic [0:0] f1128_clk;
  logic [0:0] f1128_rst;
  logic [31:0] f1128_rdata;
  sr_buffer_32_1 f1128(.wen(f1128_wen), .wdata(f1128_wdata), .clk(f1128_clk), .rst(f1128_rst), .rdata(f1128_rdata));
  assign f1128_clk = clk;
  assign f1128_rst = rst;
  // Bindings to f1128

  // f1130
  logic [0:0] f1130_wen;
  logic [31:0] f1130_wdata;
  logic [0:0] f1130_clk;
  logic [0:0] f1130_rst;
  logic [31:0] f1130_rdata;
  sr_buffer_32_1 f1130(.wen(f1130_wen), .wdata(f1130_wdata), .clk(f1130_clk), .rst(f1130_rst), .rdata(f1130_rdata));
  assign f1130_clk = clk;
  assign f1130_rst = rst;
  // Bindings to f1130

  // f1132
  logic [0:0] f1132_wen;
  logic [31:0] f1132_wdata;
  logic [0:0] f1132_clk;
  logic [0:0] f1132_rst;
  logic [31:0] f1132_rdata;
  sr_buffer_32_1 f1132(.wen(f1132_wen), .wdata(f1132_wdata), .clk(f1132_clk), .rst(f1132_rst), .rdata(f1132_rdata));
  assign f1132_clk = clk;
  assign f1132_rst = rst;
  // Bindings to f1132

  // f1134
  logic [0:0] f1134_wen;
  logic [31:0] f1134_wdata;
  logic [0:0] f1134_clk;
  logic [0:0] f1134_rst;
  logic [31:0] f1134_rdata;
  sr_buffer_32_1 f1134(.wen(f1134_wen), .wdata(f1134_wdata), .clk(f1134_clk), .rst(f1134_rst), .rdata(f1134_rdata));
  assign f1134_clk = clk;
  assign f1134_rst = rst;
  // Bindings to f1134

  // f1136
  logic [0:0] f1136_wen;
  logic [31:0] f1136_wdata;
  logic [0:0] f1136_clk;
  logic [0:0] f1136_rst;
  logic [31:0] f1136_rdata;
  sr_buffer_32_1 f1136(.wen(f1136_wen), .wdata(f1136_wdata), .clk(f1136_clk), .rst(f1136_rst), .rdata(f1136_rdata));
  assign f1136_clk = clk;
  assign f1136_rst = rst;
  // Bindings to f1136

  // f1138
  logic [0:0] f1138_wen;
  logic [31:0] f1138_wdata;
  logic [0:0] f1138_clk;
  logic [0:0] f1138_rst;
  logic [31:0] f1138_rdata;
  sr_buffer_32_1 f1138(.wen(f1138_wen), .wdata(f1138_wdata), .clk(f1138_clk), .rst(f1138_rst), .rdata(f1138_rdata));
  assign f1138_clk = clk;
  assign f1138_rst = rst;
  // Bindings to f1138

  // f1140
  logic [0:0] f1140_wen;
  logic [31:0] f1140_wdata;
  logic [0:0] f1140_clk;
  logic [0:0] f1140_rst;
  logic [31:0] f1140_rdata;
  sr_buffer_32_1 f1140(.wen(f1140_wen), .wdata(f1140_wdata), .clk(f1140_clk), .rst(f1140_rst), .rdata(f1140_rdata));
  assign f1140_clk = clk;
  assign f1140_rst = rst;
  // Bindings to f1140

  // f1142
  logic [0:0] f1142_wen;
  logic [31:0] f1142_wdata;
  logic [0:0] f1142_clk;
  logic [0:0] f1142_rst;
  logic [31:0] f1142_rdata;
  sr_buffer_32_1 f1142(.wen(f1142_wen), .wdata(f1142_wdata), .clk(f1142_clk), .rst(f1142_rst), .rdata(f1142_rdata));
  assign f1142_clk = clk;
  assign f1142_rst = rst;
  // Bindings to f1142

  // f1144
  logic [0:0] f1144_wen;
  logic [31:0] f1144_wdata;
  logic [0:0] f1144_clk;
  logic [0:0] f1144_rst;
  logic [31:0] f1144_rdata;
  sr_buffer_32_1 f1144(.wen(f1144_wen), .wdata(f1144_wdata), .clk(f1144_clk), .rst(f1144_rst), .rdata(f1144_rdata));
  assign f1144_clk = clk;
  assign f1144_rst = rst;
  // Bindings to f1144

  // f1146
  logic [0:0] f1146_wen;
  logic [31:0] f1146_wdata;
  logic [0:0] f1146_clk;
  logic [0:0] f1146_rst;
  logic [31:0] f1146_rdata;
  sr_buffer_32_1 f1146(.wen(f1146_wen), .wdata(f1146_wdata), .clk(f1146_clk), .rst(f1146_rst), .rdata(f1146_rdata));
  assign f1146_clk = clk;
  assign f1146_rst = rst;
  // Bindings to f1146

  // f1148
  logic [0:0] f1148_wen;
  logic [31:0] f1148_wdata;
  logic [0:0] f1148_clk;
  logic [0:0] f1148_rst;
  logic [31:0] f1148_rdata;
  sr_buffer_32_1 f1148(.wen(f1148_wen), .wdata(f1148_wdata), .clk(f1148_clk), .rst(f1148_rst), .rdata(f1148_rdata));
  assign f1148_clk = clk;
  assign f1148_rst = rst;
  // Bindings to f1148

  // f1150
  logic [0:0] f1150_wen;
  logic [31:0] f1150_wdata;
  logic [0:0] f1150_clk;
  logic [0:0] f1150_rst;
  logic [31:0] f1150_rdata;
  sr_buffer_32_1 f1150(.wen(f1150_wen), .wdata(f1150_wdata), .clk(f1150_clk), .rst(f1150_rst), .rdata(f1150_rdata));
  assign f1150_clk = clk;
  assign f1150_rst = rst;
  // Bindings to f1150

  // f1152
  logic [0:0] f1152_wen;
  logic [31:0] f1152_wdata;
  logic [0:0] f1152_clk;
  logic [0:0] f1152_rst;
  logic [31:0] f1152_rdata;
  sr_buffer_32_1 f1152(.wen(f1152_wen), .wdata(f1152_wdata), .clk(f1152_clk), .rst(f1152_rst), .rdata(f1152_rdata));
  assign f1152_clk = clk;
  assign f1152_rst = rst;
  // Bindings to f1152

  // f1154
  logic [0:0] f1154_wen;
  logic [31:0] f1154_wdata;
  logic [0:0] f1154_clk;
  logic [0:0] f1154_rst;
  logic [31:0] f1154_rdata;
  sr_buffer_32_1 f1154(.wen(f1154_wen), .wdata(f1154_wdata), .clk(f1154_clk), .rst(f1154_rst), .rdata(f1154_rdata));
  assign f1154_clk = clk;
  assign f1154_rst = rst;
  // Bindings to f1154

  // f1156
  logic [0:0] f1156_wen;
  logic [31:0] f1156_wdata;
  logic [0:0] f1156_clk;
  logic [0:0] f1156_rst;
  logic [31:0] f1156_rdata;
  sr_buffer_32_1 f1156(.wen(f1156_wen), .wdata(f1156_wdata), .clk(f1156_clk), .rst(f1156_rst), .rdata(f1156_rdata));
  assign f1156_clk = clk;
  assign f1156_rst = rst;
  // Bindings to f1156

  // f1158
  logic [0:0] f1158_wen;
  logic [31:0] f1158_wdata;
  logic [0:0] f1158_clk;
  logic [0:0] f1158_rst;
  logic [31:0] f1158_rdata;
  sr_buffer_32_1 f1158(.wen(f1158_wen), .wdata(f1158_wdata), .clk(f1158_clk), .rst(f1158_rst), .rdata(f1158_rdata));
  assign f1158_clk = clk;
  assign f1158_rst = rst;
  // Bindings to f1158

  // f1160
  logic [0:0] f1160_wen;
  logic [31:0] f1160_wdata;
  logic [0:0] f1160_clk;
  logic [0:0] f1160_rst;
  logic [31:0] f1160_rdata;
  sr_buffer_32_1 f1160(.wen(f1160_wen), .wdata(f1160_wdata), .clk(f1160_clk), .rst(f1160_rst), .rdata(f1160_rdata));
  assign f1160_clk = clk;
  assign f1160_rst = rst;
  // Bindings to f1160

  // f1162
  logic [0:0] f1162_wen;
  logic [31:0] f1162_wdata;
  logic [0:0] f1162_clk;
  logic [0:0] f1162_rst;
  logic [31:0] f1162_rdata;
  sr_buffer_32_1 f1162(.wen(f1162_wen), .wdata(f1162_wdata), .clk(f1162_clk), .rst(f1162_rst), .rdata(f1162_rdata));
  assign f1162_clk = clk;
  assign f1162_rst = rst;
  // Bindings to f1162

  // f1164
  logic [0:0] f1164_wen;
  logic [31:0] f1164_wdata;
  logic [0:0] f1164_clk;
  logic [0:0] f1164_rst;
  logic [31:0] f1164_rdata;
  sr_buffer_32_1 f1164(.wen(f1164_wen), .wdata(f1164_wdata), .clk(f1164_clk), .rst(f1164_rst), .rdata(f1164_rdata));
  assign f1164_clk = clk;
  assign f1164_rst = rst;
  // Bindings to f1164

  // f1166
  logic [0:0] f1166_wen;
  logic [31:0] f1166_wdata;
  logic [0:0] f1166_clk;
  logic [0:0] f1166_rst;
  logic [31:0] f1166_rdata;
  sr_buffer_32_1 f1166(.wen(f1166_wen), .wdata(f1166_wdata), .clk(f1166_clk), .rst(f1166_rst), .rdata(f1166_rdata));
  assign f1166_clk = clk;
  assign f1166_rst = rst;
  // Bindings to f1166

  // f1168
  logic [0:0] f1168_wen;
  logic [31:0] f1168_wdata;
  logic [0:0] f1168_clk;
  logic [0:0] f1168_rst;
  logic [31:0] f1168_rdata;
  sr_buffer_32_1 f1168(.wen(f1168_wen), .wdata(f1168_wdata), .clk(f1168_clk), .rst(f1168_rst), .rdata(f1168_rdata));
  assign f1168_clk = clk;
  assign f1168_rst = rst;
  // Bindings to f1168

  // f1170
  logic [0:0] f1170_wen;
  logic [31:0] f1170_wdata;
  logic [0:0] f1170_clk;
  logic [0:0] f1170_rst;
  logic [31:0] f1170_rdata;
  sr_buffer_32_1 f1170(.wen(f1170_wen), .wdata(f1170_wdata), .clk(f1170_clk), .rst(f1170_rst), .rdata(f1170_rdata));
  assign f1170_clk = clk;
  assign f1170_rst = rst;
  // Bindings to f1170

  // f1172
  logic [0:0] f1172_wen;
  logic [31:0] f1172_wdata;
  logic [0:0] f1172_clk;
  logic [0:0] f1172_rst;
  logic [31:0] f1172_rdata;
  sr_buffer_32_1 f1172(.wen(f1172_wen), .wdata(f1172_wdata), .clk(f1172_clk), .rst(f1172_rst), .rdata(f1172_rdata));
  assign f1172_clk = clk;
  assign f1172_rst = rst;
  // Bindings to f1172

  // f1174
  logic [0:0] f1174_wen;
  logic [31:0] f1174_wdata;
  logic [0:0] f1174_clk;
  logic [0:0] f1174_rst;
  logic [31:0] f1174_rdata;
  sr_buffer_32_1 f1174(.wen(f1174_wen), .wdata(f1174_wdata), .clk(f1174_clk), .rst(f1174_rst), .rdata(f1174_rdata));
  assign f1174_clk = clk;
  assign f1174_rst = rst;
  // Bindings to f1174

  // f1176
  logic [0:0] f1176_wen;
  logic [31:0] f1176_wdata;
  logic [0:0] f1176_clk;
  logic [0:0] f1176_rst;
  logic [31:0] f1176_rdata;
  sr_buffer_32_1 f1176(.wen(f1176_wen), .wdata(f1176_wdata), .clk(f1176_clk), .rst(f1176_rst), .rdata(f1176_rdata));
  assign f1176_clk = clk;
  assign f1176_rst = rst;
  // Bindings to f1176

  // f1178
  logic [0:0] f1178_wen;
  logic [31:0] f1178_wdata;
  logic [0:0] f1178_clk;
  logic [0:0] f1178_rst;
  logic [31:0] f1178_rdata;
  sr_buffer_32_1 f1178(.wen(f1178_wen), .wdata(f1178_wdata), .clk(f1178_clk), .rst(f1178_rst), .rdata(f1178_rdata));
  assign f1178_clk = clk;
  assign f1178_rst = rst;
  // Bindings to f1178

  // f1180
  logic [0:0] f1180_wen;
  logic [31:0] f1180_wdata;
  logic [0:0] f1180_clk;
  logic [0:0] f1180_rst;
  logic [31:0] f1180_rdata;
  sr_buffer_32_1 f1180(.wen(f1180_wen), .wdata(f1180_wdata), .clk(f1180_clk), .rst(f1180_rst), .rdata(f1180_rdata));
  assign f1180_clk = clk;
  assign f1180_rst = rst;
  // Bindings to f1180

  // f1182
  logic [0:0] f1182_wen;
  logic [31:0] f1182_wdata;
  logic [0:0] f1182_clk;
  logic [0:0] f1182_rst;
  logic [31:0] f1182_rdata;
  sr_buffer_32_1 f1182(.wen(f1182_wen), .wdata(f1182_wdata), .clk(f1182_clk), .rst(f1182_rst), .rdata(f1182_rdata));
  assign f1182_clk = clk;
  assign f1182_rst = rst;
  // Bindings to f1182

  // f1184
  logic [0:0] f1184_wen;
  logic [31:0] f1184_wdata;
  logic [0:0] f1184_clk;
  logic [0:0] f1184_rst;
  logic [31:0] f1184_rdata;
  sr_buffer_32_1 f1184(.wen(f1184_wen), .wdata(f1184_wdata), .clk(f1184_clk), .rst(f1184_rst), .rdata(f1184_rdata));
  assign f1184_clk = clk;
  assign f1184_rst = rst;
  // Bindings to f1184

  // f1186
  logic [0:0] f1186_wen;
  logic [31:0] f1186_wdata;
  logic [0:0] f1186_clk;
  logic [0:0] f1186_rst;
  logic [31:0] f1186_rdata;
  sr_buffer_32_1 f1186(.wen(f1186_wen), .wdata(f1186_wdata), .clk(f1186_clk), .rst(f1186_rst), .rdata(f1186_rdata));
  assign f1186_clk = clk;
  assign f1186_rst = rst;
  // Bindings to f1186

  // f1188
  logic [0:0] f1188_wen;
  logic [31:0] f1188_wdata;
  logic [0:0] f1188_clk;
  logic [0:0] f1188_rst;
  logic [31:0] f1188_rdata;
  sr_buffer_32_1 f1188(.wen(f1188_wen), .wdata(f1188_wdata), .clk(f1188_clk), .rst(f1188_rst), .rdata(f1188_rdata));
  assign f1188_clk = clk;
  assign f1188_rst = rst;
  // Bindings to f1188

  // f1190
  logic [0:0] f1190_wen;
  logic [31:0] f1190_wdata;
  logic [0:0] f1190_clk;
  logic [0:0] f1190_rst;
  logic [31:0] f1190_rdata;
  sr_buffer_32_1 f1190(.wen(f1190_wen), .wdata(f1190_wdata), .clk(f1190_clk), .rst(f1190_rst), .rdata(f1190_rdata));
  assign f1190_clk = clk;
  assign f1190_rst = rst;
  // Bindings to f1190

  // f1192
  logic [0:0] f1192_wen;
  logic [31:0] f1192_wdata;
  logic [0:0] f1192_clk;
  logic [0:0] f1192_rst;
  logic [31:0] f1192_rdata;
  sr_buffer_32_1 f1192(.wen(f1192_wen), .wdata(f1192_wdata), .clk(f1192_clk), .rst(f1192_rst), .rdata(f1192_rdata));
  assign f1192_clk = clk;
  assign f1192_rst = rst;
  // Bindings to f1192

  // f1194
  logic [0:0] f1194_wen;
  logic [31:0] f1194_wdata;
  logic [0:0] f1194_clk;
  logic [0:0] f1194_rst;
  logic [31:0] f1194_rdata;
  sr_buffer_32_1 f1194(.wen(f1194_wen), .wdata(f1194_wdata), .clk(f1194_clk), .rst(f1194_rst), .rdata(f1194_rdata));
  assign f1194_clk = clk;
  assign f1194_rst = rst;
  // Bindings to f1194

  // f1196
  logic [0:0] f1196_wen;
  logic [31:0] f1196_wdata;
  logic [0:0] f1196_clk;
  logic [0:0] f1196_rst;
  logic [31:0] f1196_rdata;
  sr_buffer_32_1 f1196(.wen(f1196_wen), .wdata(f1196_wdata), .clk(f1196_clk), .rst(f1196_rst), .rdata(f1196_rdata));
  assign f1196_clk = clk;
  assign f1196_rst = rst;
  // Bindings to f1196

  // f1198
  logic [0:0] f1198_wen;
  logic [31:0] f1198_wdata;
  logic [0:0] f1198_clk;
  logic [0:0] f1198_rst;
  logic [31:0] f1198_rdata;
  sr_buffer_32_1 f1198(.wen(f1198_wen), .wdata(f1198_wdata), .clk(f1198_clk), .rst(f1198_rst), .rdata(f1198_rdata));
  assign f1198_clk = clk;
  assign f1198_rst = rst;
  // Bindings to f1198

  // f1200
  logic [0:0] f1200_wen;
  logic [31:0] f1200_wdata;
  logic [0:0] f1200_clk;
  logic [0:0] f1200_rst;
  logic [31:0] f1200_rdata;
  sr_buffer_32_1 f1200(.wen(f1200_wen), .wdata(f1200_wdata), .clk(f1200_clk), .rst(f1200_rst), .rdata(f1200_rdata));
  assign f1200_clk = clk;
  assign f1200_rst = rst;
  // Bindings to f1200

  // f1202
  logic [0:0] f1202_wen;
  logic [31:0] f1202_wdata;
  logic [0:0] f1202_clk;
  logic [0:0] f1202_rst;
  logic [31:0] f1202_rdata;
  sr_buffer_32_1 f1202(.wen(f1202_wen), .wdata(f1202_wdata), .clk(f1202_clk), .rst(f1202_rst), .rdata(f1202_rdata));
  assign f1202_clk = clk;
  assign f1202_rst = rst;
  // Bindings to f1202

  // f1204
  logic [0:0] f1204_wen;
  logic [31:0] f1204_wdata;
  logic [0:0] f1204_clk;
  logic [0:0] f1204_rst;
  logic [31:0] f1204_rdata;
  sr_buffer_32_1 f1204(.wen(f1204_wen), .wdata(f1204_wdata), .clk(f1204_clk), .rst(f1204_rst), .rdata(f1204_rdata));
  assign f1204_clk = clk;
  assign f1204_rst = rst;
  // Bindings to f1204

  // f1206
  logic [0:0] f1206_wen;
  logic [31:0] f1206_wdata;
  logic [0:0] f1206_clk;
  logic [0:0] f1206_rst;
  logic [31:0] f1206_rdata;
  sr_buffer_32_1 f1206(.wen(f1206_wen), .wdata(f1206_wdata), .clk(f1206_clk), .rst(f1206_rst), .rdata(f1206_rdata));
  assign f1206_clk = clk;
  assign f1206_rst = rst;
  // Bindings to f1206

  // f1208
  logic [0:0] f1208_wen;
  logic [31:0] f1208_wdata;
  logic [0:0] f1208_clk;
  logic [0:0] f1208_rst;
  logic [31:0] f1208_rdata;
  sr_buffer_32_1 f1208(.wen(f1208_wen), .wdata(f1208_wdata), .clk(f1208_clk), .rst(f1208_rst), .rdata(f1208_rdata));
  assign f1208_clk = clk;
  assign f1208_rst = rst;
  // Bindings to f1208

  // f1210
  logic [0:0] f1210_wen;
  logic [31:0] f1210_wdata;
  logic [0:0] f1210_clk;
  logic [0:0] f1210_rst;
  logic [31:0] f1210_rdata;
  sr_buffer_32_1 f1210(.wen(f1210_wen), .wdata(f1210_wdata), .clk(f1210_clk), .rst(f1210_rst), .rdata(f1210_rdata));
  assign f1210_clk = clk;
  assign f1210_rst = rst;
  // Bindings to f1210

  // f1212
  logic [0:0] f1212_wen;
  logic [31:0] f1212_wdata;
  logic [0:0] f1212_clk;
  logic [0:0] f1212_rst;
  logic [31:0] f1212_rdata;
  sr_buffer_32_1 f1212(.wen(f1212_wen), .wdata(f1212_wdata), .clk(f1212_clk), .rst(f1212_rst), .rdata(f1212_rdata));
  assign f1212_clk = clk;
  assign f1212_rst = rst;
  // Bindings to f1212

  // f1214
  logic [0:0] f1214_wen;
  logic [31:0] f1214_wdata;
  logic [0:0] f1214_clk;
  logic [0:0] f1214_rst;
  logic [31:0] f1214_rdata;
  sr_buffer_32_1 f1214(.wen(f1214_wen), .wdata(f1214_wdata), .clk(f1214_clk), .rst(f1214_rst), .rdata(f1214_rdata));
  assign f1214_clk = clk;
  assign f1214_rst = rst;
  // Bindings to f1214

  // f1216
  logic [0:0] f1216_wen;
  logic [31:0] f1216_wdata;
  logic [0:0] f1216_clk;
  logic [0:0] f1216_rst;
  logic [31:0] f1216_rdata;
  sr_buffer_32_1 f1216(.wen(f1216_wen), .wdata(f1216_wdata), .clk(f1216_clk), .rst(f1216_rst), .rdata(f1216_rdata));
  assign f1216_clk = clk;
  assign f1216_rst = rst;
  // Bindings to f1216

  // f1218
  logic [0:0] f1218_wen;
  logic [31:0] f1218_wdata;
  logic [0:0] f1218_clk;
  logic [0:0] f1218_rst;
  logic [31:0] f1218_rdata;
  sr_buffer_32_1 f1218(.wen(f1218_wen), .wdata(f1218_wdata), .clk(f1218_clk), .rst(f1218_rst), .rdata(f1218_rdata));
  assign f1218_clk = clk;
  assign f1218_rst = rst;
  // Bindings to f1218

  // f1220
  logic [0:0] f1220_wen;
  logic [31:0] f1220_wdata;
  logic [0:0] f1220_clk;
  logic [0:0] f1220_rst;
  logic [31:0] f1220_rdata;
  sr_buffer_32_1 f1220(.wen(f1220_wen), .wdata(f1220_wdata), .clk(f1220_clk), .rst(f1220_rst), .rdata(f1220_rdata));
  assign f1220_clk = clk;
  assign f1220_rst = rst;
  // Bindings to f1220

  // f1222
  logic [0:0] f1222_wen;
  logic [31:0] f1222_wdata;
  logic [0:0] f1222_clk;
  logic [0:0] f1222_rst;
  logic [31:0] f1222_rdata;
  sr_buffer_32_1 f1222(.wen(f1222_wen), .wdata(f1222_wdata), .clk(f1222_clk), .rst(f1222_rst), .rdata(f1222_rdata));
  assign f1222_clk = clk;
  assign f1222_rst = rst;
  // Bindings to f1222

  // f1224
  logic [0:0] f1224_wen;
  logic [31:0] f1224_wdata;
  logic [0:0] f1224_clk;
  logic [0:0] f1224_rst;
  logic [31:0] f1224_rdata;
  sr_buffer_32_1 f1224(.wen(f1224_wen), .wdata(f1224_wdata), .clk(f1224_clk), .rst(f1224_rst), .rdata(f1224_rdata));
  assign f1224_clk = clk;
  assign f1224_rst = rst;
  // Bindings to f1224

  // f1226
  logic [0:0] f1226_wen;
  logic [31:0] f1226_wdata;
  logic [0:0] f1226_clk;
  logic [0:0] f1226_rst;
  logic [31:0] f1226_rdata;
  sr_buffer_32_1 f1226(.wen(f1226_wen), .wdata(f1226_wdata), .clk(f1226_clk), .rst(f1226_rst), .rdata(f1226_rdata));
  assign f1226_clk = clk;
  assign f1226_rst = rst;
  // Bindings to f1226

  // f1228
  logic [0:0] f1228_wen;
  logic [31:0] f1228_wdata;
  logic [0:0] f1228_clk;
  logic [0:0] f1228_rst;
  logic [31:0] f1228_rdata;
  sr_buffer_32_1 f1228(.wen(f1228_wen), .wdata(f1228_wdata), .clk(f1228_clk), .rst(f1228_rst), .rdata(f1228_rdata));
  assign f1228_clk = clk;
  assign f1228_rst = rst;
  // Bindings to f1228

  // f1230
  logic [0:0] f1230_wen;
  logic [31:0] f1230_wdata;
  logic [0:0] f1230_clk;
  logic [0:0] f1230_rst;
  logic [31:0] f1230_rdata;
  sr_buffer_32_1 f1230(.wen(f1230_wen), .wdata(f1230_wdata), .clk(f1230_clk), .rst(f1230_rst), .rdata(f1230_rdata));
  assign f1230_clk = clk;
  assign f1230_rst = rst;
  // Bindings to f1230

  // f1232
  logic [0:0] f1232_wen;
  logic [31:0] f1232_wdata;
  logic [0:0] f1232_clk;
  logic [0:0] f1232_rst;
  logic [31:0] f1232_rdata;
  sr_buffer_32_1 f1232(.wen(f1232_wen), .wdata(f1232_wdata), .clk(f1232_clk), .rst(f1232_rst), .rdata(f1232_rdata));
  assign f1232_clk = clk;
  assign f1232_rst = rst;
  // Bindings to f1232

  // f1234
  logic [0:0] f1234_wen;
  logic [31:0] f1234_wdata;
  logic [0:0] f1234_clk;
  logic [0:0] f1234_rst;
  logic [31:0] f1234_rdata;
  sr_buffer_32_1 f1234(.wen(f1234_wen), .wdata(f1234_wdata), .clk(f1234_clk), .rst(f1234_rst), .rdata(f1234_rdata));
  assign f1234_clk = clk;
  assign f1234_rst = rst;
  // Bindings to f1234

  // f1236
  logic [0:0] f1236_wen;
  logic [31:0] f1236_wdata;
  logic [0:0] f1236_clk;
  logic [0:0] f1236_rst;
  logic [31:0] f1236_rdata;
  sr_buffer_32_1 f1236(.wen(f1236_wen), .wdata(f1236_wdata), .clk(f1236_clk), .rst(f1236_rst), .rdata(f1236_rdata));
  assign f1236_clk = clk;
  assign f1236_rst = rst;
  // Bindings to f1236

  // f1238
  logic [0:0] f1238_wen;
  logic [31:0] f1238_wdata;
  logic [0:0] f1238_clk;
  logic [0:0] f1238_rst;
  logic [31:0] f1238_rdata;
  sr_buffer_32_1 f1238(.wen(f1238_wen), .wdata(f1238_wdata), .clk(f1238_clk), .rst(f1238_rst), .rdata(f1238_rdata));
  assign f1238_clk = clk;
  assign f1238_rst = rst;
  // Bindings to f1238

  // f1240
  logic [0:0] f1240_wen;
  logic [31:0] f1240_wdata;
  logic [0:0] f1240_clk;
  logic [0:0] f1240_rst;
  logic [31:0] f1240_rdata;
  sr_buffer_32_1 f1240(.wen(f1240_wen), .wdata(f1240_wdata), .clk(f1240_clk), .rst(f1240_rst), .rdata(f1240_rdata));
  assign f1240_clk = clk;
  assign f1240_rst = rst;
  // Bindings to f1240

  // f1242
  logic [0:0] f1242_wen;
  logic [31:0] f1242_wdata;
  logic [0:0] f1242_clk;
  logic [0:0] f1242_rst;
  logic [31:0] f1242_rdata;
  sr_buffer_32_1 f1242(.wen(f1242_wen), .wdata(f1242_wdata), .clk(f1242_clk), .rst(f1242_rst), .rdata(f1242_rdata));
  assign f1242_clk = clk;
  assign f1242_rst = rst;
  // Bindings to f1242

  // f1244
  logic [0:0] f1244_wen;
  logic [31:0] f1244_wdata;
  logic [0:0] f1244_clk;
  logic [0:0] f1244_rst;
  logic [31:0] f1244_rdata;
  sr_buffer_32_1 f1244(.wen(f1244_wen), .wdata(f1244_wdata), .clk(f1244_clk), .rst(f1244_rst), .rdata(f1244_rdata));
  assign f1244_clk = clk;
  assign f1244_rst = rst;
  // Bindings to f1244

  // f1246
  logic [0:0] f1246_wen;
  logic [31:0] f1246_wdata;
  logic [0:0] f1246_clk;
  logic [0:0] f1246_rst;
  logic [31:0] f1246_rdata;
  sr_buffer_32_1 f1246(.wen(f1246_wen), .wdata(f1246_wdata), .clk(f1246_clk), .rst(f1246_rst), .rdata(f1246_rdata));
  assign f1246_clk = clk;
  assign f1246_rst = rst;
  // Bindings to f1246

  // f1248
  logic [0:0] f1248_wen;
  logic [31:0] f1248_wdata;
  logic [0:0] f1248_clk;
  logic [0:0] f1248_rst;
  logic [31:0] f1248_rdata;
  sr_buffer_32_1 f1248(.wen(f1248_wen), .wdata(f1248_wdata), .clk(f1248_clk), .rst(f1248_rst), .rdata(f1248_rdata));
  assign f1248_clk = clk;
  assign f1248_rst = rst;
  // Bindings to f1248

  // f1250
  logic [0:0] f1250_wen;
  logic [31:0] f1250_wdata;
  logic [0:0] f1250_clk;
  logic [0:0] f1250_rst;
  logic [31:0] f1250_rdata;
  sr_buffer_32_1 f1250(.wen(f1250_wen), .wdata(f1250_wdata), .clk(f1250_clk), .rst(f1250_rst), .rdata(f1250_rdata));
  assign f1250_clk = clk;
  assign f1250_rst = rst;
  // Bindings to f1250

  // f1252
  logic [0:0] f1252_wen;
  logic [31:0] f1252_wdata;
  logic [0:0] f1252_clk;
  logic [0:0] f1252_rst;
  logic [31:0] f1252_rdata;
  sr_buffer_32_1 f1252(.wen(f1252_wen), .wdata(f1252_wdata), .clk(f1252_clk), .rst(f1252_rst), .rdata(f1252_rdata));
  assign f1252_clk = clk;
  assign f1252_rst = rst;
  // Bindings to f1252



endmodule


module bright_bright_update_0_write0_to_bright_laplace_diff_0_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_16431 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f2494
  logic [0:0] f2494_wen;
  logic [31:0] f2494_wdata;
  logic [0:0] f2494_clk;
  logic [0:0] f2494_rst;
  logic [31:0] f2494_rdata;
  sr_buffer_32_1 f2494(.wen(f2494_wen), .wdata(f2494_wdata), .clk(f2494_clk), .rst(f2494_rst), .rdata(f2494_rdata));
  assign f2494_clk = clk;
  assign f2494_rst = rst;
  // Bindings to f2494

  // f2496
  logic [0:0] f2496_wen;
  logic [31:0] f2496_wdata;
  logic [0:0] f2496_clk;
  logic [0:0] f2496_rst;
  logic [31:0] f2496_rdata;
  sr_buffer_32_1 f2496(.wen(f2496_wen), .wdata(f2496_wdata), .clk(f2496_clk), .rst(f2496_rst), .rdata(f2496_rdata));
  assign f2496_clk = clk;
  assign f2496_rst = rst;
  // Bindings to f2496

  // f2498
  logic [0:0] f2498_wen;
  logic [31:0] f2498_wdata;
  logic [0:0] f2498_clk;
  logic [0:0] f2498_rst;
  logic [31:0] f2498_rdata;
  sr_buffer_32_1 f2498(.wen(f2498_wen), .wdata(f2498_wdata), .clk(f2498_clk), .rst(f2498_rst), .rdata(f2498_rdata));
  assign f2498_clk = clk;
  assign f2498_rst = rst;
  // Bindings to f2498

  // f2500
  logic [0:0] f2500_wen;
  logic [31:0] f2500_wdata;
  logic [0:0] f2500_clk;
  logic [0:0] f2500_rst;
  logic [31:0] f2500_rdata;
  sr_buffer_32_1 f2500(.wen(f2500_wen), .wdata(f2500_wdata), .clk(f2500_clk), .rst(f2500_rst), .rdata(f2500_rdata));
  assign f2500_clk = clk;
  assign f2500_rst = rst;
  // Bindings to f2500

  // f2502
  logic [0:0] f2502_wen;
  logic [31:0] f2502_wdata;
  logic [0:0] f2502_clk;
  logic [0:0] f2502_rst;
  logic [31:0] f2502_rdata;
  sr_buffer_32_1 f2502(.wen(f2502_wen), .wdata(f2502_wdata), .clk(f2502_clk), .rst(f2502_rst), .rdata(f2502_rdata));
  assign f2502_clk = clk;
  assign f2502_rst = rst;
  // Bindings to f2502

  // f2504
  logic [0:0] f2504_wen;
  logic [31:0] f2504_wdata;
  logic [0:0] f2504_clk;
  logic [0:0] f2504_rst;
  logic [31:0] f2504_rdata;
  sr_buffer_32_1 f2504(.wen(f2504_wen), .wdata(f2504_wdata), .clk(f2504_clk), .rst(f2504_rst), .rdata(f2504_rdata));
  assign f2504_clk = clk;
  assign f2504_rst = rst;
  // Bindings to f2504

  // f2506
  logic [0:0] f2506_wen;
  logic [31:0] f2506_wdata;
  logic [0:0] f2506_clk;
  logic [0:0] f2506_rst;
  logic [31:0] f2506_rdata;
  sr_buffer_32_1 f2506(.wen(f2506_wen), .wdata(f2506_wdata), .clk(f2506_clk), .rst(f2506_rst), .rdata(f2506_rdata));
  assign f2506_clk = clk;
  assign f2506_rst = rst;
  // Bindings to f2506

  // f2508
  logic [0:0] f2508_wen;
  logic [31:0] f2508_wdata;
  logic [0:0] f2508_clk;
  logic [0:0] f2508_rst;
  logic [31:0] f2508_rdata;
  sr_buffer_32_1 f2508(.wen(f2508_wen), .wdata(f2508_wdata), .clk(f2508_clk), .rst(f2508_rst), .rdata(f2508_rdata));
  assign f2508_clk = clk;
  assign f2508_rst = rst;
  // Bindings to f2508

  // f2510
  logic [0:0] f2510_wen;
  logic [31:0] f2510_wdata;
  logic [0:0] f2510_clk;
  logic [0:0] f2510_rst;
  logic [31:0] f2510_rdata;
  sr_buffer_32_1 f2510(.wen(f2510_wen), .wdata(f2510_wdata), .clk(f2510_clk), .rst(f2510_rst), .rdata(f2510_rdata));
  assign f2510_clk = clk;
  assign f2510_rst = rst;
  // Bindings to f2510

  // f2512
  logic [0:0] f2512_wen;
  logic [31:0] f2512_wdata;
  logic [0:0] f2512_clk;
  logic [0:0] f2512_rst;
  logic [31:0] f2512_rdata;
  sr_buffer_32_1 f2512(.wen(f2512_wen), .wdata(f2512_wdata), .clk(f2512_clk), .rst(f2512_rst), .rdata(f2512_rdata));
  assign f2512_clk = clk;
  assign f2512_rst = rst;
  // Bindings to f2512

  // f2514
  logic [0:0] f2514_wen;
  logic [31:0] f2514_wdata;
  logic [0:0] f2514_clk;
  logic [0:0] f2514_rst;
  logic [31:0] f2514_rdata;
  sr_buffer_32_1 f2514(.wen(f2514_wen), .wdata(f2514_wdata), .clk(f2514_clk), .rst(f2514_rst), .rdata(f2514_rdata));
  assign f2514_clk = clk;
  assign f2514_rst = rst;
  // Bindings to f2514

  // f2516
  logic [0:0] f2516_wen;
  logic [31:0] f2516_wdata;
  logic [0:0] f2516_clk;
  logic [0:0] f2516_rst;
  logic [31:0] f2516_rdata;
  sr_buffer_32_1 f2516(.wen(f2516_wen), .wdata(f2516_wdata), .clk(f2516_clk), .rst(f2516_rst), .rdata(f2516_rdata));
  assign f2516_clk = clk;
  assign f2516_rst = rst;
  // Bindings to f2516

  // f2518
  logic [0:0] f2518_wen;
  logic [31:0] f2518_wdata;
  logic [0:0] f2518_clk;
  logic [0:0] f2518_rst;
  logic [31:0] f2518_rdata;
  sr_buffer_32_1 f2518(.wen(f2518_wen), .wdata(f2518_wdata), .clk(f2518_clk), .rst(f2518_rst), .rdata(f2518_rdata));
  assign f2518_clk = clk;
  assign f2518_rst = rst;
  // Bindings to f2518

  // f2520
  logic [0:0] f2520_wen;
  logic [31:0] f2520_wdata;
  logic [0:0] f2520_clk;
  logic [0:0] f2520_rst;
  logic [31:0] f2520_rdata;
  sr_buffer_32_1 f2520(.wen(f2520_wen), .wdata(f2520_wdata), .clk(f2520_clk), .rst(f2520_rst), .rdata(f2520_rdata));
  assign f2520_clk = clk;
  assign f2520_rst = rst;
  // Bindings to f2520

  // f2522
  logic [0:0] f2522_wen;
  logic [31:0] f2522_wdata;
  logic [0:0] f2522_clk;
  logic [0:0] f2522_rst;
  logic [31:0] f2522_rdata;
  sr_buffer_32_1 f2522(.wen(f2522_wen), .wdata(f2522_wdata), .clk(f2522_clk), .rst(f2522_rst), .rdata(f2522_rdata));
  assign f2522_clk = clk;
  assign f2522_rst = rst;
  // Bindings to f2522

  // f2524
  logic [0:0] f2524_wen;
  logic [31:0] f2524_wdata;
  logic [0:0] f2524_clk;
  logic [0:0] f2524_rst;
  logic [31:0] f2524_rdata;
  sr_buffer_32_1 f2524(.wen(f2524_wen), .wdata(f2524_wdata), .clk(f2524_clk), .rst(f2524_rst), .rdata(f2524_rdata));
  assign f2524_clk = clk;
  assign f2524_rst = rst;
  // Bindings to f2524

  // f2526
  logic [0:0] f2526_wen;
  logic [31:0] f2526_wdata;
  logic [0:0] f2526_clk;
  logic [0:0] f2526_rst;
  logic [31:0] f2526_rdata;
  sr_buffer_32_1 f2526(.wen(f2526_wen), .wdata(f2526_wdata), .clk(f2526_clk), .rst(f2526_rst), .rdata(f2526_rdata));
  assign f2526_clk = clk;
  assign f2526_rst = rst;
  // Bindings to f2526

  // f2528
  logic [0:0] f2528_wen;
  logic [31:0] f2528_wdata;
  logic [0:0] f2528_clk;
  logic [0:0] f2528_rst;
  logic [31:0] f2528_rdata;
  sr_buffer_32_1 f2528(.wen(f2528_wen), .wdata(f2528_wdata), .clk(f2528_clk), .rst(f2528_rst), .rdata(f2528_rdata));
  assign f2528_clk = clk;
  assign f2528_rst = rst;
  // Bindings to f2528

  // f2530
  logic [0:0] f2530_wen;
  logic [31:0] f2530_wdata;
  logic [0:0] f2530_clk;
  logic [0:0] f2530_rst;
  logic [31:0] f2530_rdata;
  sr_buffer_32_1 f2530(.wen(f2530_wen), .wdata(f2530_wdata), .clk(f2530_clk), .rst(f2530_rst), .rdata(f2530_rdata));
  assign f2530_clk = clk;
  assign f2530_rst = rst;
  // Bindings to f2530

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f458
  logic [0:0] f458_wen;
  logic [31:0] f458_wdata;
  logic [0:0] f458_clk;
  logic [0:0] f458_rst;
  logic [31:0] f458_rdata;
  sr_buffer_32_1 f458(.wen(f458_wen), .wdata(f458_wdata), .clk(f458_clk), .rst(f458_rst), .rdata(f458_rdata));
  assign f458_clk = clk;
  assign f458_rst = rst;
  // Bindings to f458

  // f460
  logic [0:0] f460_wen;
  logic [31:0] f460_wdata;
  logic [0:0] f460_clk;
  logic [0:0] f460_rst;
  logic [31:0] f460_rdata;
  sr_buffer_32_1 f460(.wen(f460_wen), .wdata(f460_wdata), .clk(f460_clk), .rst(f460_rst), .rdata(f460_rdata));
  assign f460_clk = clk;
  assign f460_rst = rst;
  // Bindings to f460

  // f462
  logic [0:0] f462_wen;
  logic [31:0] f462_wdata;
  logic [0:0] f462_clk;
  logic [0:0] f462_rst;
  logic [31:0] f462_rdata;
  sr_buffer_32_1 f462(.wen(f462_wen), .wdata(f462_wdata), .clk(f462_clk), .rst(f462_rst), .rdata(f462_rdata));
  assign f462_clk = clk;
  assign f462_rst = rst;
  // Bindings to f462

  // f464
  logic [0:0] f464_wen;
  logic [31:0] f464_wdata;
  logic [0:0] f464_clk;
  logic [0:0] f464_rst;
  logic [31:0] f464_rdata;
  sr_buffer_32_1 f464(.wen(f464_wen), .wdata(f464_wdata), .clk(f464_clk), .rst(f464_rst), .rdata(f464_rdata));
  assign f464_clk = clk;
  assign f464_rst = rst;
  // Bindings to f464

  // f466
  logic [0:0] f466_wen;
  logic [31:0] f466_wdata;
  logic [0:0] f466_clk;
  logic [0:0] f466_rst;
  logic [31:0] f466_rdata;
  sr_buffer_32_1 f466(.wen(f466_wen), .wdata(f466_wdata), .clk(f466_clk), .rst(f466_rst), .rdata(f466_rdata));
  assign f466_clk = clk;
  assign f466_rst = rst;
  // Bindings to f466

  // f468
  logic [0:0] f468_wen;
  logic [31:0] f468_wdata;
  logic [0:0] f468_clk;
  logic [0:0] f468_rst;
  logic [31:0] f468_rdata;
  sr_buffer_32_1 f468(.wen(f468_wen), .wdata(f468_wdata), .clk(f468_clk), .rst(f468_rst), .rdata(f468_rdata));
  assign f468_clk = clk;
  assign f468_rst = rst;
  // Bindings to f468

  // f470
  logic [0:0] f470_wen;
  logic [31:0] f470_wdata;
  logic [0:0] f470_clk;
  logic [0:0] f470_rst;
  logic [31:0] f470_rdata;
  sr_buffer_32_1 f470(.wen(f470_wen), .wdata(f470_wdata), .clk(f470_clk), .rst(f470_rst), .rdata(f470_rdata));
  assign f470_clk = clk;
  assign f470_rst = rst;
  // Bindings to f470

  // f472
  logic [0:0] f472_wen;
  logic [31:0] f472_wdata;
  logic [0:0] f472_clk;
  logic [0:0] f472_rst;
  logic [31:0] f472_rdata;
  sr_buffer_32_1 f472(.wen(f472_wen), .wdata(f472_wdata), .clk(f472_clk), .rst(f472_rst), .rdata(f472_rdata));
  assign f472_clk = clk;
  assign f472_rst = rst;
  // Bindings to f472

  // f474
  logic [0:0] f474_wen;
  logic [31:0] f474_wdata;
  logic [0:0] f474_clk;
  logic [0:0] f474_rst;
  logic [31:0] f474_rdata;
  sr_buffer_32_1 f474(.wen(f474_wen), .wdata(f474_wdata), .clk(f474_clk), .rst(f474_rst), .rdata(f474_rdata));
  assign f474_clk = clk;
  assign f474_rst = rst;
  // Bindings to f474

  // f476
  logic [0:0] f476_wen;
  logic [31:0] f476_wdata;
  logic [0:0] f476_clk;
  logic [0:0] f476_rst;
  logic [31:0] f476_rdata;
  sr_buffer_32_1 f476(.wen(f476_wen), .wdata(f476_wdata), .clk(f476_clk), .rst(f476_rst), .rdata(f476_rdata));
  assign f476_clk = clk;
  assign f476_rst = rst;
  // Bindings to f476

  // f478
  logic [0:0] f478_wen;
  logic [31:0] f478_wdata;
  logic [0:0] f478_clk;
  logic [0:0] f478_rst;
  logic [31:0] f478_rdata;
  sr_buffer_32_1 f478(.wen(f478_wen), .wdata(f478_wdata), .clk(f478_clk), .rst(f478_rst), .rdata(f478_rdata));
  assign f478_clk = clk;
  assign f478_rst = rst;
  // Bindings to f478

  // f480
  logic [0:0] f480_wen;
  logic [31:0] f480_wdata;
  logic [0:0] f480_clk;
  logic [0:0] f480_rst;
  logic [31:0] f480_rdata;
  sr_buffer_32_1 f480(.wen(f480_wen), .wdata(f480_wdata), .clk(f480_clk), .rst(f480_rst), .rdata(f480_rdata));
  assign f480_clk = clk;
  assign f480_rst = rst;
  // Bindings to f480

  // f482
  logic [0:0] f482_wen;
  logic [31:0] f482_wdata;
  logic [0:0] f482_clk;
  logic [0:0] f482_rst;
  logic [31:0] f482_rdata;
  sr_buffer_32_1 f482(.wen(f482_wen), .wdata(f482_wdata), .clk(f482_clk), .rst(f482_rst), .rdata(f482_rdata));
  assign f482_clk = clk;
  assign f482_rst = rst;
  // Bindings to f482

  // f484
  logic [0:0] f484_wen;
  logic [31:0] f484_wdata;
  logic [0:0] f484_clk;
  logic [0:0] f484_rst;
  logic [31:0] f484_rdata;
  sr_buffer_32_1 f484(.wen(f484_wen), .wdata(f484_wdata), .clk(f484_clk), .rst(f484_rst), .rdata(f484_rdata));
  assign f484_clk = clk;
  assign f484_rst = rst;
  // Bindings to f484

  // f486
  logic [0:0] f486_wen;
  logic [31:0] f486_wdata;
  logic [0:0] f486_clk;
  logic [0:0] f486_rst;
  logic [31:0] f486_rdata;
  sr_buffer_32_1 f486(.wen(f486_wen), .wdata(f486_wdata), .clk(f486_clk), .rst(f486_rst), .rdata(f486_rdata));
  assign f486_clk = clk;
  assign f486_rst = rst;
  // Bindings to f486

  // f502
  logic [0:0] f502_wen;
  logic [31:0] f502_wdata;
  logic [0:0] f502_clk;
  logic [0:0] f502_rst;
  logic [31:0] f502_rdata;
  sr_buffer_32_1 f502(.wen(f502_wen), .wdata(f502_wdata), .clk(f502_clk), .rst(f502_rst), .rdata(f502_rdata));
  assign f502_clk = clk;
  assign f502_rst = rst;
  // Bindings to f502

  // f504
  logic [0:0] f504_wen;
  logic [31:0] f504_wdata;
  logic [0:0] f504_clk;
  logic [0:0] f504_rst;
  logic [31:0] f504_rdata;
  sr_buffer_32_1 f504(.wen(f504_wen), .wdata(f504_wdata), .clk(f504_clk), .rst(f504_rst), .rdata(f504_rdata));
  assign f504_clk = clk;
  assign f504_rst = rst;
  // Bindings to f504

  // f506
  logic [0:0] f506_wen;
  logic [31:0] f506_wdata;
  logic [0:0] f506_clk;
  logic [0:0] f506_rst;
  logic [31:0] f506_rdata;
  sr_buffer_32_1 f506(.wen(f506_wen), .wdata(f506_wdata), .clk(f506_clk), .rst(f506_rst), .rdata(f506_rdata));
  assign f506_clk = clk;
  assign f506_rst = rst;
  // Bindings to f506

  // f508
  logic [0:0] f508_wen;
  logic [31:0] f508_wdata;
  logic [0:0] f508_clk;
  logic [0:0] f508_rst;
  logic [31:0] f508_rdata;
  sr_buffer_32_1 f508(.wen(f508_wen), .wdata(f508_wdata), .clk(f508_clk), .rst(f508_rst), .rdata(f508_rdata));
  assign f508_clk = clk;
  assign f508_rst = rst;
  // Bindings to f508

  // f510
  logic [0:0] f510_wen;
  logic [31:0] f510_wdata;
  logic [0:0] f510_clk;
  logic [0:0] f510_rst;
  logic [31:0] f510_rdata;
  sr_buffer_32_1 f510(.wen(f510_wen), .wdata(f510_wdata), .clk(f510_clk), .rst(f510_rst), .rdata(f510_rdata));
  assign f510_clk = clk;
  assign f510_rst = rst;
  // Bindings to f510

  // f512
  logic [0:0] f512_wen;
  logic [31:0] f512_wdata;
  logic [0:0] f512_clk;
  logic [0:0] f512_rst;
  logic [31:0] f512_rdata;
  sr_buffer_32_1 f512(.wen(f512_wen), .wdata(f512_wdata), .clk(f512_clk), .rst(f512_rst), .rdata(f512_rdata));
  assign f512_clk = clk;
  assign f512_rst = rst;
  // Bindings to f512

  // f514
  logic [0:0] f514_wen;
  logic [31:0] f514_wdata;
  logic [0:0] f514_clk;
  logic [0:0] f514_rst;
  logic [31:0] f514_rdata;
  sr_buffer_32_1 f514(.wen(f514_wen), .wdata(f514_wdata), .clk(f514_clk), .rst(f514_rst), .rdata(f514_rdata));
  assign f514_clk = clk;
  assign f514_rst = rst;
  // Bindings to f514

  // f516
  logic [0:0] f516_wen;
  logic [31:0] f516_wdata;
  logic [0:0] f516_clk;
  logic [0:0] f516_rst;
  logic [31:0] f516_rdata;
  sr_buffer_32_1 f516(.wen(f516_wen), .wdata(f516_wdata), .clk(f516_clk), .rst(f516_rst), .rdata(f516_rdata));
  assign f516_clk = clk;
  assign f516_rst = rst;
  // Bindings to f516

  // f518
  logic [0:0] f518_wen;
  logic [31:0] f518_wdata;
  logic [0:0] f518_clk;
  logic [0:0] f518_rst;
  logic [31:0] f518_rdata;
  sr_buffer_32_1 f518(.wen(f518_wen), .wdata(f518_wdata), .clk(f518_clk), .rst(f518_rst), .rdata(f518_rdata));
  assign f518_clk = clk;
  assign f518_rst = rst;
  // Bindings to f518

  // f520
  logic [0:0] f520_wen;
  logic [31:0] f520_wdata;
  logic [0:0] f520_clk;
  logic [0:0] f520_rst;
  logic [31:0] f520_rdata;
  sr_buffer_32_1 f520(.wen(f520_wen), .wdata(f520_wdata), .clk(f520_clk), .rst(f520_rst), .rdata(f520_rdata));
  assign f520_clk = clk;
  assign f520_rst = rst;
  // Bindings to f520

  // f522
  logic [0:0] f522_wen;
  logic [31:0] f522_wdata;
  logic [0:0] f522_clk;
  logic [0:0] f522_rst;
  logic [31:0] f522_rdata;
  sr_buffer_32_1 f522(.wen(f522_wen), .wdata(f522_wdata), .clk(f522_clk), .rst(f522_rst), .rdata(f522_rdata));
  assign f522_clk = clk;
  assign f522_rst = rst;
  // Bindings to f522

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f314
  logic [0:0] f314_wen;
  logic [31:0] f314_wdata;
  logic [0:0] f314_clk;
  logic [0:0] f314_rst;
  logic [31:0] f314_rdata;
  sr_buffer_32_1 f314(.wen(f314_wen), .wdata(f314_wdata), .clk(f314_clk), .rst(f314_rst), .rdata(f314_rdata));
  assign f314_clk = clk;
  assign f314_rst = rst;
  // Bindings to f314

  // f316
  logic [0:0] f316_wen;
  logic [31:0] f316_wdata;
  logic [0:0] f316_clk;
  logic [0:0] f316_rst;
  logic [31:0] f316_rdata;
  sr_buffer_32_1 f316(.wen(f316_wen), .wdata(f316_wdata), .clk(f316_clk), .rst(f316_rst), .rdata(f316_rdata));
  assign f316_clk = clk;
  assign f316_rst = rst;
  // Bindings to f316

  // f318
  logic [0:0] f318_wen;
  logic [31:0] f318_wdata;
  logic [0:0] f318_clk;
  logic [0:0] f318_rst;
  logic [31:0] f318_rdata;
  sr_buffer_32_1 f318(.wen(f318_wen), .wdata(f318_wdata), .clk(f318_clk), .rst(f318_rst), .rdata(f318_rdata));
  assign f318_clk = clk;
  assign f318_rst = rst;
  // Bindings to f318

  // f320
  logic [0:0] f320_wen;
  logic [31:0] f320_wdata;
  logic [0:0] f320_clk;
  logic [0:0] f320_rst;
  logic [31:0] f320_rdata;
  sr_buffer_32_1 f320(.wen(f320_wen), .wdata(f320_wdata), .clk(f320_clk), .rst(f320_rst), .rdata(f320_rdata));
  assign f320_clk = clk;
  assign f320_rst = rst;
  // Bindings to f320

  // f322
  logic [0:0] f322_wen;
  logic [31:0] f322_wdata;
  logic [0:0] f322_clk;
  logic [0:0] f322_rst;
  logic [31:0] f322_rdata;
  sr_buffer_32_1 f322(.wen(f322_wen), .wdata(f322_wdata), .clk(f322_clk), .rst(f322_rst), .rdata(f322_rdata));
  assign f322_clk = clk;
  assign f322_rst = rst;
  // Bindings to f322

  // f324
  logic [0:0] f324_wen;
  logic [31:0] f324_wdata;
  logic [0:0] f324_clk;
  logic [0:0] f324_rst;
  logic [31:0] f324_rdata;
  sr_buffer_32_1 f324(.wen(f324_wen), .wdata(f324_wdata), .clk(f324_clk), .rst(f324_rst), .rdata(f324_rdata));
  assign f324_clk = clk;
  assign f324_rst = rst;
  // Bindings to f324

  // f326
  logic [0:0] f326_wen;
  logic [31:0] f326_wdata;
  logic [0:0] f326_clk;
  logic [0:0] f326_rst;
  logic [31:0] f326_rdata;
  sr_buffer_32_1 f326(.wen(f326_wen), .wdata(f326_wdata), .clk(f326_clk), .rst(f326_rst), .rdata(f326_rdata));
  assign f326_clk = clk;
  assign f326_rst = rst;
  // Bindings to f326

  // f328
  logic [0:0] f328_wen;
  logic [31:0] f328_wdata;
  logic [0:0] f328_clk;
  logic [0:0] f328_rst;
  logic [31:0] f328_rdata;
  sr_buffer_32_1 f328(.wen(f328_wen), .wdata(f328_wdata), .clk(f328_clk), .rst(f328_rst), .rdata(f328_rdata));
  assign f328_clk = clk;
  assign f328_rst = rst;
  // Bindings to f328

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f386
  logic [0:0] f386_wen;
  logic [31:0] f386_wdata;
  logic [0:0] f386_clk;
  logic [0:0] f386_rst;
  logic [31:0] f386_rdata;
  sr_buffer_32_1 f386(.wen(f386_wen), .wdata(f386_wdata), .clk(f386_clk), .rst(f386_rst), .rdata(f386_rdata));
  assign f386_clk = clk;
  assign f386_rst = rst;
  // Bindings to f386

  // f388
  logic [0:0] f388_wen;
  logic [31:0] f388_wdata;
  logic [0:0] f388_clk;
  logic [0:0] f388_rst;
  logic [31:0] f388_rdata;
  sr_buffer_32_1 f388(.wen(f388_wen), .wdata(f388_wdata), .clk(f388_clk), .rst(f388_rst), .rdata(f388_rdata));
  assign f388_clk = clk;
  assign f388_rst = rst;
  // Bindings to f388

  // f390
  logic [0:0] f390_wen;
  logic [31:0] f390_wdata;
  logic [0:0] f390_clk;
  logic [0:0] f390_rst;
  logic [31:0] f390_rdata;
  sr_buffer_32_1 f390(.wen(f390_wen), .wdata(f390_wdata), .clk(f390_clk), .rst(f390_rst), .rdata(f390_rdata));
  assign f390_clk = clk;
  assign f390_rst = rst;
  // Bindings to f390

  // f392
  logic [0:0] f392_wen;
  logic [31:0] f392_wdata;
  logic [0:0] f392_clk;
  logic [0:0] f392_rst;
  logic [31:0] f392_rdata;
  sr_buffer_32_1 f392(.wen(f392_wen), .wdata(f392_wdata), .clk(f392_clk), .rst(f392_rst), .rdata(f392_rdata));
  assign f392_clk = clk;
  assign f392_rst = rst;
  // Bindings to f392

  // f394
  logic [0:0] f394_wen;
  logic [31:0] f394_wdata;
  logic [0:0] f394_clk;
  logic [0:0] f394_rst;
  logic [31:0] f394_rdata;
  sr_buffer_32_1 f394(.wen(f394_wen), .wdata(f394_wdata), .clk(f394_clk), .rst(f394_rst), .rdata(f394_rdata));
  assign f394_clk = clk;
  assign f394_rst = rst;
  // Bindings to f394

  // f396
  logic [0:0] f396_wen;
  logic [31:0] f396_wdata;
  logic [0:0] f396_clk;
  logic [0:0] f396_rst;
  logic [31:0] f396_rdata;
  sr_buffer_32_1 f396(.wen(f396_wen), .wdata(f396_wdata), .clk(f396_clk), .rst(f396_rst), .rdata(f396_rdata));
  assign f396_clk = clk;
  assign f396_rst = rst;
  // Bindings to f396

  // f398
  logic [0:0] f398_wen;
  logic [31:0] f398_wdata;
  logic [0:0] f398_clk;
  logic [0:0] f398_rst;
  logic [31:0] f398_rdata;
  sr_buffer_32_1 f398(.wen(f398_wen), .wdata(f398_wdata), .clk(f398_clk), .rst(f398_rst), .rdata(f398_rdata));
  assign f398_clk = clk;
  assign f398_rst = rst;
  // Bindings to f398

  // f400
  logic [0:0] f400_wen;
  logic [31:0] f400_wdata;
  logic [0:0] f400_clk;
  logic [0:0] f400_rst;
  logic [31:0] f400_rdata;
  sr_buffer_32_1 f400(.wen(f400_wen), .wdata(f400_wdata), .clk(f400_clk), .rst(f400_rst), .rdata(f400_rdata));
  assign f400_clk = clk;
  assign f400_rst = rst;
  // Bindings to f400

  // f402
  logic [0:0] f402_wen;
  logic [31:0] f402_wdata;
  logic [0:0] f402_clk;
  logic [0:0] f402_rst;
  logic [31:0] f402_rdata;
  sr_buffer_32_1 f402(.wen(f402_wen), .wdata(f402_wdata), .clk(f402_clk), .rst(f402_rst), .rdata(f402_rdata));
  assign f402_clk = clk;
  assign f402_rst = rst;
  // Bindings to f402

  // f404
  logic [0:0] f404_wen;
  logic [31:0] f404_wdata;
  logic [0:0] f404_clk;
  logic [0:0] f404_rst;
  logic [31:0] f404_rdata;
  sr_buffer_32_1 f404(.wen(f404_wen), .wdata(f404_wdata), .clk(f404_clk), .rst(f404_rst), .rdata(f404_rdata));
  assign f404_clk = clk;
  assign f404_rst = rst;
  // Bindings to f404

  // f406
  logic [0:0] f406_wen;
  logic [31:0] f406_wdata;
  logic [0:0] f406_clk;
  logic [0:0] f406_rst;
  logic [31:0] f406_rdata;
  sr_buffer_32_1 f406(.wen(f406_wen), .wdata(f406_wdata), .clk(f406_clk), .rst(f406_rst), .rdata(f406_rdata));
  assign f406_clk = clk;
  assign f406_rst = rst;
  // Bindings to f406

  // f408
  logic [0:0] f408_wen;
  logic [31:0] f408_wdata;
  logic [0:0] f408_clk;
  logic [0:0] f408_rst;
  logic [31:0] f408_rdata;
  sr_buffer_32_1 f408(.wen(f408_wen), .wdata(f408_wdata), .clk(f408_clk), .rst(f408_rst), .rdata(f408_rdata));
  assign f408_clk = clk;
  assign f408_rst = rst;
  // Bindings to f408

  // f410
  logic [0:0] f410_wen;
  logic [31:0] f410_wdata;
  logic [0:0] f410_clk;
  logic [0:0] f410_rst;
  logic [31:0] f410_rdata;
  sr_buffer_32_1 f410(.wen(f410_wen), .wdata(f410_wdata), .clk(f410_clk), .rst(f410_rst), .rdata(f410_rdata));
  assign f410_clk = clk;
  assign f410_rst = rst;
  // Bindings to f410

  // f412
  logic [0:0] f412_wen;
  logic [31:0] f412_wdata;
  logic [0:0] f412_clk;
  logic [0:0] f412_rst;
  logic [31:0] f412_rdata;
  sr_buffer_32_1 f412(.wen(f412_wen), .wdata(f412_wdata), .clk(f412_clk), .rst(f412_rst), .rdata(f412_rdata));
  assign f412_clk = clk;
  assign f412_rst = rst;
  // Bindings to f412

  // f414
  logic [0:0] f414_wen;
  logic [31:0] f414_wdata;
  logic [0:0] f414_clk;
  logic [0:0] f414_rst;
  logic [31:0] f414_rdata;
  sr_buffer_32_1 f414(.wen(f414_wen), .wdata(f414_wdata), .clk(f414_clk), .rst(f414_rst), .rdata(f414_rdata));
  assign f414_clk = clk;
  assign f414_rst = rst;
  // Bindings to f414

  // f416
  logic [0:0] f416_wen;
  logic [31:0] f416_wdata;
  logic [0:0] f416_clk;
  logic [0:0] f416_rst;
  logic [31:0] f416_rdata;
  sr_buffer_32_1 f416(.wen(f416_wen), .wdata(f416_wdata), .clk(f416_clk), .rst(f416_rst), .rdata(f416_rdata));
  assign f416_clk = clk;
  assign f416_rst = rst;
  // Bindings to f416

  // f418
  logic [0:0] f418_wen;
  logic [31:0] f418_wdata;
  logic [0:0] f418_clk;
  logic [0:0] f418_rst;
  logic [31:0] f418_rdata;
  sr_buffer_32_1 f418(.wen(f418_wen), .wdata(f418_wdata), .clk(f418_clk), .rst(f418_rst), .rdata(f418_rdata));
  assign f418_clk = clk;
  assign f418_rst = rst;
  // Bindings to f418

  // f420
  logic [0:0] f420_wen;
  logic [31:0] f420_wdata;
  logic [0:0] f420_clk;
  logic [0:0] f420_rst;
  logic [31:0] f420_rdata;
  sr_buffer_32_1 f420(.wen(f420_wen), .wdata(f420_wdata), .clk(f420_clk), .rst(f420_rst), .rdata(f420_rdata));
  assign f420_clk = clk;
  assign f420_rst = rst;
  // Bindings to f420

  // f422
  logic [0:0] f422_wen;
  logic [31:0] f422_wdata;
  logic [0:0] f422_clk;
  logic [0:0] f422_rst;
  logic [31:0] f422_rdata;
  sr_buffer_32_1 f422(.wen(f422_wen), .wdata(f422_wdata), .clk(f422_clk), .rst(f422_rst), .rdata(f422_rdata));
  assign f422_clk = clk;
  assign f422_rst = rst;
  // Bindings to f422

  // f424
  logic [0:0] f424_wen;
  logic [31:0] f424_wdata;
  logic [0:0] f424_clk;
  logic [0:0] f424_rst;
  logic [31:0] f424_rdata;
  sr_buffer_32_1 f424(.wen(f424_wen), .wdata(f424_wdata), .clk(f424_clk), .rst(f424_rst), .rdata(f424_rdata));
  assign f424_clk = clk;
  assign f424_rst = rst;
  // Bindings to f424

  // f426
  logic [0:0] f426_wen;
  logic [31:0] f426_wdata;
  logic [0:0] f426_clk;
  logic [0:0] f426_rst;
  logic [31:0] f426_rdata;
  sr_buffer_32_1 f426(.wen(f426_wen), .wdata(f426_wdata), .clk(f426_clk), .rst(f426_rst), .rdata(f426_rdata));
  assign f426_clk = clk;
  assign f426_rst = rst;
  // Bindings to f426

  // f428
  logic [0:0] f428_wen;
  logic [31:0] f428_wdata;
  logic [0:0] f428_clk;
  logic [0:0] f428_rst;
  logic [31:0] f428_rdata;
  sr_buffer_32_1 f428(.wen(f428_wen), .wdata(f428_wdata), .clk(f428_clk), .rst(f428_rst), .rdata(f428_rdata));
  assign f428_clk = clk;
  assign f428_rst = rst;
  // Bindings to f428

  // f430
  logic [0:0] f430_wen;
  logic [31:0] f430_wdata;
  logic [0:0] f430_clk;
  logic [0:0] f430_rst;
  logic [31:0] f430_rdata;
  sr_buffer_32_1 f430(.wen(f430_wen), .wdata(f430_wdata), .clk(f430_clk), .rst(f430_rst), .rdata(f430_rdata));
  assign f430_clk = clk;
  assign f430_rst = rst;
  // Bindings to f430

  // f432
  logic [0:0] f432_wen;
  logic [31:0] f432_wdata;
  logic [0:0] f432_clk;
  logic [0:0] f432_rst;
  logic [31:0] f432_rdata;
  sr_buffer_32_1 f432(.wen(f432_wen), .wdata(f432_wdata), .clk(f432_clk), .rst(f432_rst), .rdata(f432_rdata));
  assign f432_clk = clk;
  assign f432_rst = rst;
  // Bindings to f432

  // f434
  logic [0:0] f434_wen;
  logic [31:0] f434_wdata;
  logic [0:0] f434_clk;
  logic [0:0] f434_rst;
  logic [31:0] f434_rdata;
  sr_buffer_32_1 f434(.wen(f434_wen), .wdata(f434_wdata), .clk(f434_clk), .rst(f434_rst), .rdata(f434_rdata));
  assign f434_clk = clk;
  assign f434_rst = rst;
  // Bindings to f434

  // f436
  logic [0:0] f436_wen;
  logic [31:0] f436_wdata;
  logic [0:0] f436_clk;
  logic [0:0] f436_rst;
  logic [31:0] f436_rdata;
  sr_buffer_32_1 f436(.wen(f436_wen), .wdata(f436_wdata), .clk(f436_clk), .rst(f436_rst), .rdata(f436_rdata));
  assign f436_clk = clk;
  assign f436_rst = rst;
  // Bindings to f436

  // f438
  logic [0:0] f438_wen;
  logic [31:0] f438_wdata;
  logic [0:0] f438_clk;
  logic [0:0] f438_rst;
  logic [31:0] f438_rdata;
  sr_buffer_32_1 f438(.wen(f438_wen), .wdata(f438_wdata), .clk(f438_clk), .rst(f438_rst), .rdata(f438_rdata));
  assign f438_clk = clk;
  assign f438_rst = rst;
  // Bindings to f438

  // f440
  logic [0:0] f440_wen;
  logic [31:0] f440_wdata;
  logic [0:0] f440_clk;
  logic [0:0] f440_rst;
  logic [31:0] f440_rdata;
  sr_buffer_32_1 f440(.wen(f440_wen), .wdata(f440_wdata), .clk(f440_clk), .rst(f440_rst), .rdata(f440_rdata));
  assign f440_clk = clk;
  assign f440_rst = rst;
  // Bindings to f440

  // f442
  logic [0:0] f442_wen;
  logic [31:0] f442_wdata;
  logic [0:0] f442_clk;
  logic [0:0] f442_rst;
  logic [31:0] f442_rdata;
  sr_buffer_32_1 f442(.wen(f442_wen), .wdata(f442_wdata), .clk(f442_clk), .rst(f442_rst), .rdata(f442_rdata));
  assign f442_clk = clk;
  assign f442_rst = rst;
  // Bindings to f442

  // f444
  logic [0:0] f444_wen;
  logic [31:0] f444_wdata;
  logic [0:0] f444_clk;
  logic [0:0] f444_rst;
  logic [31:0] f444_rdata;
  sr_buffer_32_1 f444(.wen(f444_wen), .wdata(f444_wdata), .clk(f444_clk), .rst(f444_rst), .rdata(f444_rdata));
  assign f444_clk = clk;
  assign f444_rst = rst;
  // Bindings to f444

  // f446
  logic [0:0] f446_wen;
  logic [31:0] f446_wdata;
  logic [0:0] f446_clk;
  logic [0:0] f446_rst;
  logic [31:0] f446_rdata;
  sr_buffer_32_1 f446(.wen(f446_wen), .wdata(f446_wdata), .clk(f446_clk), .rst(f446_rst), .rdata(f446_rdata));
  assign f446_clk = clk;
  assign f446_rst = rst;
  // Bindings to f446

  // f448
  logic [0:0] f448_wen;
  logic [31:0] f448_wdata;
  logic [0:0] f448_clk;
  logic [0:0] f448_rst;
  logic [31:0] f448_rdata;
  sr_buffer_32_1 f448(.wen(f448_wen), .wdata(f448_wdata), .clk(f448_clk), .rst(f448_rst), .rdata(f448_rdata));
  assign f448_clk = clk;
  assign f448_rst = rst;
  // Bindings to f448

  // f450
  logic [0:0] f450_wen;
  logic [31:0] f450_wdata;
  logic [0:0] f450_clk;
  logic [0:0] f450_rst;
  logic [31:0] f450_rdata;
  sr_buffer_32_1 f450(.wen(f450_wen), .wdata(f450_wdata), .clk(f450_clk), .rst(f450_rst), .rdata(f450_rdata));
  assign f450_clk = clk;
  assign f450_rst = rst;
  // Bindings to f450

  // f452
  logic [0:0] f452_wen;
  logic [31:0] f452_wdata;
  logic [0:0] f452_clk;
  logic [0:0] f452_rst;
  logic [31:0] f452_rdata;
  sr_buffer_32_1 f452(.wen(f452_wen), .wdata(f452_wdata), .clk(f452_clk), .rst(f452_rst), .rdata(f452_rdata));
  assign f452_clk = clk;
  assign f452_rst = rst;
  // Bindings to f452

  // f454
  logic [0:0] f454_wen;
  logic [31:0] f454_wdata;
  logic [0:0] f454_clk;
  logic [0:0] f454_rst;
  logic [31:0] f454_rdata;
  sr_buffer_32_1 f454(.wen(f454_wen), .wdata(f454_wdata), .clk(f454_clk), .rst(f454_rst), .rdata(f454_rdata));
  assign f454_clk = clk;
  assign f454_rst = rst;
  // Bindings to f454

  // f456
  logic [0:0] f456_wen;
  logic [31:0] f456_wdata;
  logic [0:0] f456_clk;
  logic [0:0] f456_rst;
  logic [31:0] f456_rdata;
  sr_buffer_32_1 f456(.wen(f456_wen), .wdata(f456_wdata), .clk(f456_clk), .rst(f456_rst), .rdata(f456_rdata));
  assign f456_clk = clk;
  assign f456_rst = rst;
  // Bindings to f456

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f488
  logic [0:0] f488_wen;
  logic [31:0] f488_wdata;
  logic [0:0] f488_clk;
  logic [0:0] f488_rst;
  logic [31:0] f488_rdata;
  sr_buffer_32_1 f488(.wen(f488_wen), .wdata(f488_wdata), .clk(f488_clk), .rst(f488_rst), .rdata(f488_rdata));
  assign f488_clk = clk;
  assign f488_rst = rst;
  // Bindings to f488

  // f490
  logic [0:0] f490_wen;
  logic [31:0] f490_wdata;
  logic [0:0] f490_clk;
  logic [0:0] f490_rst;
  logic [31:0] f490_rdata;
  sr_buffer_32_1 f490(.wen(f490_wen), .wdata(f490_wdata), .clk(f490_clk), .rst(f490_rst), .rdata(f490_rdata));
  assign f490_clk = clk;
  assign f490_rst = rst;
  // Bindings to f490

  // f492
  logic [0:0] f492_wen;
  logic [31:0] f492_wdata;
  logic [0:0] f492_clk;
  logic [0:0] f492_rst;
  logic [31:0] f492_rdata;
  sr_buffer_32_1 f492(.wen(f492_wen), .wdata(f492_wdata), .clk(f492_clk), .rst(f492_rst), .rdata(f492_rdata));
  assign f492_clk = clk;
  assign f492_rst = rst;
  // Bindings to f492

  // f494
  logic [0:0] f494_wen;
  logic [31:0] f494_wdata;
  logic [0:0] f494_clk;
  logic [0:0] f494_rst;
  logic [31:0] f494_rdata;
  sr_buffer_32_1 f494(.wen(f494_wen), .wdata(f494_wdata), .clk(f494_clk), .rst(f494_rst), .rdata(f494_rdata));
  assign f494_clk = clk;
  assign f494_rst = rst;
  // Bindings to f494

  // f496
  logic [0:0] f496_wen;
  logic [31:0] f496_wdata;
  logic [0:0] f496_clk;
  logic [0:0] f496_rst;
  logic [31:0] f496_rdata;
  sr_buffer_32_1 f496(.wen(f496_wen), .wdata(f496_wdata), .clk(f496_clk), .rst(f496_rst), .rdata(f496_rdata));
  assign f496_clk = clk;
  assign f496_rst = rst;
  // Bindings to f496

  // f498
  logic [0:0] f498_wen;
  logic [31:0] f498_wdata;
  logic [0:0] f498_clk;
  logic [0:0] f498_rst;
  logic [31:0] f498_rdata;
  sr_buffer_32_1 f498(.wen(f498_wen), .wdata(f498_wdata), .clk(f498_clk), .rst(f498_rst), .rdata(f498_rdata));
  assign f498_clk = clk;
  assign f498_rst = rst;
  // Bindings to f498

  // f500
  logic [0:0] f500_wen;
  logic [31:0] f500_wdata;
  logic [0:0] f500_clk;
  logic [0:0] f500_rst;
  logic [31:0] f500_rdata;
  sr_buffer_32_1 f500(.wen(f500_wen), .wdata(f500_wdata), .clk(f500_clk), .rst(f500_rst), .rdata(f500_rdata));
  assign f500_clk = clk;
  assign f500_rst = rst;
  // Bindings to f500

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f346
  logic [0:0] f346_wen;
  logic [31:0] f346_wdata;
  logic [0:0] f346_clk;
  logic [0:0] f346_rst;
  logic [31:0] f346_rdata;
  sr_buffer_32_1 f346(.wen(f346_wen), .wdata(f346_wdata), .clk(f346_clk), .rst(f346_rst), .rdata(f346_rdata));
  assign f346_clk = clk;
  assign f346_rst = rst;
  // Bindings to f346

  // f348
  logic [0:0] f348_wen;
  logic [31:0] f348_wdata;
  logic [0:0] f348_clk;
  logic [0:0] f348_rst;
  logic [31:0] f348_rdata;
  sr_buffer_32_1 f348(.wen(f348_wen), .wdata(f348_wdata), .clk(f348_clk), .rst(f348_rst), .rdata(f348_rdata));
  assign f348_clk = clk;
  assign f348_rst = rst;
  // Bindings to f348

  // f350
  logic [0:0] f350_wen;
  logic [31:0] f350_wdata;
  logic [0:0] f350_clk;
  logic [0:0] f350_rst;
  logic [31:0] f350_rdata;
  sr_buffer_32_1 f350(.wen(f350_wen), .wdata(f350_wdata), .clk(f350_clk), .rst(f350_rst), .rdata(f350_rdata));
  assign f350_clk = clk;
  assign f350_rst = rst;
  // Bindings to f350

  // f352
  logic [0:0] f352_wen;
  logic [31:0] f352_wdata;
  logic [0:0] f352_clk;
  logic [0:0] f352_rst;
  logic [31:0] f352_rdata;
  sr_buffer_32_1 f352(.wen(f352_wen), .wdata(f352_wdata), .clk(f352_clk), .rst(f352_rst), .rdata(f352_rdata));
  assign f352_clk = clk;
  assign f352_rst = rst;
  // Bindings to f352

  // f354
  logic [0:0] f354_wen;
  logic [31:0] f354_wdata;
  logic [0:0] f354_clk;
  logic [0:0] f354_rst;
  logic [31:0] f354_rdata;
  sr_buffer_32_1 f354(.wen(f354_wen), .wdata(f354_wdata), .clk(f354_clk), .rst(f354_rst), .rdata(f354_rdata));
  assign f354_clk = clk;
  assign f354_rst = rst;
  // Bindings to f354

  // f356
  logic [0:0] f356_wen;
  logic [31:0] f356_wdata;
  logic [0:0] f356_clk;
  logic [0:0] f356_rst;
  logic [31:0] f356_rdata;
  sr_buffer_32_1 f356(.wen(f356_wen), .wdata(f356_wdata), .clk(f356_clk), .rst(f356_rst), .rdata(f356_rdata));
  assign f356_clk = clk;
  assign f356_rst = rst;
  // Bindings to f356

  // f358
  logic [0:0] f358_wen;
  logic [31:0] f358_wdata;
  logic [0:0] f358_clk;
  logic [0:0] f358_rst;
  logic [31:0] f358_rdata;
  sr_buffer_32_1 f358(.wen(f358_wen), .wdata(f358_wdata), .clk(f358_clk), .rst(f358_rst), .rdata(f358_rdata));
  assign f358_clk = clk;
  assign f358_rst = rst;
  // Bindings to f358

  // f360
  logic [0:0] f360_wen;
  logic [31:0] f360_wdata;
  logic [0:0] f360_clk;
  logic [0:0] f360_rst;
  logic [31:0] f360_rdata;
  sr_buffer_32_1 f360(.wen(f360_wen), .wdata(f360_wdata), .clk(f360_clk), .rst(f360_rst), .rdata(f360_rdata));
  assign f360_clk = clk;
  assign f360_rst = rst;
  // Bindings to f360

  // f362
  logic [0:0] f362_wen;
  logic [31:0] f362_wdata;
  logic [0:0] f362_clk;
  logic [0:0] f362_rst;
  logic [31:0] f362_rdata;
  sr_buffer_32_1 f362(.wen(f362_wen), .wdata(f362_wdata), .clk(f362_clk), .rst(f362_rst), .rdata(f362_rdata));
  assign f362_clk = clk;
  assign f362_rst = rst;
  // Bindings to f362

  // f364
  logic [0:0] f364_wen;
  logic [31:0] f364_wdata;
  logic [0:0] f364_clk;
  logic [0:0] f364_rst;
  logic [31:0] f364_rdata;
  sr_buffer_32_1 f364(.wen(f364_wen), .wdata(f364_wdata), .clk(f364_clk), .rst(f364_rst), .rdata(f364_rdata));
  assign f364_clk = clk;
  assign f364_rst = rst;
  // Bindings to f364

  // f366
  logic [0:0] f366_wen;
  logic [31:0] f366_wdata;
  logic [0:0] f366_clk;
  logic [0:0] f366_rst;
  logic [31:0] f366_rdata;
  sr_buffer_32_1 f366(.wen(f366_wen), .wdata(f366_wdata), .clk(f366_clk), .rst(f366_rst), .rdata(f366_rdata));
  assign f366_clk = clk;
  assign f366_rst = rst;
  // Bindings to f366

  // f368
  logic [0:0] f368_wen;
  logic [31:0] f368_wdata;
  logic [0:0] f368_clk;
  logic [0:0] f368_rst;
  logic [31:0] f368_rdata;
  sr_buffer_32_1 f368(.wen(f368_wen), .wdata(f368_wdata), .clk(f368_clk), .rst(f368_rst), .rdata(f368_rdata));
  assign f368_clk = clk;
  assign f368_rst = rst;
  // Bindings to f368

  // f370
  logic [0:0] f370_wen;
  logic [31:0] f370_wdata;
  logic [0:0] f370_clk;
  logic [0:0] f370_rst;
  logic [31:0] f370_rdata;
  sr_buffer_32_1 f370(.wen(f370_wen), .wdata(f370_wdata), .clk(f370_clk), .rst(f370_rst), .rdata(f370_rdata));
  assign f370_clk = clk;
  assign f370_rst = rst;
  // Bindings to f370

  // f372
  logic [0:0] f372_wen;
  logic [31:0] f372_wdata;
  logic [0:0] f372_clk;
  logic [0:0] f372_rst;
  logic [31:0] f372_rdata;
  sr_buffer_32_1 f372(.wen(f372_wen), .wdata(f372_wdata), .clk(f372_clk), .rst(f372_rst), .rdata(f372_rdata));
  assign f372_clk = clk;
  assign f372_rst = rst;
  // Bindings to f372

  // f374
  logic [0:0] f374_wen;
  logic [31:0] f374_wdata;
  logic [0:0] f374_clk;
  logic [0:0] f374_rst;
  logic [31:0] f374_rdata;
  sr_buffer_32_1 f374(.wen(f374_wen), .wdata(f374_wdata), .clk(f374_clk), .rst(f374_rst), .rdata(f374_rdata));
  assign f374_clk = clk;
  assign f374_rst = rst;
  // Bindings to f374

  // f376
  logic [0:0] f376_wen;
  logic [31:0] f376_wdata;
  logic [0:0] f376_clk;
  logic [0:0] f376_rst;
  logic [31:0] f376_rdata;
  sr_buffer_32_1 f376(.wen(f376_wen), .wdata(f376_wdata), .clk(f376_clk), .rst(f376_rst), .rdata(f376_rdata));
  assign f376_clk = clk;
  assign f376_rst = rst;
  // Bindings to f376

  // f378
  logic [0:0] f378_wen;
  logic [31:0] f378_wdata;
  logic [0:0] f378_clk;
  logic [0:0] f378_rst;
  logic [31:0] f378_rdata;
  sr_buffer_32_1 f378(.wen(f378_wen), .wdata(f378_wdata), .clk(f378_clk), .rst(f378_rst), .rdata(f378_rdata));
  assign f378_clk = clk;
  assign f378_rst = rst;
  // Bindings to f378

  // f380
  logic [0:0] f380_wen;
  logic [31:0] f380_wdata;
  logic [0:0] f380_clk;
  logic [0:0] f380_rst;
  logic [31:0] f380_rdata;
  sr_buffer_32_1 f380(.wen(f380_wen), .wdata(f380_wdata), .clk(f380_clk), .rst(f380_rst), .rdata(f380_rdata));
  assign f380_clk = clk;
  assign f380_rst = rst;
  // Bindings to f380

  // f382
  logic [0:0] f382_wen;
  logic [31:0] f382_wdata;
  logic [0:0] f382_clk;
  logic [0:0] f382_rst;
  logic [31:0] f382_rdata;
  sr_buffer_32_1 f382(.wen(f382_wen), .wdata(f382_wdata), .clk(f382_clk), .rst(f382_rst), .rdata(f382_rdata));
  assign f382_clk = clk;
  assign f382_rst = rst;
  // Bindings to f382

  // f384
  logic [0:0] f384_wen;
  logic [31:0] f384_wdata;
  logic [0:0] f384_clk;
  logic [0:0] f384_rst;
  logic [31:0] f384_rdata;
  sr_buffer_32_1 f384(.wen(f384_wen), .wdata(f384_wdata), .clk(f384_clk), .rst(f384_rst), .rdata(f384_rdata));
  assign f384_clk = clk;
  assign f384_rst = rst;
  // Bindings to f384

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f330
  logic [0:0] f330_wen;
  logic [31:0] f330_wdata;
  logic [0:0] f330_clk;
  logic [0:0] f330_rst;
  logic [31:0] f330_rdata;
  sr_buffer_32_1 f330(.wen(f330_wen), .wdata(f330_wdata), .clk(f330_clk), .rst(f330_rst), .rdata(f330_rdata));
  assign f330_clk = clk;
  assign f330_rst = rst;
  // Bindings to f330

  // f332
  logic [0:0] f332_wen;
  logic [31:0] f332_wdata;
  logic [0:0] f332_clk;
  logic [0:0] f332_rst;
  logic [31:0] f332_rdata;
  sr_buffer_32_1 f332(.wen(f332_wen), .wdata(f332_wdata), .clk(f332_clk), .rst(f332_rst), .rdata(f332_rdata));
  assign f332_clk = clk;
  assign f332_rst = rst;
  // Bindings to f332

  // f334
  logic [0:0] f334_wen;
  logic [31:0] f334_wdata;
  logic [0:0] f334_clk;
  logic [0:0] f334_rst;
  logic [31:0] f334_rdata;
  sr_buffer_32_1 f334(.wen(f334_wen), .wdata(f334_wdata), .clk(f334_clk), .rst(f334_rst), .rdata(f334_rdata));
  assign f334_clk = clk;
  assign f334_rst = rst;
  // Bindings to f334

  // f336
  logic [0:0] f336_wen;
  logic [31:0] f336_wdata;
  logic [0:0] f336_clk;
  logic [0:0] f336_rst;
  logic [31:0] f336_rdata;
  sr_buffer_32_1 f336(.wen(f336_wen), .wdata(f336_wdata), .clk(f336_clk), .rst(f336_rst), .rdata(f336_rdata));
  assign f336_clk = clk;
  assign f336_rst = rst;
  // Bindings to f336

  // f338
  logic [0:0] f338_wen;
  logic [31:0] f338_wdata;
  logic [0:0] f338_clk;
  logic [0:0] f338_rst;
  logic [31:0] f338_rdata;
  sr_buffer_32_1 f338(.wen(f338_wen), .wdata(f338_wdata), .clk(f338_clk), .rst(f338_rst), .rdata(f338_rdata));
  assign f338_clk = clk;
  assign f338_rst = rst;
  // Bindings to f338

  // f340
  logic [0:0] f340_wen;
  logic [31:0] f340_wdata;
  logic [0:0] f340_clk;
  logic [0:0] f340_rst;
  logic [31:0] f340_rdata;
  sr_buffer_32_1 f340(.wen(f340_wen), .wdata(f340_wdata), .clk(f340_clk), .rst(f340_rst), .rdata(f340_rdata));
  assign f340_clk = clk;
  assign f340_rst = rst;
  // Bindings to f340

  // f342
  logic [0:0] f342_wen;
  logic [31:0] f342_wdata;
  logic [0:0] f342_clk;
  logic [0:0] f342_rst;
  logic [31:0] f342_rdata;
  sr_buffer_32_1 f342(.wen(f342_wen), .wdata(f342_wdata), .clk(f342_clk), .rst(f342_rst), .rdata(f342_rdata));
  assign f342_clk = clk;
  assign f342_rst = rst;
  // Bindings to f342

  // f344
  logic [0:0] f344_wen;
  logic [31:0] f344_wdata;
  logic [0:0] f344_clk;
  logic [0:0] f344_rst;
  logic [31:0] f344_rdata;
  sr_buffer_32_1 f344(.wen(f344_wen), .wdata(f344_wdata), .clk(f344_clk), .rst(f344_rst), .rdata(f344_rdata));
  assign f344_clk = clk;
  assign f344_rst = rst;
  // Bindings to f344

  // f524
  logic [0:0] f524_wen;
  logic [31:0] f524_wdata;
  logic [0:0] f524_clk;
  logic [0:0] f524_rst;
  logic [31:0] f524_rdata;
  sr_buffer_32_1 f524(.wen(f524_wen), .wdata(f524_wdata), .clk(f524_clk), .rst(f524_rst), .rdata(f524_rdata));
  assign f524_clk = clk;
  assign f524_rst = rst;
  // Bindings to f524

  // f526
  logic [0:0] f526_wen;
  logic [31:0] f526_wdata;
  logic [0:0] f526_clk;
  logic [0:0] f526_rst;
  logic [31:0] f526_rdata;
  sr_buffer_32_1 f526(.wen(f526_wen), .wdata(f526_wdata), .clk(f526_clk), .rst(f526_rst), .rdata(f526_rdata));
  assign f526_clk = clk;
  assign f526_rst = rst;
  // Bindings to f526

  // f528
  logic [0:0] f528_wen;
  logic [31:0] f528_wdata;
  logic [0:0] f528_clk;
  logic [0:0] f528_rst;
  logic [31:0] f528_rdata;
  sr_buffer_32_1 f528(.wen(f528_wen), .wdata(f528_wdata), .clk(f528_clk), .rst(f528_rst), .rdata(f528_rdata));
  assign f528_clk = clk;
  assign f528_rst = rst;
  // Bindings to f528

  // f530
  logic [0:0] f530_wen;
  logic [31:0] f530_wdata;
  logic [0:0] f530_clk;
  logic [0:0] f530_rst;
  logic [31:0] f530_rdata;
  sr_buffer_32_1 f530(.wen(f530_wen), .wdata(f530_wdata), .clk(f530_clk), .rst(f530_rst), .rdata(f530_rdata));
  assign f530_clk = clk;
  assign f530_rst = rst;
  // Bindings to f530

  // f532
  logic [0:0] f532_wen;
  logic [31:0] f532_wdata;
  logic [0:0] f532_clk;
  logic [0:0] f532_rst;
  logic [31:0] f532_rdata;
  sr_buffer_32_1 f532(.wen(f532_wen), .wdata(f532_wdata), .clk(f532_clk), .rst(f532_rst), .rdata(f532_rdata));
  assign f532_clk = clk;
  assign f532_rst = rst;
  // Bindings to f532

  // f534
  logic [0:0] f534_wen;
  logic [31:0] f534_wdata;
  logic [0:0] f534_clk;
  logic [0:0] f534_rst;
  logic [31:0] f534_rdata;
  sr_buffer_32_1 f534(.wen(f534_wen), .wdata(f534_wdata), .clk(f534_clk), .rst(f534_rst), .rdata(f534_rdata));
  assign f534_clk = clk;
  assign f534_rst = rst;
  // Bindings to f534

  // f536
  logic [0:0] f536_wen;
  logic [31:0] f536_wdata;
  logic [0:0] f536_clk;
  logic [0:0] f536_rst;
  logic [31:0] f536_rdata;
  sr_buffer_32_1 f536(.wen(f536_wen), .wdata(f536_wdata), .clk(f536_clk), .rst(f536_rst), .rdata(f536_rdata));
  assign f536_clk = clk;
  assign f536_rst = rst;
  // Bindings to f536

  // f538
  logic [0:0] f538_wen;
  logic [31:0] f538_wdata;
  logic [0:0] f538_clk;
  logic [0:0] f538_rst;
  logic [31:0] f538_rdata;
  sr_buffer_32_1 f538(.wen(f538_wen), .wdata(f538_wdata), .clk(f538_clk), .rst(f538_rst), .rdata(f538_rdata));
  assign f538_clk = clk;
  assign f538_rst = rst;
  // Bindings to f538

  // f540
  logic [0:0] f540_wen;
  logic [31:0] f540_wdata;
  logic [0:0] f540_clk;
  logic [0:0] f540_rst;
  logic [31:0] f540_rdata;
  sr_buffer_32_1 f540(.wen(f540_wen), .wdata(f540_wdata), .clk(f540_clk), .rst(f540_rst), .rdata(f540_rdata));
  assign f540_clk = clk;
  assign f540_rst = rst;
  // Bindings to f540

  // f542
  logic [0:0] f542_wen;
  logic [31:0] f542_wdata;
  logic [0:0] f542_clk;
  logic [0:0] f542_rst;
  logic [31:0] f542_rdata;
  sr_buffer_32_1 f542(.wen(f542_wen), .wdata(f542_wdata), .clk(f542_clk), .rst(f542_rst), .rdata(f542_rdata));
  assign f542_clk = clk;
  assign f542_rst = rst;
  // Bindings to f542

  // f544
  logic [0:0] f544_wen;
  logic [31:0] f544_wdata;
  logic [0:0] f544_clk;
  logic [0:0] f544_rst;
  logic [31:0] f544_rdata;
  sr_buffer_32_1 f544(.wen(f544_wen), .wdata(f544_wdata), .clk(f544_clk), .rst(f544_rst), .rdata(f544_rdata));
  assign f544_clk = clk;
  assign f544_rst = rst;
  // Bindings to f544

  // f546
  logic [0:0] f546_wen;
  logic [31:0] f546_wdata;
  logic [0:0] f546_clk;
  logic [0:0] f546_rst;
  logic [31:0] f546_rdata;
  sr_buffer_32_1 f546(.wen(f546_wen), .wdata(f546_wdata), .clk(f546_clk), .rst(f546_rst), .rdata(f546_rdata));
  assign f546_clk = clk;
  assign f546_rst = rst;
  // Bindings to f546

  // f548
  logic [0:0] f548_wen;
  logic [31:0] f548_wdata;
  logic [0:0] f548_clk;
  logic [0:0] f548_rst;
  logic [31:0] f548_rdata;
  sr_buffer_32_1 f548(.wen(f548_wen), .wdata(f548_wdata), .clk(f548_clk), .rst(f548_rst), .rdata(f548_rdata));
  assign f548_clk = clk;
  assign f548_rst = rst;
  // Bindings to f548

  // f550
  logic [0:0] f550_wen;
  logic [31:0] f550_wdata;
  logic [0:0] f550_clk;
  logic [0:0] f550_rst;
  logic [31:0] f550_rdata;
  sr_buffer_32_1 f550(.wen(f550_wen), .wdata(f550_wdata), .clk(f550_clk), .rst(f550_rst), .rdata(f550_rdata));
  assign f550_clk = clk;
  assign f550_rst = rst;
  // Bindings to f550

  // f552
  logic [0:0] f552_wen;
  logic [31:0] f552_wdata;
  logic [0:0] f552_clk;
  logic [0:0] f552_rst;
  logic [31:0] f552_rdata;
  sr_buffer_32_1 f552(.wen(f552_wen), .wdata(f552_wdata), .clk(f552_clk), .rst(f552_rst), .rdata(f552_rdata));
  assign f552_clk = clk;
  assign f552_rst = rst;
  // Bindings to f552

  // f554
  logic [0:0] f554_wen;
  logic [31:0] f554_wdata;
  logic [0:0] f554_clk;
  logic [0:0] f554_rst;
  logic [31:0] f554_rdata;
  sr_buffer_32_1 f554(.wen(f554_wen), .wdata(f554_wdata), .clk(f554_clk), .rst(f554_rst), .rdata(f554_rdata));
  assign f554_clk = clk;
  assign f554_rst = rst;
  // Bindings to f554

  // f556
  logic [0:0] f556_wen;
  logic [31:0] f556_wdata;
  logic [0:0] f556_clk;
  logic [0:0] f556_rst;
  logic [31:0] f556_rdata;
  sr_buffer_32_1 f556(.wen(f556_wen), .wdata(f556_wdata), .clk(f556_clk), .rst(f556_rst), .rdata(f556_rdata));
  assign f556_clk = clk;
  assign f556_rst = rst;
  // Bindings to f556

  // f558
  logic [0:0] f558_wen;
  logic [31:0] f558_wdata;
  logic [0:0] f558_clk;
  logic [0:0] f558_rst;
  logic [31:0] f558_rdata;
  sr_buffer_32_1 f558(.wen(f558_wen), .wdata(f558_wdata), .clk(f558_clk), .rst(f558_rst), .rdata(f558_rdata));
  assign f558_clk = clk;
  assign f558_rst = rst;
  // Bindings to f558

  // f560
  logic [0:0] f560_wen;
  logic [31:0] f560_wdata;
  logic [0:0] f560_clk;
  logic [0:0] f560_rst;
  logic [31:0] f560_rdata;
  sr_buffer_32_1 f560(.wen(f560_wen), .wdata(f560_wdata), .clk(f560_clk), .rst(f560_rst), .rdata(f560_rdata));
  assign f560_clk = clk;
  assign f560_rst = rst;
  // Bindings to f560

  // f562
  logic [0:0] f562_wen;
  logic [31:0] f562_wdata;
  logic [0:0] f562_clk;
  logic [0:0] f562_rst;
  logic [31:0] f562_rdata;
  sr_buffer_32_1 f562(.wen(f562_wen), .wdata(f562_wdata), .clk(f562_clk), .rst(f562_rst), .rdata(f562_rdata));
  assign f562_clk = clk;
  assign f562_rst = rst;
  // Bindings to f562

  // f564
  logic [0:0] f564_wen;
  logic [31:0] f564_wdata;
  logic [0:0] f564_clk;
  logic [0:0] f564_rst;
  logic [31:0] f564_rdata;
  sr_buffer_32_1 f564(.wen(f564_wen), .wdata(f564_wdata), .clk(f564_clk), .rst(f564_rst), .rdata(f564_rdata));
  assign f564_clk = clk;
  assign f564_rst = rst;
  // Bindings to f564

  // f566
  logic [0:0] f566_wen;
  logic [31:0] f566_wdata;
  logic [0:0] f566_clk;
  logic [0:0] f566_rst;
  logic [31:0] f566_rdata;
  sr_buffer_32_1 f566(.wen(f566_wen), .wdata(f566_wdata), .clk(f566_clk), .rst(f566_rst), .rdata(f566_rdata));
  assign f566_clk = clk;
  assign f566_rst = rst;
  // Bindings to f566

  // f568
  logic [0:0] f568_wen;
  logic [31:0] f568_wdata;
  logic [0:0] f568_clk;
  logic [0:0] f568_rst;
  logic [31:0] f568_rdata;
  sr_buffer_32_1 f568(.wen(f568_wen), .wdata(f568_wdata), .clk(f568_clk), .rst(f568_rst), .rdata(f568_rdata));
  assign f568_clk = clk;
  assign f568_rst = rst;
  // Bindings to f568

  // f570
  logic [0:0] f570_wen;
  logic [31:0] f570_wdata;
  logic [0:0] f570_clk;
  logic [0:0] f570_rst;
  logic [31:0] f570_rdata;
  sr_buffer_32_1 f570(.wen(f570_wen), .wdata(f570_wdata), .clk(f570_clk), .rst(f570_rst), .rdata(f570_rdata));
  assign f570_clk = clk;
  assign f570_rst = rst;
  // Bindings to f570

  // f572
  logic [0:0] f572_wen;
  logic [31:0] f572_wdata;
  logic [0:0] f572_clk;
  logic [0:0] f572_rst;
  logic [31:0] f572_rdata;
  sr_buffer_32_1 f572(.wen(f572_wen), .wdata(f572_wdata), .clk(f572_clk), .rst(f572_rst), .rdata(f572_rdata));
  assign f572_clk = clk;
  assign f572_rst = rst;
  // Bindings to f572

  // f574
  logic [0:0] f574_wen;
  logic [31:0] f574_wdata;
  logic [0:0] f574_clk;
  logic [0:0] f574_rst;
  logic [31:0] f574_rdata;
  sr_buffer_32_1 f574(.wen(f574_wen), .wdata(f574_wdata), .clk(f574_clk), .rst(f574_rst), .rdata(f574_rdata));
  assign f574_clk = clk;
  assign f574_rst = rst;
  // Bindings to f574

  // f576
  logic [0:0] f576_wen;
  logic [31:0] f576_wdata;
  logic [0:0] f576_clk;
  logic [0:0] f576_rst;
  logic [31:0] f576_rdata;
  sr_buffer_32_1 f576(.wen(f576_wen), .wdata(f576_wdata), .clk(f576_clk), .rst(f576_rst), .rdata(f576_rdata));
  assign f576_clk = clk;
  assign f576_rst = rst;
  // Bindings to f576

  // f578
  logic [0:0] f578_wen;
  logic [31:0] f578_wdata;
  logic [0:0] f578_clk;
  logic [0:0] f578_rst;
  logic [31:0] f578_rdata;
  sr_buffer_32_1 f578(.wen(f578_wen), .wdata(f578_wdata), .clk(f578_clk), .rst(f578_rst), .rdata(f578_rdata));
  assign f578_clk = clk;
  assign f578_rst = rst;
  // Bindings to f578

  // f580
  logic [0:0] f580_wen;
  logic [31:0] f580_wdata;
  logic [0:0] f580_clk;
  logic [0:0] f580_rst;
  logic [31:0] f580_rdata;
  sr_buffer_32_1 f580(.wen(f580_wen), .wdata(f580_wdata), .clk(f580_clk), .rst(f580_rst), .rdata(f580_rdata));
  assign f580_clk = clk;
  assign f580_rst = rst;
  // Bindings to f580

  // f582
  logic [0:0] f582_wen;
  logic [31:0] f582_wdata;
  logic [0:0] f582_clk;
  logic [0:0] f582_rst;
  logic [31:0] f582_rdata;
  sr_buffer_32_1 f582(.wen(f582_wen), .wdata(f582_wdata), .clk(f582_clk), .rst(f582_rst), .rdata(f582_rdata));
  assign f582_clk = clk;
  assign f582_rst = rst;
  // Bindings to f582

  // f584
  logic [0:0] f584_wen;
  logic [31:0] f584_wdata;
  logic [0:0] f584_clk;
  logic [0:0] f584_rst;
  logic [31:0] f584_rdata;
  sr_buffer_32_1 f584(.wen(f584_wen), .wdata(f584_wdata), .clk(f584_clk), .rst(f584_rst), .rdata(f584_rdata));
  assign f584_clk = clk;
  assign f584_rst = rst;
  // Bindings to f584

  // f586
  logic [0:0] f586_wen;
  logic [31:0] f586_wdata;
  logic [0:0] f586_clk;
  logic [0:0] f586_rst;
  logic [31:0] f586_rdata;
  sr_buffer_32_1 f586(.wen(f586_wen), .wdata(f586_wdata), .clk(f586_clk), .rst(f586_rst), .rdata(f586_rdata));
  assign f586_clk = clk;
  assign f586_rst = rst;
  // Bindings to f586

  // f588
  logic [0:0] f588_wen;
  logic [31:0] f588_wdata;
  logic [0:0] f588_clk;
  logic [0:0] f588_rst;
  logic [31:0] f588_rdata;
  sr_buffer_32_1 f588(.wen(f588_wen), .wdata(f588_wdata), .clk(f588_clk), .rst(f588_rst), .rdata(f588_rdata));
  assign f588_clk = clk;
  assign f588_rst = rst;
  // Bindings to f588

  // f590
  logic [0:0] f590_wen;
  logic [31:0] f590_wdata;
  logic [0:0] f590_clk;
  logic [0:0] f590_rst;
  logic [31:0] f590_rdata;
  sr_buffer_32_1 f590(.wen(f590_wen), .wdata(f590_wdata), .clk(f590_clk), .rst(f590_rst), .rdata(f590_rdata));
  assign f590_clk = clk;
  assign f590_rst = rst;
  // Bindings to f590

  // f592
  logic [0:0] f592_wen;
  logic [31:0] f592_wdata;
  logic [0:0] f592_clk;
  logic [0:0] f592_rst;
  logic [31:0] f592_rdata;
  sr_buffer_32_1 f592(.wen(f592_wen), .wdata(f592_wdata), .clk(f592_clk), .rst(f592_rst), .rdata(f592_rdata));
  assign f592_clk = clk;
  assign f592_rst = rst;
  // Bindings to f592

  // f594
  logic [0:0] f594_wen;
  logic [31:0] f594_wdata;
  logic [0:0] f594_clk;
  logic [0:0] f594_rst;
  logic [31:0] f594_rdata;
  sr_buffer_32_1 f594(.wen(f594_wen), .wdata(f594_wdata), .clk(f594_clk), .rst(f594_rst), .rdata(f594_rdata));
  assign f594_clk = clk;
  assign f594_rst = rst;
  // Bindings to f594

  // f596
  logic [0:0] f596_wen;
  logic [31:0] f596_wdata;
  logic [0:0] f596_clk;
  logic [0:0] f596_rst;
  logic [31:0] f596_rdata;
  sr_buffer_32_1 f596(.wen(f596_wen), .wdata(f596_wdata), .clk(f596_clk), .rst(f596_rst), .rdata(f596_rdata));
  assign f596_clk = clk;
  assign f596_rst = rst;
  // Bindings to f596

  // f598
  logic [0:0] f598_wen;
  logic [31:0] f598_wdata;
  logic [0:0] f598_clk;
  logic [0:0] f598_rst;
  logic [31:0] f598_rdata;
  sr_buffer_32_1 f598(.wen(f598_wen), .wdata(f598_wdata), .clk(f598_clk), .rst(f598_rst), .rdata(f598_rdata));
  assign f598_clk = clk;
  assign f598_rst = rst;
  // Bindings to f598

  // f600
  logic [0:0] f600_wen;
  logic [31:0] f600_wdata;
  logic [0:0] f600_clk;
  logic [0:0] f600_rst;
  logic [31:0] f600_rdata;
  sr_buffer_32_1 f600(.wen(f600_wen), .wdata(f600_wdata), .clk(f600_clk), .rst(f600_rst), .rdata(f600_rdata));
  assign f600_clk = clk;
  assign f600_rst = rst;
  // Bindings to f600

  // f602
  logic [0:0] f602_wen;
  logic [31:0] f602_wdata;
  logic [0:0] f602_clk;
  logic [0:0] f602_rst;
  logic [31:0] f602_rdata;
  sr_buffer_32_1 f602(.wen(f602_wen), .wdata(f602_wdata), .clk(f602_clk), .rst(f602_rst), .rdata(f602_rdata));
  assign f602_clk = clk;
  assign f602_rst = rst;
  // Bindings to f602

  // f604
  logic [0:0] f604_wen;
  logic [31:0] f604_wdata;
  logic [0:0] f604_clk;
  logic [0:0] f604_rst;
  logic [31:0] f604_rdata;
  sr_buffer_32_1 f604(.wen(f604_wen), .wdata(f604_wdata), .clk(f604_clk), .rst(f604_rst), .rdata(f604_rdata));
  assign f604_clk = clk;
  assign f604_rst = rst;
  // Bindings to f604

  // f606
  logic [0:0] f606_wen;
  logic [31:0] f606_wdata;
  logic [0:0] f606_clk;
  logic [0:0] f606_rst;
  logic [31:0] f606_rdata;
  sr_buffer_32_1 f606(.wen(f606_wen), .wdata(f606_wdata), .clk(f606_clk), .rst(f606_rst), .rdata(f606_rdata));
  assign f606_clk = clk;
  assign f606_rst = rst;
  // Bindings to f606

  // f608
  logic [0:0] f608_wen;
  logic [31:0] f608_wdata;
  logic [0:0] f608_clk;
  logic [0:0] f608_rst;
  logic [31:0] f608_rdata;
  sr_buffer_32_1 f608(.wen(f608_wen), .wdata(f608_wdata), .clk(f608_clk), .rst(f608_rst), .rdata(f608_rdata));
  assign f608_clk = clk;
  assign f608_rst = rst;
  // Bindings to f608

  // f610
  logic [0:0] f610_wen;
  logic [31:0] f610_wdata;
  logic [0:0] f610_clk;
  logic [0:0] f610_rst;
  logic [31:0] f610_rdata;
  sr_buffer_32_1 f610(.wen(f610_wen), .wdata(f610_wdata), .clk(f610_clk), .rst(f610_rst), .rdata(f610_rdata));
  assign f610_clk = clk;
  assign f610_rst = rst;
  // Bindings to f610

  // f612
  logic [0:0] f612_wen;
  logic [31:0] f612_wdata;
  logic [0:0] f612_clk;
  logic [0:0] f612_rst;
  logic [31:0] f612_rdata;
  sr_buffer_32_1 f612(.wen(f612_wen), .wdata(f612_wdata), .clk(f612_clk), .rst(f612_rst), .rdata(f612_rdata));
  assign f612_clk = clk;
  assign f612_rst = rst;
  // Bindings to f612

  // f614
  logic [0:0] f614_wen;
  logic [31:0] f614_wdata;
  logic [0:0] f614_clk;
  logic [0:0] f614_rst;
  logic [31:0] f614_rdata;
  sr_buffer_32_1 f614(.wen(f614_wen), .wdata(f614_wdata), .clk(f614_clk), .rst(f614_rst), .rdata(f614_rdata));
  assign f614_clk = clk;
  assign f614_rst = rst;
  // Bindings to f614

  // f616
  logic [0:0] f616_wen;
  logic [31:0] f616_wdata;
  logic [0:0] f616_clk;
  logic [0:0] f616_rst;
  logic [31:0] f616_rdata;
  sr_buffer_32_1 f616(.wen(f616_wen), .wdata(f616_wdata), .clk(f616_clk), .rst(f616_rst), .rdata(f616_rdata));
  assign f616_clk = clk;
  assign f616_rst = rst;
  // Bindings to f616

  // f618
  logic [0:0] f618_wen;
  logic [31:0] f618_wdata;
  logic [0:0] f618_clk;
  logic [0:0] f618_rst;
  logic [31:0] f618_rdata;
  sr_buffer_32_1 f618(.wen(f618_wen), .wdata(f618_wdata), .clk(f618_clk), .rst(f618_rst), .rdata(f618_rdata));
  assign f618_clk = clk;
  assign f618_rst = rst;
  // Bindings to f618

  // f620
  logic [0:0] f620_wen;
  logic [31:0] f620_wdata;
  logic [0:0] f620_clk;
  logic [0:0] f620_rst;
  logic [31:0] f620_rdata;
  sr_buffer_32_1 f620(.wen(f620_wen), .wdata(f620_wdata), .clk(f620_clk), .rst(f620_rst), .rdata(f620_rdata));
  assign f620_clk = clk;
  assign f620_rst = rst;
  // Bindings to f620

  // f622
  logic [0:0] f622_wen;
  logic [31:0] f622_wdata;
  logic [0:0] f622_clk;
  logic [0:0] f622_rst;
  logic [31:0] f622_rdata;
  sr_buffer_32_1 f622(.wen(f622_wen), .wdata(f622_wdata), .clk(f622_clk), .rst(f622_rst), .rdata(f622_rdata));
  assign f622_clk = clk;
  assign f622_rst = rst;
  // Bindings to f622

  // f624
  logic [0:0] f624_wen;
  logic [31:0] f624_wdata;
  logic [0:0] f624_clk;
  logic [0:0] f624_rst;
  logic [31:0] f624_rdata;
  sr_buffer_32_1 f624(.wen(f624_wen), .wdata(f624_wdata), .clk(f624_clk), .rst(f624_rst), .rdata(f624_rdata));
  assign f624_clk = clk;
  assign f624_rst = rst;
  // Bindings to f624

  // f626
  logic [0:0] f626_wen;
  logic [31:0] f626_wdata;
  logic [0:0] f626_clk;
  logic [0:0] f626_rst;
  logic [31:0] f626_rdata;
  sr_buffer_32_1 f626(.wen(f626_wen), .wdata(f626_wdata), .clk(f626_clk), .rst(f626_rst), .rdata(f626_rdata));
  assign f626_clk = clk;
  assign f626_rst = rst;
  // Bindings to f626

  // f628
  logic [0:0] f628_wen;
  logic [31:0] f628_wdata;
  logic [0:0] f628_clk;
  logic [0:0] f628_rst;
  logic [31:0] f628_rdata;
  sr_buffer_32_1 f628(.wen(f628_wen), .wdata(f628_wdata), .clk(f628_clk), .rst(f628_rst), .rdata(f628_rdata));
  assign f628_clk = clk;
  assign f628_rst = rst;
  // Bindings to f628

  // f630
  logic [0:0] f630_wen;
  logic [31:0] f630_wdata;
  logic [0:0] f630_clk;
  logic [0:0] f630_rst;
  logic [31:0] f630_rdata;
  sr_buffer_32_1 f630(.wen(f630_wen), .wdata(f630_wdata), .clk(f630_clk), .rst(f630_rst), .rdata(f630_rdata));
  assign f630_clk = clk;
  assign f630_rst = rst;
  // Bindings to f630

  // f632
  logic [0:0] f632_wen;
  logic [31:0] f632_wdata;
  logic [0:0] f632_clk;
  logic [0:0] f632_rst;
  logic [31:0] f632_rdata;
  sr_buffer_32_1 f632(.wen(f632_wen), .wdata(f632_wdata), .clk(f632_clk), .rst(f632_rst), .rdata(f632_rdata));
  assign f632_clk = clk;
  assign f632_rst = rst;
  // Bindings to f632

  // f634
  logic [0:0] f634_wen;
  logic [31:0] f634_wdata;
  logic [0:0] f634_clk;
  logic [0:0] f634_rst;
  logic [31:0] f634_rdata;
  sr_buffer_32_1 f634(.wen(f634_wen), .wdata(f634_wdata), .clk(f634_clk), .rst(f634_rst), .rdata(f634_rdata));
  assign f634_clk = clk;
  assign f634_rst = rst;
  // Bindings to f634

  // f636
  logic [0:0] f636_wen;
  logic [31:0] f636_wdata;
  logic [0:0] f636_clk;
  logic [0:0] f636_rst;
  logic [31:0] f636_rdata;
  sr_buffer_32_1 f636(.wen(f636_wen), .wdata(f636_wdata), .clk(f636_clk), .rst(f636_rst), .rdata(f636_rdata));
  assign f636_clk = clk;
  assign f636_rst = rst;
  // Bindings to f636

  // f638
  logic [0:0] f638_wen;
  logic [31:0] f638_wdata;
  logic [0:0] f638_clk;
  logic [0:0] f638_rst;
  logic [31:0] f638_rdata;
  sr_buffer_32_1 f638(.wen(f638_wen), .wdata(f638_wdata), .clk(f638_clk), .rst(f638_rst), .rdata(f638_rdata));
  assign f638_clk = clk;
  assign f638_rst = rst;
  // Bindings to f638

  // f640
  logic [0:0] f640_wen;
  logic [31:0] f640_wdata;
  logic [0:0] f640_clk;
  logic [0:0] f640_rst;
  logic [31:0] f640_rdata;
  sr_buffer_32_1 f640(.wen(f640_wen), .wdata(f640_wdata), .clk(f640_clk), .rst(f640_rst), .rdata(f640_rdata));
  assign f640_clk = clk;
  assign f640_rst = rst;
  // Bindings to f640

  // f642
  logic [0:0] f642_wen;
  logic [31:0] f642_wdata;
  logic [0:0] f642_clk;
  logic [0:0] f642_rst;
  logic [31:0] f642_rdata;
  sr_buffer_32_1 f642(.wen(f642_wen), .wdata(f642_wdata), .clk(f642_clk), .rst(f642_rst), .rdata(f642_rdata));
  assign f642_clk = clk;
  assign f642_rst = rst;
  // Bindings to f642

  // f644
  logic [0:0] f644_wen;
  logic [31:0] f644_wdata;
  logic [0:0] f644_clk;
  logic [0:0] f644_rst;
  logic [31:0] f644_rdata;
  sr_buffer_32_1 f644(.wen(f644_wen), .wdata(f644_wdata), .clk(f644_clk), .rst(f644_rst), .rdata(f644_rdata));
  assign f644_clk = clk;
  assign f644_rst = rst;
  // Bindings to f644

  // f646
  logic [0:0] f646_wen;
  logic [31:0] f646_wdata;
  logic [0:0] f646_clk;
  logic [0:0] f646_rst;
  logic [31:0] f646_rdata;
  sr_buffer_32_1 f646(.wen(f646_wen), .wdata(f646_wdata), .clk(f646_clk), .rst(f646_rst), .rdata(f646_rdata));
  assign f646_clk = clk;
  assign f646_rst = rst;
  // Bindings to f646

  // f648
  logic [0:0] f648_wen;
  logic [31:0] f648_wdata;
  logic [0:0] f648_clk;
  logic [0:0] f648_rst;
  logic [31:0] f648_rdata;
  sr_buffer_32_1 f648(.wen(f648_wen), .wdata(f648_wdata), .clk(f648_clk), .rst(f648_rst), .rdata(f648_rdata));
  assign f648_clk = clk;
  assign f648_rst = rst;
  // Bindings to f648

  // f650
  logic [0:0] f650_wen;
  logic [31:0] f650_wdata;
  logic [0:0] f650_clk;
  logic [0:0] f650_rst;
  logic [31:0] f650_rdata;
  sr_buffer_32_1 f650(.wen(f650_wen), .wdata(f650_wdata), .clk(f650_clk), .rst(f650_rst), .rdata(f650_rdata));
  assign f650_clk = clk;
  assign f650_rst = rst;
  // Bindings to f650

  // f652
  logic [0:0] f652_wen;
  logic [31:0] f652_wdata;
  logic [0:0] f652_clk;
  logic [0:0] f652_rst;
  logic [31:0] f652_rdata;
  sr_buffer_32_1 f652(.wen(f652_wen), .wdata(f652_wdata), .clk(f652_clk), .rst(f652_rst), .rdata(f652_rdata));
  assign f652_clk = clk;
  assign f652_rst = rst;
  // Bindings to f652

  // f654
  logic [0:0] f654_wen;
  logic [31:0] f654_wdata;
  logic [0:0] f654_clk;
  logic [0:0] f654_rst;
  logic [31:0] f654_rdata;
  sr_buffer_32_1 f654(.wen(f654_wen), .wdata(f654_wdata), .clk(f654_clk), .rst(f654_rst), .rdata(f654_rdata));
  assign f654_clk = clk;
  assign f654_rst = rst;
  // Bindings to f654

  // f656
  logic [0:0] f656_wen;
  logic [31:0] f656_wdata;
  logic [0:0] f656_clk;
  logic [0:0] f656_rst;
  logic [31:0] f656_rdata;
  sr_buffer_32_1 f656(.wen(f656_wen), .wdata(f656_wdata), .clk(f656_clk), .rst(f656_rst), .rdata(f656_rdata));
  assign f656_clk = clk;
  assign f656_rst = rst;
  // Bindings to f656

  // f658
  logic [0:0] f658_wen;
  logic [31:0] f658_wdata;
  logic [0:0] f658_clk;
  logic [0:0] f658_rst;
  logic [31:0] f658_rdata;
  sr_buffer_32_1 f658(.wen(f658_wen), .wdata(f658_wdata), .clk(f658_clk), .rst(f658_rst), .rdata(f658_rdata));
  assign f658_clk = clk;
  assign f658_rst = rst;
  // Bindings to f658

  // f660
  logic [0:0] f660_wen;
  logic [31:0] f660_wdata;
  logic [0:0] f660_clk;
  logic [0:0] f660_rst;
  logic [31:0] f660_rdata;
  sr_buffer_32_1 f660(.wen(f660_wen), .wdata(f660_wdata), .clk(f660_clk), .rst(f660_rst), .rdata(f660_rdata));
  assign f660_clk = clk;
  assign f660_rst = rst;
  // Bindings to f660

  // f662
  logic [0:0] f662_wen;
  logic [31:0] f662_wdata;
  logic [0:0] f662_clk;
  logic [0:0] f662_rst;
  logic [31:0] f662_rdata;
  sr_buffer_32_1 f662(.wen(f662_wen), .wdata(f662_wdata), .clk(f662_clk), .rst(f662_rst), .rdata(f662_rdata));
  assign f662_clk = clk;
  assign f662_rst = rst;
  // Bindings to f662

  // f664
  logic [0:0] f664_wen;
  logic [31:0] f664_wdata;
  logic [0:0] f664_clk;
  logic [0:0] f664_rst;
  logic [31:0] f664_rdata;
  sr_buffer_32_1 f664(.wen(f664_wen), .wdata(f664_wdata), .clk(f664_clk), .rst(f664_rst), .rdata(f664_rdata));
  assign f664_clk = clk;
  assign f664_rst = rst;
  // Bindings to f664

  // f666
  logic [0:0] f666_wen;
  logic [31:0] f666_wdata;
  logic [0:0] f666_clk;
  logic [0:0] f666_rst;
  logic [31:0] f666_rdata;
  sr_buffer_32_1 f666(.wen(f666_wen), .wdata(f666_wdata), .clk(f666_clk), .rst(f666_rst), .rdata(f666_rdata));
  assign f666_clk = clk;
  assign f666_rst = rst;
  // Bindings to f666

  // f668
  logic [0:0] f668_wen;
  logic [31:0] f668_wdata;
  logic [0:0] f668_clk;
  logic [0:0] f668_rst;
  logic [31:0] f668_rdata;
  sr_buffer_32_1 f668(.wen(f668_wen), .wdata(f668_wdata), .clk(f668_clk), .rst(f668_rst), .rdata(f668_rdata));
  assign f668_clk = clk;
  assign f668_rst = rst;
  // Bindings to f668

  // f670
  logic [0:0] f670_wen;
  logic [31:0] f670_wdata;
  logic [0:0] f670_clk;
  logic [0:0] f670_rst;
  logic [31:0] f670_rdata;
  sr_buffer_32_1 f670(.wen(f670_wen), .wdata(f670_wdata), .clk(f670_clk), .rst(f670_rst), .rdata(f670_rdata));
  assign f670_clk = clk;
  assign f670_rst = rst;
  // Bindings to f670

  // f672
  logic [0:0] f672_wen;
  logic [31:0] f672_wdata;
  logic [0:0] f672_clk;
  logic [0:0] f672_rst;
  logic [31:0] f672_rdata;
  sr_buffer_32_1 f672(.wen(f672_wen), .wdata(f672_wdata), .clk(f672_clk), .rst(f672_rst), .rdata(f672_rdata));
  assign f672_clk = clk;
  assign f672_rst = rst;
  // Bindings to f672

  // f674
  logic [0:0] f674_wen;
  logic [31:0] f674_wdata;
  logic [0:0] f674_clk;
  logic [0:0] f674_rst;
  logic [31:0] f674_rdata;
  sr_buffer_32_1 f674(.wen(f674_wen), .wdata(f674_wdata), .clk(f674_clk), .rst(f674_rst), .rdata(f674_rdata));
  assign f674_clk = clk;
  assign f674_rst = rst;
  // Bindings to f674

  // f676
  logic [0:0] f676_wen;
  logic [31:0] f676_wdata;
  logic [0:0] f676_clk;
  logic [0:0] f676_rst;
  logic [31:0] f676_rdata;
  sr_buffer_32_1 f676(.wen(f676_wen), .wdata(f676_wdata), .clk(f676_clk), .rst(f676_rst), .rdata(f676_rdata));
  assign f676_clk = clk;
  assign f676_rst = rst;
  // Bindings to f676

  // f678
  logic [0:0] f678_wen;
  logic [31:0] f678_wdata;
  logic [0:0] f678_clk;
  logic [0:0] f678_rst;
  logic [31:0] f678_rdata;
  sr_buffer_32_1 f678(.wen(f678_wen), .wdata(f678_wdata), .clk(f678_clk), .rst(f678_rst), .rdata(f678_rdata));
  assign f678_clk = clk;
  assign f678_rst = rst;
  // Bindings to f678

  // f680
  logic [0:0] f680_wen;
  logic [31:0] f680_wdata;
  logic [0:0] f680_clk;
  logic [0:0] f680_rst;
  logic [31:0] f680_rdata;
  sr_buffer_32_1 f680(.wen(f680_wen), .wdata(f680_wdata), .clk(f680_clk), .rst(f680_rst), .rdata(f680_rdata));
  assign f680_clk = clk;
  assign f680_rst = rst;
  // Bindings to f680

  // f682
  logic [0:0] f682_wen;
  logic [31:0] f682_wdata;
  logic [0:0] f682_clk;
  logic [0:0] f682_rst;
  logic [31:0] f682_rdata;
  sr_buffer_32_1 f682(.wen(f682_wen), .wdata(f682_wdata), .clk(f682_clk), .rst(f682_rst), .rdata(f682_rdata));
  assign f682_clk = clk;
  assign f682_rst = rst;
  // Bindings to f682

  // f684
  logic [0:0] f684_wen;
  logic [31:0] f684_wdata;
  logic [0:0] f684_clk;
  logic [0:0] f684_rst;
  logic [31:0] f684_rdata;
  sr_buffer_32_1 f684(.wen(f684_wen), .wdata(f684_wdata), .clk(f684_clk), .rst(f684_rst), .rdata(f684_rdata));
  assign f684_clk = clk;
  assign f684_rst = rst;
  // Bindings to f684

  // f686
  logic [0:0] f686_wen;
  logic [31:0] f686_wdata;
  logic [0:0] f686_clk;
  logic [0:0] f686_rst;
  logic [31:0] f686_rdata;
  sr_buffer_32_1 f686(.wen(f686_wen), .wdata(f686_wdata), .clk(f686_clk), .rst(f686_rst), .rdata(f686_rdata));
  assign f686_clk = clk;
  assign f686_rst = rst;
  // Bindings to f686

  // f688
  logic [0:0] f688_wen;
  logic [31:0] f688_wdata;
  logic [0:0] f688_clk;
  logic [0:0] f688_rst;
  logic [31:0] f688_rdata;
  sr_buffer_32_1 f688(.wen(f688_wen), .wdata(f688_wdata), .clk(f688_clk), .rst(f688_rst), .rdata(f688_rdata));
  assign f688_clk = clk;
  assign f688_rst = rst;
  // Bindings to f688

  // f690
  logic [0:0] f690_wen;
  logic [31:0] f690_wdata;
  logic [0:0] f690_clk;
  logic [0:0] f690_rst;
  logic [31:0] f690_rdata;
  sr_buffer_32_1 f690(.wen(f690_wen), .wdata(f690_wdata), .clk(f690_clk), .rst(f690_rst), .rdata(f690_rdata));
  assign f690_clk = clk;
  assign f690_rst = rst;
  // Bindings to f690

  // f692
  logic [0:0] f692_wen;
  logic [31:0] f692_wdata;
  logic [0:0] f692_clk;
  logic [0:0] f692_rst;
  logic [31:0] f692_rdata;
  sr_buffer_32_1 f692(.wen(f692_wen), .wdata(f692_wdata), .clk(f692_clk), .rst(f692_rst), .rdata(f692_rdata));
  assign f692_clk = clk;
  assign f692_rst = rst;
  // Bindings to f692

  // f694
  logic [0:0] f694_wen;
  logic [31:0] f694_wdata;
  logic [0:0] f694_clk;
  logic [0:0] f694_rst;
  logic [31:0] f694_rdata;
  sr_buffer_32_1 f694(.wen(f694_wen), .wdata(f694_wdata), .clk(f694_clk), .rst(f694_rst), .rdata(f694_rdata));
  assign f694_clk = clk;
  assign f694_rst = rst;
  // Bindings to f694

  // f696
  logic [0:0] f696_wen;
  logic [31:0] f696_wdata;
  logic [0:0] f696_clk;
  logic [0:0] f696_rst;
  logic [31:0] f696_rdata;
  sr_buffer_32_1 f696(.wen(f696_wen), .wdata(f696_wdata), .clk(f696_clk), .rst(f696_rst), .rdata(f696_rdata));
  assign f696_clk = clk;
  assign f696_rst = rst;
  // Bindings to f696

  // f698
  logic [0:0] f698_wen;
  logic [31:0] f698_wdata;
  logic [0:0] f698_clk;
  logic [0:0] f698_rst;
  logic [31:0] f698_rdata;
  sr_buffer_32_1 f698(.wen(f698_wen), .wdata(f698_wdata), .clk(f698_clk), .rst(f698_rst), .rdata(f698_rdata));
  assign f698_clk = clk;
  assign f698_rst = rst;
  // Bindings to f698

  // f700
  logic [0:0] f700_wen;
  logic [31:0] f700_wdata;
  logic [0:0] f700_clk;
  logic [0:0] f700_rst;
  logic [31:0] f700_rdata;
  sr_buffer_32_1 f700(.wen(f700_wen), .wdata(f700_wdata), .clk(f700_clk), .rst(f700_rst), .rdata(f700_rdata));
  assign f700_clk = clk;
  assign f700_rst = rst;
  // Bindings to f700

  // f702
  logic [0:0] f702_wen;
  logic [31:0] f702_wdata;
  logic [0:0] f702_clk;
  logic [0:0] f702_rst;
  logic [31:0] f702_rdata;
  sr_buffer_32_1 f702(.wen(f702_wen), .wdata(f702_wdata), .clk(f702_clk), .rst(f702_rst), .rdata(f702_rdata));
  assign f702_clk = clk;
  assign f702_rst = rst;
  // Bindings to f702

  // f704
  logic [0:0] f704_wen;
  logic [31:0] f704_wdata;
  logic [0:0] f704_clk;
  logic [0:0] f704_rst;
  logic [31:0] f704_rdata;
  sr_buffer_32_1 f704(.wen(f704_wen), .wdata(f704_wdata), .clk(f704_clk), .rst(f704_rst), .rdata(f704_rdata));
  assign f704_clk = clk;
  assign f704_rst = rst;
  // Bindings to f704

  // f706
  logic [0:0] f706_wen;
  logic [31:0] f706_wdata;
  logic [0:0] f706_clk;
  logic [0:0] f706_rst;
  logic [31:0] f706_rdata;
  sr_buffer_32_1 f706(.wen(f706_wen), .wdata(f706_wdata), .clk(f706_clk), .rst(f706_rst), .rdata(f706_rdata));
  assign f706_clk = clk;
  assign f706_rst = rst;
  // Bindings to f706

  // f708
  logic [0:0] f708_wen;
  logic [31:0] f708_wdata;
  logic [0:0] f708_clk;
  logic [0:0] f708_rst;
  logic [31:0] f708_rdata;
  sr_buffer_32_1 f708(.wen(f708_wen), .wdata(f708_wdata), .clk(f708_clk), .rst(f708_rst), .rdata(f708_rdata));
  assign f708_clk = clk;
  assign f708_rst = rst;
  // Bindings to f708

  // f710
  logic [0:0] f710_wen;
  logic [31:0] f710_wdata;
  logic [0:0] f710_clk;
  logic [0:0] f710_rst;
  logic [31:0] f710_rdata;
  sr_buffer_32_1 f710(.wen(f710_wen), .wdata(f710_wdata), .clk(f710_clk), .rst(f710_rst), .rdata(f710_rdata));
  assign f710_clk = clk;
  assign f710_rst = rst;
  // Bindings to f710

  // f712
  logic [0:0] f712_wen;
  logic [31:0] f712_wdata;
  logic [0:0] f712_clk;
  logic [0:0] f712_rst;
  logic [31:0] f712_rdata;
  sr_buffer_32_1 f712(.wen(f712_wen), .wdata(f712_wdata), .clk(f712_clk), .rst(f712_rst), .rdata(f712_rdata));
  assign f712_clk = clk;
  assign f712_rst = rst;
  // Bindings to f712

  // f714
  logic [0:0] f714_wen;
  logic [31:0] f714_wdata;
  logic [0:0] f714_clk;
  logic [0:0] f714_rst;
  logic [31:0] f714_rdata;
  sr_buffer_32_1 f714(.wen(f714_wen), .wdata(f714_wdata), .clk(f714_clk), .rst(f714_rst), .rdata(f714_rdata));
  assign f714_clk = clk;
  assign f714_rst = rst;
  // Bindings to f714

  // f716
  logic [0:0] f716_wen;
  logic [31:0] f716_wdata;
  logic [0:0] f716_clk;
  logic [0:0] f716_rst;
  logic [31:0] f716_rdata;
  sr_buffer_32_1 f716(.wen(f716_wen), .wdata(f716_wdata), .clk(f716_clk), .rst(f716_rst), .rdata(f716_rdata));
  assign f716_clk = clk;
  assign f716_rst = rst;
  // Bindings to f716

  // f718
  logic [0:0] f718_wen;
  logic [31:0] f718_wdata;
  logic [0:0] f718_clk;
  logic [0:0] f718_rst;
  logic [31:0] f718_rdata;
  sr_buffer_32_1 f718(.wen(f718_wen), .wdata(f718_wdata), .clk(f718_clk), .rst(f718_rst), .rdata(f718_rdata));
  assign f718_clk = clk;
  assign f718_rst = rst;
  // Bindings to f718

  // f720
  logic [0:0] f720_wen;
  logic [31:0] f720_wdata;
  logic [0:0] f720_clk;
  logic [0:0] f720_rst;
  logic [31:0] f720_rdata;
  sr_buffer_32_1 f720(.wen(f720_wen), .wdata(f720_wdata), .clk(f720_clk), .rst(f720_rst), .rdata(f720_rdata));
  assign f720_clk = clk;
  assign f720_rst = rst;
  // Bindings to f720

  // f722
  logic [0:0] f722_wen;
  logic [31:0] f722_wdata;
  logic [0:0] f722_clk;
  logic [0:0] f722_rst;
  logic [31:0] f722_rdata;
  sr_buffer_32_1 f722(.wen(f722_wen), .wdata(f722_wdata), .clk(f722_clk), .rst(f722_rst), .rdata(f722_rdata));
  assign f722_clk = clk;
  assign f722_rst = rst;
  // Bindings to f722

  // f724
  logic [0:0] f724_wen;
  logic [31:0] f724_wdata;
  logic [0:0] f724_clk;
  logic [0:0] f724_rst;
  logic [31:0] f724_rdata;
  sr_buffer_32_1 f724(.wen(f724_wen), .wdata(f724_wdata), .clk(f724_clk), .rst(f724_rst), .rdata(f724_rdata));
  assign f724_clk = clk;
  assign f724_rst = rst;
  // Bindings to f724

  // f726
  logic [0:0] f726_wen;
  logic [31:0] f726_wdata;
  logic [0:0] f726_clk;
  logic [0:0] f726_rst;
  logic [31:0] f726_rdata;
  sr_buffer_32_1 f726(.wen(f726_wen), .wdata(f726_wdata), .clk(f726_clk), .rst(f726_rst), .rdata(f726_rdata));
  assign f726_clk = clk;
  assign f726_rst = rst;
  // Bindings to f726

  // f728
  logic [0:0] f728_wen;
  logic [31:0] f728_wdata;
  logic [0:0] f728_clk;
  logic [0:0] f728_rst;
  logic [31:0] f728_rdata;
  sr_buffer_32_1 f728(.wen(f728_wen), .wdata(f728_wdata), .clk(f728_clk), .rst(f728_rst), .rdata(f728_rdata));
  assign f728_clk = clk;
  assign f728_rst = rst;
  // Bindings to f728

  // f730
  logic [0:0] f730_wen;
  logic [31:0] f730_wdata;
  logic [0:0] f730_clk;
  logic [0:0] f730_rst;
  logic [31:0] f730_rdata;
  sr_buffer_32_1 f730(.wen(f730_wen), .wdata(f730_wdata), .clk(f730_clk), .rst(f730_rst), .rdata(f730_rdata));
  assign f730_clk = clk;
  assign f730_rst = rst;
  // Bindings to f730

  // f732
  logic [0:0] f732_wen;
  logic [31:0] f732_wdata;
  logic [0:0] f732_clk;
  logic [0:0] f732_rst;
  logic [31:0] f732_rdata;
  sr_buffer_32_1 f732(.wen(f732_wen), .wdata(f732_wdata), .clk(f732_clk), .rst(f732_rst), .rdata(f732_rdata));
  assign f732_clk = clk;
  assign f732_rst = rst;
  // Bindings to f732

  // f734
  logic [0:0] f734_wen;
  logic [31:0] f734_wdata;
  logic [0:0] f734_clk;
  logic [0:0] f734_rst;
  logic [31:0] f734_rdata;
  sr_buffer_32_1 f734(.wen(f734_wen), .wdata(f734_wdata), .clk(f734_clk), .rst(f734_rst), .rdata(f734_rdata));
  assign f734_clk = clk;
  assign f734_rst = rst;
  // Bindings to f734

  // f736
  logic [0:0] f736_wen;
  logic [31:0] f736_wdata;
  logic [0:0] f736_clk;
  logic [0:0] f736_rst;
  logic [31:0] f736_rdata;
  sr_buffer_32_1 f736(.wen(f736_wen), .wdata(f736_wdata), .clk(f736_clk), .rst(f736_rst), .rdata(f736_rdata));
  assign f736_clk = clk;
  assign f736_rst = rst;
  // Bindings to f736

  // f738
  logic [0:0] f738_wen;
  logic [31:0] f738_wdata;
  logic [0:0] f738_clk;
  logic [0:0] f738_rst;
  logic [31:0] f738_rdata;
  sr_buffer_32_1 f738(.wen(f738_wen), .wdata(f738_wdata), .clk(f738_clk), .rst(f738_rst), .rdata(f738_rdata));
  assign f738_clk = clk;
  assign f738_rst = rst;
  // Bindings to f738

  // f740
  logic [0:0] f740_wen;
  logic [31:0] f740_wdata;
  logic [0:0] f740_clk;
  logic [0:0] f740_rst;
  logic [31:0] f740_rdata;
  sr_buffer_32_1 f740(.wen(f740_wen), .wdata(f740_wdata), .clk(f740_clk), .rst(f740_rst), .rdata(f740_rdata));
  assign f740_clk = clk;
  assign f740_rst = rst;
  // Bindings to f740

  // f742
  logic [0:0] f742_wen;
  logic [31:0] f742_wdata;
  logic [0:0] f742_clk;
  logic [0:0] f742_rst;
  logic [31:0] f742_rdata;
  sr_buffer_32_1 f742(.wen(f742_wen), .wdata(f742_wdata), .clk(f742_clk), .rst(f742_rst), .rdata(f742_rdata));
  assign f742_clk = clk;
  assign f742_rst = rst;
  // Bindings to f742

  // f744
  logic [0:0] f744_wen;
  logic [31:0] f744_wdata;
  logic [0:0] f744_clk;
  logic [0:0] f744_rst;
  logic [31:0] f744_rdata;
  sr_buffer_32_1 f744(.wen(f744_wen), .wdata(f744_wdata), .clk(f744_clk), .rst(f744_rst), .rdata(f744_rdata));
  assign f744_clk = clk;
  assign f744_rst = rst;
  // Bindings to f744

  // f746
  logic [0:0] f746_wen;
  logic [31:0] f746_wdata;
  logic [0:0] f746_clk;
  logic [0:0] f746_rst;
  logic [31:0] f746_rdata;
  sr_buffer_32_1 f746(.wen(f746_wen), .wdata(f746_wdata), .clk(f746_clk), .rst(f746_rst), .rdata(f746_rdata));
  assign f746_clk = clk;
  assign f746_rst = rst;
  // Bindings to f746

  // f748
  logic [0:0] f748_wen;
  logic [31:0] f748_wdata;
  logic [0:0] f748_clk;
  logic [0:0] f748_rst;
  logic [31:0] f748_rdata;
  sr_buffer_32_1 f748(.wen(f748_wen), .wdata(f748_wdata), .clk(f748_clk), .rst(f748_rst), .rdata(f748_rdata));
  assign f748_clk = clk;
  assign f748_rst = rst;
  // Bindings to f748

  // f750
  logic [0:0] f750_wen;
  logic [31:0] f750_wdata;
  logic [0:0] f750_clk;
  logic [0:0] f750_rst;
  logic [31:0] f750_rdata;
  sr_buffer_32_1 f750(.wen(f750_wen), .wdata(f750_wdata), .clk(f750_clk), .rst(f750_rst), .rdata(f750_rdata));
  assign f750_clk = clk;
  assign f750_rst = rst;
  // Bindings to f750

  // f752
  logic [0:0] f752_wen;
  logic [31:0] f752_wdata;
  logic [0:0] f752_clk;
  logic [0:0] f752_rst;
  logic [31:0] f752_rdata;
  sr_buffer_32_1 f752(.wen(f752_wen), .wdata(f752_wdata), .clk(f752_clk), .rst(f752_rst), .rdata(f752_rdata));
  assign f752_clk = clk;
  assign f752_rst = rst;
  // Bindings to f752

  // f754
  logic [0:0] f754_wen;
  logic [31:0] f754_wdata;
  logic [0:0] f754_clk;
  logic [0:0] f754_rst;
  logic [31:0] f754_rdata;
  sr_buffer_32_1 f754(.wen(f754_wen), .wdata(f754_wdata), .clk(f754_clk), .rst(f754_rst), .rdata(f754_rdata));
  assign f754_clk = clk;
  assign f754_rst = rst;
  // Bindings to f754

  // f756
  logic [0:0] f756_wen;
  logic [31:0] f756_wdata;
  logic [0:0] f756_clk;
  logic [0:0] f756_rst;
  logic [31:0] f756_rdata;
  sr_buffer_32_1 f756(.wen(f756_wen), .wdata(f756_wdata), .clk(f756_clk), .rst(f756_rst), .rdata(f756_rdata));
  assign f756_clk = clk;
  assign f756_rst = rst;
  // Bindings to f756

  // f758
  logic [0:0] f758_wen;
  logic [31:0] f758_wdata;
  logic [0:0] f758_clk;
  logic [0:0] f758_rst;
  logic [31:0] f758_rdata;
  sr_buffer_32_1 f758(.wen(f758_wen), .wdata(f758_wdata), .clk(f758_clk), .rst(f758_rst), .rdata(f758_rdata));
  assign f758_clk = clk;
  assign f758_rst = rst;
  // Bindings to f758

  // f760
  logic [0:0] f760_wen;
  logic [31:0] f760_wdata;
  logic [0:0] f760_clk;
  logic [0:0] f760_rst;
  logic [31:0] f760_rdata;
  sr_buffer_32_1 f760(.wen(f760_wen), .wdata(f760_wdata), .clk(f760_clk), .rst(f760_rst), .rdata(f760_rdata));
  assign f760_clk = clk;
  assign f760_rst = rst;
  // Bindings to f760

  // f762
  logic [0:0] f762_wen;
  logic [31:0] f762_wdata;
  logic [0:0] f762_clk;
  logic [0:0] f762_rst;
  logic [31:0] f762_rdata;
  sr_buffer_32_1 f762(.wen(f762_wen), .wdata(f762_wdata), .clk(f762_clk), .rst(f762_rst), .rdata(f762_rdata));
  assign f762_clk = clk;
  assign f762_rst = rst;
  // Bindings to f762

  // f764
  logic [0:0] f764_wen;
  logic [31:0] f764_wdata;
  logic [0:0] f764_clk;
  logic [0:0] f764_rst;
  logic [31:0] f764_rdata;
  sr_buffer_32_1 f764(.wen(f764_wen), .wdata(f764_wdata), .clk(f764_clk), .rst(f764_rst), .rdata(f764_rdata));
  assign f764_clk = clk;
  assign f764_rst = rst;
  // Bindings to f764

  // f766
  logic [0:0] f766_wen;
  logic [31:0] f766_wdata;
  logic [0:0] f766_clk;
  logic [0:0] f766_rst;
  logic [31:0] f766_rdata;
  sr_buffer_32_1 f766(.wen(f766_wen), .wdata(f766_wdata), .clk(f766_clk), .rst(f766_rst), .rdata(f766_rdata));
  assign f766_clk = clk;
  assign f766_rst = rst;
  // Bindings to f766

  // f768
  logic [0:0] f768_wen;
  logic [31:0] f768_wdata;
  logic [0:0] f768_clk;
  logic [0:0] f768_rst;
  logic [31:0] f768_rdata;
  sr_buffer_32_1 f768(.wen(f768_wen), .wdata(f768_wdata), .clk(f768_clk), .rst(f768_rst), .rdata(f768_rdata));
  assign f768_clk = clk;
  assign f768_rst = rst;
  // Bindings to f768

  // f770
  logic [0:0] f770_wen;
  logic [31:0] f770_wdata;
  logic [0:0] f770_clk;
  logic [0:0] f770_rst;
  logic [31:0] f770_rdata;
  sr_buffer_32_1 f770(.wen(f770_wen), .wdata(f770_wdata), .clk(f770_clk), .rst(f770_rst), .rdata(f770_rdata));
  assign f770_clk = clk;
  assign f770_rst = rst;
  // Bindings to f770

  // f772
  logic [0:0] f772_wen;
  logic [31:0] f772_wdata;
  logic [0:0] f772_clk;
  logic [0:0] f772_rst;
  logic [31:0] f772_rdata;
  sr_buffer_32_1 f772(.wen(f772_wen), .wdata(f772_wdata), .clk(f772_clk), .rst(f772_rst), .rdata(f772_rdata));
  assign f772_clk = clk;
  assign f772_rst = rst;
  // Bindings to f772

  // f774
  logic [0:0] f774_wen;
  logic [31:0] f774_wdata;
  logic [0:0] f774_clk;
  logic [0:0] f774_rst;
  logic [31:0] f774_rdata;
  sr_buffer_32_1 f774(.wen(f774_wen), .wdata(f774_wdata), .clk(f774_clk), .rst(f774_rst), .rdata(f774_rdata));
  assign f774_clk = clk;
  assign f774_rst = rst;
  // Bindings to f774

  // f776
  logic [0:0] f776_wen;
  logic [31:0] f776_wdata;
  logic [0:0] f776_clk;
  logic [0:0] f776_rst;
  logic [31:0] f776_rdata;
  sr_buffer_32_1 f776(.wen(f776_wen), .wdata(f776_wdata), .clk(f776_clk), .rst(f776_rst), .rdata(f776_rdata));
  assign f776_clk = clk;
  assign f776_rst = rst;
  // Bindings to f776

  // f778
  logic [0:0] f778_wen;
  logic [31:0] f778_wdata;
  logic [0:0] f778_clk;
  logic [0:0] f778_rst;
  logic [31:0] f778_rdata;
  sr_buffer_32_1 f778(.wen(f778_wen), .wdata(f778_wdata), .clk(f778_clk), .rst(f778_rst), .rdata(f778_rdata));
  assign f778_clk = clk;
  assign f778_rst = rst;
  // Bindings to f778

  // f780
  logic [0:0] f780_wen;
  logic [31:0] f780_wdata;
  logic [0:0] f780_clk;
  logic [0:0] f780_rst;
  logic [31:0] f780_rdata;
  sr_buffer_32_1 f780(.wen(f780_wen), .wdata(f780_wdata), .clk(f780_clk), .rst(f780_rst), .rdata(f780_rdata));
  assign f780_clk = clk;
  assign f780_rst = rst;
  // Bindings to f780

  // f782
  logic [0:0] f782_wen;
  logic [31:0] f782_wdata;
  logic [0:0] f782_clk;
  logic [0:0] f782_rst;
  logic [31:0] f782_rdata;
  sr_buffer_32_1 f782(.wen(f782_wen), .wdata(f782_wdata), .clk(f782_clk), .rst(f782_rst), .rdata(f782_rdata));
  assign f782_clk = clk;
  assign f782_rst = rst;
  // Bindings to f782

  // f784
  logic [0:0] f784_wen;
  logic [31:0] f784_wdata;
  logic [0:0] f784_clk;
  logic [0:0] f784_rst;
  logic [31:0] f784_rdata;
  sr_buffer_32_1 f784(.wen(f784_wen), .wdata(f784_wdata), .clk(f784_clk), .rst(f784_rst), .rdata(f784_rdata));
  assign f784_clk = clk;
  assign f784_rst = rst;
  // Bindings to f784

  // f786
  logic [0:0] f786_wen;
  logic [31:0] f786_wdata;
  logic [0:0] f786_clk;
  logic [0:0] f786_rst;
  logic [31:0] f786_rdata;
  sr_buffer_32_1 f786(.wen(f786_wen), .wdata(f786_wdata), .clk(f786_clk), .rst(f786_rst), .rdata(f786_rdata));
  assign f786_clk = clk;
  assign f786_rst = rst;
  // Bindings to f786

  // f788
  logic [0:0] f788_wen;
  logic [31:0] f788_wdata;
  logic [0:0] f788_clk;
  logic [0:0] f788_rst;
  logic [31:0] f788_rdata;
  sr_buffer_32_1 f788(.wen(f788_wen), .wdata(f788_wdata), .clk(f788_clk), .rst(f788_rst), .rdata(f788_rdata));
  assign f788_clk = clk;
  assign f788_rst = rst;
  // Bindings to f788

  // f790
  logic [0:0] f790_wen;
  logic [31:0] f790_wdata;
  logic [0:0] f790_clk;
  logic [0:0] f790_rst;
  logic [31:0] f790_rdata;
  sr_buffer_32_1 f790(.wen(f790_wen), .wdata(f790_wdata), .clk(f790_clk), .rst(f790_rst), .rdata(f790_rdata));
  assign f790_clk = clk;
  assign f790_rst = rst;
  // Bindings to f790

  // f792
  logic [0:0] f792_wen;
  logic [31:0] f792_wdata;
  logic [0:0] f792_clk;
  logic [0:0] f792_rst;
  logic [31:0] f792_rdata;
  sr_buffer_32_1 f792(.wen(f792_wen), .wdata(f792_wdata), .clk(f792_clk), .rst(f792_rst), .rdata(f792_rdata));
  assign f792_clk = clk;
  assign f792_rst = rst;
  // Bindings to f792

  // f794
  logic [0:0] f794_wen;
  logic [31:0] f794_wdata;
  logic [0:0] f794_clk;
  logic [0:0] f794_rst;
  logic [31:0] f794_rdata;
  sr_buffer_32_1 f794(.wen(f794_wen), .wdata(f794_wdata), .clk(f794_clk), .rst(f794_rst), .rdata(f794_rdata));
  assign f794_clk = clk;
  assign f794_rst = rst;
  // Bindings to f794

  // f796
  logic [0:0] f796_wen;
  logic [31:0] f796_wdata;
  logic [0:0] f796_clk;
  logic [0:0] f796_rst;
  logic [31:0] f796_rdata;
  sr_buffer_32_1 f796(.wen(f796_wen), .wdata(f796_wdata), .clk(f796_clk), .rst(f796_rst), .rdata(f796_rdata));
  assign f796_clk = clk;
  assign f796_rst = rst;
  // Bindings to f796

  // f798
  logic [0:0] f798_wen;
  logic [31:0] f798_wdata;
  logic [0:0] f798_clk;
  logic [0:0] f798_rst;
  logic [31:0] f798_rdata;
  sr_buffer_32_1 f798(.wen(f798_wen), .wdata(f798_wdata), .clk(f798_clk), .rst(f798_rst), .rdata(f798_rdata));
  assign f798_clk = clk;
  assign f798_rst = rst;
  // Bindings to f798

  // f800
  logic [0:0] f800_wen;
  logic [31:0] f800_wdata;
  logic [0:0] f800_clk;
  logic [0:0] f800_rst;
  logic [31:0] f800_rdata;
  sr_buffer_32_1 f800(.wen(f800_wen), .wdata(f800_wdata), .clk(f800_clk), .rst(f800_rst), .rdata(f800_rdata));
  assign f800_clk = clk;
  assign f800_rst = rst;
  // Bindings to f800

  // f802
  logic [0:0] f802_wen;
  logic [31:0] f802_wdata;
  logic [0:0] f802_clk;
  logic [0:0] f802_rst;
  logic [31:0] f802_rdata;
  sr_buffer_32_1 f802(.wen(f802_wen), .wdata(f802_wdata), .clk(f802_clk), .rst(f802_rst), .rdata(f802_rdata));
  assign f802_clk = clk;
  assign f802_rst = rst;
  // Bindings to f802

  // f804
  logic [0:0] f804_wen;
  logic [31:0] f804_wdata;
  logic [0:0] f804_clk;
  logic [0:0] f804_rst;
  logic [31:0] f804_rdata;
  sr_buffer_32_1 f804(.wen(f804_wen), .wdata(f804_wdata), .clk(f804_clk), .rst(f804_rst), .rdata(f804_rdata));
  assign f804_clk = clk;
  assign f804_rst = rst;
  // Bindings to f804

  // f806
  logic [0:0] f806_wen;
  logic [31:0] f806_wdata;
  logic [0:0] f806_clk;
  logic [0:0] f806_rst;
  logic [31:0] f806_rdata;
  sr_buffer_32_1 f806(.wen(f806_wen), .wdata(f806_wdata), .clk(f806_clk), .rst(f806_rst), .rdata(f806_rdata));
  assign f806_clk = clk;
  assign f806_rst = rst;
  // Bindings to f806

  // f808
  logic [0:0] f808_wen;
  logic [31:0] f808_wdata;
  logic [0:0] f808_clk;
  logic [0:0] f808_rst;
  logic [31:0] f808_rdata;
  sr_buffer_32_1 f808(.wen(f808_wen), .wdata(f808_wdata), .clk(f808_clk), .rst(f808_rst), .rdata(f808_rdata));
  assign f808_clk = clk;
  assign f808_rst = rst;
  // Bindings to f808

  // f810
  logic [0:0] f810_wen;
  logic [31:0] f810_wdata;
  logic [0:0] f810_clk;
  logic [0:0] f810_rst;
  logic [31:0] f810_rdata;
  sr_buffer_32_1 f810(.wen(f810_wen), .wdata(f810_wdata), .clk(f810_clk), .rst(f810_rst), .rdata(f810_rdata));
  assign f810_clk = clk;
  assign f810_rst = rst;
  // Bindings to f810

  // f812
  logic [0:0] f812_wen;
  logic [31:0] f812_wdata;
  logic [0:0] f812_clk;
  logic [0:0] f812_rst;
  logic [31:0] f812_rdata;
  sr_buffer_32_1 f812(.wen(f812_wen), .wdata(f812_wdata), .clk(f812_clk), .rst(f812_rst), .rdata(f812_rdata));
  assign f812_clk = clk;
  assign f812_rst = rst;
  // Bindings to f812

  // f814
  logic [0:0] f814_wen;
  logic [31:0] f814_wdata;
  logic [0:0] f814_clk;
  logic [0:0] f814_rst;
  logic [31:0] f814_rdata;
  sr_buffer_32_1 f814(.wen(f814_wen), .wdata(f814_wdata), .clk(f814_clk), .rst(f814_rst), .rdata(f814_rdata));
  assign f814_clk = clk;
  assign f814_rst = rst;
  // Bindings to f814

  // f816
  logic [0:0] f816_wen;
  logic [31:0] f816_wdata;
  logic [0:0] f816_clk;
  logic [0:0] f816_rst;
  logic [31:0] f816_rdata;
  sr_buffer_32_1 f816(.wen(f816_wen), .wdata(f816_wdata), .clk(f816_clk), .rst(f816_rst), .rdata(f816_rdata));
  assign f816_clk = clk;
  assign f816_rst = rst;
  // Bindings to f816

  // f818
  logic [0:0] f818_wen;
  logic [31:0] f818_wdata;
  logic [0:0] f818_clk;
  logic [0:0] f818_rst;
  logic [31:0] f818_rdata;
  sr_buffer_32_1 f818(.wen(f818_wen), .wdata(f818_wdata), .clk(f818_clk), .rst(f818_rst), .rdata(f818_rdata));
  assign f818_clk = clk;
  assign f818_rst = rst;
  // Bindings to f818

  // f820
  logic [0:0] f820_wen;
  logic [31:0] f820_wdata;
  logic [0:0] f820_clk;
  logic [0:0] f820_rst;
  logic [31:0] f820_rdata;
  sr_buffer_32_1 f820(.wen(f820_wen), .wdata(f820_wdata), .clk(f820_clk), .rst(f820_rst), .rdata(f820_rdata));
  assign f820_clk = clk;
  assign f820_rst = rst;
  // Bindings to f820

  // f822
  logic [0:0] f822_wen;
  logic [31:0] f822_wdata;
  logic [0:0] f822_clk;
  logic [0:0] f822_rst;
  logic [31:0] f822_rdata;
  sr_buffer_32_1 f822(.wen(f822_wen), .wdata(f822_wdata), .clk(f822_clk), .rst(f822_rst), .rdata(f822_rdata));
  assign f822_clk = clk;
  assign f822_rst = rst;
  // Bindings to f822

  // f824
  logic [0:0] f824_wen;
  logic [31:0] f824_wdata;
  logic [0:0] f824_clk;
  logic [0:0] f824_rst;
  logic [31:0] f824_rdata;
  sr_buffer_32_1 f824(.wen(f824_wen), .wdata(f824_wdata), .clk(f824_clk), .rst(f824_rst), .rdata(f824_rdata));
  assign f824_clk = clk;
  assign f824_rst = rst;
  // Bindings to f824

  // f826
  logic [0:0] f826_wen;
  logic [31:0] f826_wdata;
  logic [0:0] f826_clk;
  logic [0:0] f826_rst;
  logic [31:0] f826_rdata;
  sr_buffer_32_1 f826(.wen(f826_wen), .wdata(f826_wdata), .clk(f826_clk), .rst(f826_rst), .rdata(f826_rdata));
  assign f826_clk = clk;
  assign f826_rst = rst;
  // Bindings to f826

  // f828
  logic [0:0] f828_wen;
  logic [31:0] f828_wdata;
  logic [0:0] f828_clk;
  logic [0:0] f828_rst;
  logic [31:0] f828_rdata;
  sr_buffer_32_1 f828(.wen(f828_wen), .wdata(f828_wdata), .clk(f828_clk), .rst(f828_rst), .rdata(f828_rdata));
  assign f828_clk = clk;
  assign f828_rst = rst;
  // Bindings to f828

  // f830
  logic [0:0] f830_wen;
  logic [31:0] f830_wdata;
  logic [0:0] f830_clk;
  logic [0:0] f830_rst;
  logic [31:0] f830_rdata;
  sr_buffer_32_1 f830(.wen(f830_wen), .wdata(f830_wdata), .clk(f830_clk), .rst(f830_rst), .rdata(f830_rdata));
  assign f830_clk = clk;
  assign f830_rst = rst;
  // Bindings to f830

  // f832
  logic [0:0] f832_wen;
  logic [31:0] f832_wdata;
  logic [0:0] f832_clk;
  logic [0:0] f832_rst;
  logic [31:0] f832_rdata;
  sr_buffer_32_1 f832(.wen(f832_wen), .wdata(f832_wdata), .clk(f832_clk), .rst(f832_rst), .rdata(f832_rdata));
  assign f832_clk = clk;
  assign f832_rst = rst;
  // Bindings to f832

  // f834
  logic [0:0] f834_wen;
  logic [31:0] f834_wdata;
  logic [0:0] f834_clk;
  logic [0:0] f834_rst;
  logic [31:0] f834_rdata;
  sr_buffer_32_1 f834(.wen(f834_wen), .wdata(f834_wdata), .clk(f834_clk), .rst(f834_rst), .rdata(f834_rdata));
  assign f834_clk = clk;
  assign f834_rst = rst;
  // Bindings to f834

  // f836
  logic [0:0] f836_wen;
  logic [31:0] f836_wdata;
  logic [0:0] f836_clk;
  logic [0:0] f836_rst;
  logic [31:0] f836_rdata;
  sr_buffer_32_1 f836(.wen(f836_wen), .wdata(f836_wdata), .clk(f836_clk), .rst(f836_rst), .rdata(f836_rdata));
  assign f836_clk = clk;
  assign f836_rst = rst;
  // Bindings to f836

  // f838
  logic [0:0] f838_wen;
  logic [31:0] f838_wdata;
  logic [0:0] f838_clk;
  logic [0:0] f838_rst;
  logic [31:0] f838_rdata;
  sr_buffer_32_1 f838(.wen(f838_wen), .wdata(f838_wdata), .clk(f838_clk), .rst(f838_rst), .rdata(f838_rdata));
  assign f838_clk = clk;
  assign f838_rst = rst;
  // Bindings to f838

  // f840
  logic [0:0] f840_wen;
  logic [31:0] f840_wdata;
  logic [0:0] f840_clk;
  logic [0:0] f840_rst;
  logic [31:0] f840_rdata;
  sr_buffer_32_1 f840(.wen(f840_wen), .wdata(f840_wdata), .clk(f840_clk), .rst(f840_rst), .rdata(f840_rdata));
  assign f840_clk = clk;
  assign f840_rst = rst;
  // Bindings to f840

  // f842
  logic [0:0] f842_wen;
  logic [31:0] f842_wdata;
  logic [0:0] f842_clk;
  logic [0:0] f842_rst;
  logic [31:0] f842_rdata;
  sr_buffer_32_1 f842(.wen(f842_wen), .wdata(f842_wdata), .clk(f842_clk), .rst(f842_rst), .rdata(f842_rdata));
  assign f842_clk = clk;
  assign f842_rst = rst;
  // Bindings to f842

  // f844
  logic [0:0] f844_wen;
  logic [31:0] f844_wdata;
  logic [0:0] f844_clk;
  logic [0:0] f844_rst;
  logic [31:0] f844_rdata;
  sr_buffer_32_1 f844(.wen(f844_wen), .wdata(f844_wdata), .clk(f844_clk), .rst(f844_rst), .rdata(f844_rdata));
  assign f844_clk = clk;
  assign f844_rst = rst;
  // Bindings to f844

  // f846
  logic [0:0] f846_wen;
  logic [31:0] f846_wdata;
  logic [0:0] f846_clk;
  logic [0:0] f846_rst;
  logic [31:0] f846_rdata;
  sr_buffer_32_1 f846(.wen(f846_wen), .wdata(f846_wdata), .clk(f846_clk), .rst(f846_rst), .rdata(f846_rdata));
  assign f846_clk = clk;
  assign f846_rst = rst;
  // Bindings to f846

  // f848
  logic [0:0] f848_wen;
  logic [31:0] f848_wdata;
  logic [0:0] f848_clk;
  logic [0:0] f848_rst;
  logic [31:0] f848_rdata;
  sr_buffer_32_1 f848(.wen(f848_wen), .wdata(f848_wdata), .clk(f848_clk), .rst(f848_rst), .rdata(f848_rdata));
  assign f848_clk = clk;
  assign f848_rst = rst;
  // Bindings to f848

  // f850
  logic [0:0] f850_wen;
  logic [31:0] f850_wdata;
  logic [0:0] f850_clk;
  logic [0:0] f850_rst;
  logic [31:0] f850_rdata;
  sr_buffer_32_1 f850(.wen(f850_wen), .wdata(f850_wdata), .clk(f850_clk), .rst(f850_rst), .rdata(f850_rdata));
  assign f850_clk = clk;
  assign f850_rst = rst;
  // Bindings to f850

  // f852
  logic [0:0] f852_wen;
  logic [31:0] f852_wdata;
  logic [0:0] f852_clk;
  logic [0:0] f852_rst;
  logic [31:0] f852_rdata;
  sr_buffer_32_1 f852(.wen(f852_wen), .wdata(f852_wdata), .clk(f852_clk), .rst(f852_rst), .rdata(f852_rdata));
  assign f852_clk = clk;
  assign f852_rst = rst;
  // Bindings to f852

  // f854
  logic [0:0] f854_wen;
  logic [31:0] f854_wdata;
  logic [0:0] f854_clk;
  logic [0:0] f854_rst;
  logic [31:0] f854_rdata;
  sr_buffer_32_1 f854(.wen(f854_wen), .wdata(f854_wdata), .clk(f854_clk), .rst(f854_rst), .rdata(f854_rdata));
  assign f854_clk = clk;
  assign f854_rst = rst;
  // Bindings to f854

  // f856
  logic [0:0] f856_wen;
  logic [31:0] f856_wdata;
  logic [0:0] f856_clk;
  logic [0:0] f856_rst;
  logic [31:0] f856_rdata;
  sr_buffer_32_1 f856(.wen(f856_wen), .wdata(f856_wdata), .clk(f856_clk), .rst(f856_rst), .rdata(f856_rdata));
  assign f856_clk = clk;
  assign f856_rst = rst;
  // Bindings to f856

  // f858
  logic [0:0] f858_wen;
  logic [31:0] f858_wdata;
  logic [0:0] f858_clk;
  logic [0:0] f858_rst;
  logic [31:0] f858_rdata;
  sr_buffer_32_1 f858(.wen(f858_wen), .wdata(f858_wdata), .clk(f858_clk), .rst(f858_rst), .rdata(f858_rdata));
  assign f858_clk = clk;
  assign f858_rst = rst;
  // Bindings to f858

  // f860
  logic [0:0] f860_wen;
  logic [31:0] f860_wdata;
  logic [0:0] f860_clk;
  logic [0:0] f860_rst;
  logic [31:0] f860_rdata;
  sr_buffer_32_1 f860(.wen(f860_wen), .wdata(f860_wdata), .clk(f860_clk), .rst(f860_rst), .rdata(f860_rdata));
  assign f860_clk = clk;
  assign f860_rst = rst;
  // Bindings to f860

  // f862
  logic [0:0] f862_wen;
  logic [31:0] f862_wdata;
  logic [0:0] f862_clk;
  logic [0:0] f862_rst;
  logic [31:0] f862_rdata;
  sr_buffer_32_1 f862(.wen(f862_wen), .wdata(f862_wdata), .clk(f862_clk), .rst(f862_rst), .rdata(f862_rdata));
  assign f862_clk = clk;
  assign f862_rst = rst;
  // Bindings to f862

  // f864
  logic [0:0] f864_wen;
  logic [31:0] f864_wdata;
  logic [0:0] f864_clk;
  logic [0:0] f864_rst;
  logic [31:0] f864_rdata;
  sr_buffer_32_1 f864(.wen(f864_wen), .wdata(f864_wdata), .clk(f864_clk), .rst(f864_rst), .rdata(f864_rdata));
  assign f864_clk = clk;
  assign f864_rst = rst;
  // Bindings to f864

  // f866
  logic [0:0] f866_wen;
  logic [31:0] f866_wdata;
  logic [0:0] f866_clk;
  logic [0:0] f866_rst;
  logic [31:0] f866_rdata;
  sr_buffer_32_1 f866(.wen(f866_wen), .wdata(f866_wdata), .clk(f866_clk), .rst(f866_rst), .rdata(f866_rdata));
  assign f866_clk = clk;
  assign f866_rst = rst;
  // Bindings to f866

  // f868
  logic [0:0] f868_wen;
  logic [31:0] f868_wdata;
  logic [0:0] f868_clk;
  logic [0:0] f868_rst;
  logic [31:0] f868_rdata;
  sr_buffer_32_1 f868(.wen(f868_wen), .wdata(f868_wdata), .clk(f868_clk), .rst(f868_rst), .rdata(f868_rdata));
  assign f868_clk = clk;
  assign f868_rst = rst;
  // Bindings to f868

  // f870
  logic [0:0] f870_wen;
  logic [31:0] f870_wdata;
  logic [0:0] f870_clk;
  logic [0:0] f870_rst;
  logic [31:0] f870_rdata;
  sr_buffer_32_1 f870(.wen(f870_wen), .wdata(f870_wdata), .clk(f870_clk), .rst(f870_rst), .rdata(f870_rdata));
  assign f870_clk = clk;
  assign f870_rst = rst;
  // Bindings to f870

  // f872
  logic [0:0] f872_wen;
  logic [31:0] f872_wdata;
  logic [0:0] f872_clk;
  logic [0:0] f872_rst;
  logic [31:0] f872_rdata;
  sr_buffer_32_1 f872(.wen(f872_wen), .wdata(f872_wdata), .clk(f872_clk), .rst(f872_rst), .rdata(f872_rdata));
  assign f872_clk = clk;
  assign f872_rst = rst;
  // Bindings to f872

  // f874
  logic [0:0] f874_wen;
  logic [31:0] f874_wdata;
  logic [0:0] f874_clk;
  logic [0:0] f874_rst;
  logic [31:0] f874_rdata;
  sr_buffer_32_1 f874(.wen(f874_wen), .wdata(f874_wdata), .clk(f874_clk), .rst(f874_rst), .rdata(f874_rdata));
  assign f874_clk = clk;
  assign f874_rst = rst;
  // Bindings to f874

  // f876
  logic [0:0] f876_wen;
  logic [31:0] f876_wdata;
  logic [0:0] f876_clk;
  logic [0:0] f876_rst;
  logic [31:0] f876_rdata;
  sr_buffer_32_1 f876(.wen(f876_wen), .wdata(f876_wdata), .clk(f876_clk), .rst(f876_rst), .rdata(f876_rdata));
  assign f876_clk = clk;
  assign f876_rst = rst;
  // Bindings to f876

  // f878
  logic [0:0] f878_wen;
  logic [31:0] f878_wdata;
  logic [0:0] f878_clk;
  logic [0:0] f878_rst;
  logic [31:0] f878_rdata;
  sr_buffer_32_1 f878(.wen(f878_wen), .wdata(f878_wdata), .clk(f878_clk), .rst(f878_rst), .rdata(f878_rdata));
  assign f878_clk = clk;
  assign f878_rst = rst;
  // Bindings to f878

  // f880
  logic [0:0] f880_wen;
  logic [31:0] f880_wdata;
  logic [0:0] f880_clk;
  logic [0:0] f880_rst;
  logic [31:0] f880_rdata;
  sr_buffer_32_1 f880(.wen(f880_wen), .wdata(f880_wdata), .clk(f880_clk), .rst(f880_rst), .rdata(f880_rdata));
  assign f880_clk = clk;
  assign f880_rst = rst;
  // Bindings to f880

  // f882
  logic [0:0] f882_wen;
  logic [31:0] f882_wdata;
  logic [0:0] f882_clk;
  logic [0:0] f882_rst;
  logic [31:0] f882_rdata;
  sr_buffer_32_1 f882(.wen(f882_wen), .wdata(f882_wdata), .clk(f882_clk), .rst(f882_rst), .rdata(f882_rdata));
  assign f882_clk = clk;
  assign f882_rst = rst;
  // Bindings to f882

  // f884
  logic [0:0] f884_wen;
  logic [31:0] f884_wdata;
  logic [0:0] f884_clk;
  logic [0:0] f884_rst;
  logic [31:0] f884_rdata;
  sr_buffer_32_1 f884(.wen(f884_wen), .wdata(f884_wdata), .clk(f884_clk), .rst(f884_rst), .rdata(f884_rdata));
  assign f884_clk = clk;
  assign f884_rst = rst;
  // Bindings to f884

  // f886
  logic [0:0] f886_wen;
  logic [31:0] f886_wdata;
  logic [0:0] f886_clk;
  logic [0:0] f886_rst;
  logic [31:0] f886_rdata;
  sr_buffer_32_1 f886(.wen(f886_wen), .wdata(f886_wdata), .clk(f886_clk), .rst(f886_rst), .rdata(f886_rdata));
  assign f886_clk = clk;
  assign f886_rst = rst;
  // Bindings to f886

  // f888
  logic [0:0] f888_wen;
  logic [31:0] f888_wdata;
  logic [0:0] f888_clk;
  logic [0:0] f888_rst;
  logic [31:0] f888_rdata;
  sr_buffer_32_1 f888(.wen(f888_wen), .wdata(f888_wdata), .clk(f888_clk), .rst(f888_rst), .rdata(f888_rdata));
  assign f888_clk = clk;
  assign f888_rst = rst;
  // Bindings to f888

  // f890
  logic [0:0] f890_wen;
  logic [31:0] f890_wdata;
  logic [0:0] f890_clk;
  logic [0:0] f890_rst;
  logic [31:0] f890_rdata;
  sr_buffer_32_1 f890(.wen(f890_wen), .wdata(f890_wdata), .clk(f890_clk), .rst(f890_rst), .rdata(f890_rdata));
  assign f890_clk = clk;
  assign f890_rst = rst;
  // Bindings to f890

  // f892
  logic [0:0] f892_wen;
  logic [31:0] f892_wdata;
  logic [0:0] f892_clk;
  logic [0:0] f892_rst;
  logic [31:0] f892_rdata;
  sr_buffer_32_1 f892(.wen(f892_wen), .wdata(f892_wdata), .clk(f892_clk), .rst(f892_rst), .rdata(f892_rdata));
  assign f892_clk = clk;
  assign f892_rst = rst;
  // Bindings to f892

  // f894
  logic [0:0] f894_wen;
  logic [31:0] f894_wdata;
  logic [0:0] f894_clk;
  logic [0:0] f894_rst;
  logic [31:0] f894_rdata;
  sr_buffer_32_1 f894(.wen(f894_wen), .wdata(f894_wdata), .clk(f894_clk), .rst(f894_rst), .rdata(f894_rdata));
  assign f894_clk = clk;
  assign f894_rst = rst;
  // Bindings to f894

  // f896
  logic [0:0] f896_wen;
  logic [31:0] f896_wdata;
  logic [0:0] f896_clk;
  logic [0:0] f896_rst;
  logic [31:0] f896_rdata;
  sr_buffer_32_1 f896(.wen(f896_wen), .wdata(f896_wdata), .clk(f896_clk), .rst(f896_rst), .rdata(f896_rdata));
  assign f896_clk = clk;
  assign f896_rst = rst;
  // Bindings to f896

  // f898
  logic [0:0] f898_wen;
  logic [31:0] f898_wdata;
  logic [0:0] f898_clk;
  logic [0:0] f898_rst;
  logic [31:0] f898_rdata;
  sr_buffer_32_1 f898(.wen(f898_wen), .wdata(f898_wdata), .clk(f898_clk), .rst(f898_rst), .rdata(f898_rdata));
  assign f898_clk = clk;
  assign f898_rst = rst;
  // Bindings to f898

  // f900
  logic [0:0] f900_wen;
  logic [31:0] f900_wdata;
  logic [0:0] f900_clk;
  logic [0:0] f900_rst;
  logic [31:0] f900_rdata;
  sr_buffer_32_1 f900(.wen(f900_wen), .wdata(f900_wdata), .clk(f900_clk), .rst(f900_rst), .rdata(f900_rdata));
  assign f900_clk = clk;
  assign f900_rst = rst;
  // Bindings to f900

  // f902
  logic [0:0] f902_wen;
  logic [31:0] f902_wdata;
  logic [0:0] f902_clk;
  logic [0:0] f902_rst;
  logic [31:0] f902_rdata;
  sr_buffer_32_1 f902(.wen(f902_wen), .wdata(f902_wdata), .clk(f902_clk), .rst(f902_rst), .rdata(f902_rdata));
  assign f902_clk = clk;
  assign f902_rst = rst;
  // Bindings to f902

  // f904
  logic [0:0] f904_wen;
  logic [31:0] f904_wdata;
  logic [0:0] f904_clk;
  logic [0:0] f904_rst;
  logic [31:0] f904_rdata;
  sr_buffer_32_1 f904(.wen(f904_wen), .wdata(f904_wdata), .clk(f904_clk), .rst(f904_rst), .rdata(f904_rdata));
  assign f904_clk = clk;
  assign f904_rst = rst;
  // Bindings to f904

  // f906
  logic [0:0] f906_wen;
  logic [31:0] f906_wdata;
  logic [0:0] f906_clk;
  logic [0:0] f906_rst;
  logic [31:0] f906_rdata;
  sr_buffer_32_1 f906(.wen(f906_wen), .wdata(f906_wdata), .clk(f906_clk), .rst(f906_rst), .rdata(f906_rdata));
  assign f906_clk = clk;
  assign f906_rst = rst;
  // Bindings to f906

  // f908
  logic [0:0] f908_wen;
  logic [31:0] f908_wdata;
  logic [0:0] f908_clk;
  logic [0:0] f908_rst;
  logic [31:0] f908_rdata;
  sr_buffer_32_1 f908(.wen(f908_wen), .wdata(f908_wdata), .clk(f908_clk), .rst(f908_rst), .rdata(f908_rdata));
  assign f908_clk = clk;
  assign f908_rst = rst;
  // Bindings to f908

  // f910
  logic [0:0] f910_wen;
  logic [31:0] f910_wdata;
  logic [0:0] f910_clk;
  logic [0:0] f910_rst;
  logic [31:0] f910_rdata;
  sr_buffer_32_1 f910(.wen(f910_wen), .wdata(f910_wdata), .clk(f910_clk), .rst(f910_rst), .rdata(f910_rdata));
  assign f910_clk = clk;
  assign f910_rst = rst;
  // Bindings to f910

  // f912
  logic [0:0] f912_wen;
  logic [31:0] f912_wdata;
  logic [0:0] f912_clk;
  logic [0:0] f912_rst;
  logic [31:0] f912_rdata;
  sr_buffer_32_1 f912(.wen(f912_wen), .wdata(f912_wdata), .clk(f912_clk), .rst(f912_rst), .rdata(f912_rdata));
  assign f912_clk = clk;
  assign f912_rst = rst;
  // Bindings to f912

  // f914
  logic [0:0] f914_wen;
  logic [31:0] f914_wdata;
  logic [0:0] f914_clk;
  logic [0:0] f914_rst;
  logic [31:0] f914_rdata;
  sr_buffer_32_1 f914(.wen(f914_wen), .wdata(f914_wdata), .clk(f914_clk), .rst(f914_rst), .rdata(f914_rdata));
  assign f914_clk = clk;
  assign f914_rst = rst;
  // Bindings to f914

  // f916
  logic [0:0] f916_wen;
  logic [31:0] f916_wdata;
  logic [0:0] f916_clk;
  logic [0:0] f916_rst;
  logic [31:0] f916_rdata;
  sr_buffer_32_1 f916(.wen(f916_wen), .wdata(f916_wdata), .clk(f916_clk), .rst(f916_rst), .rdata(f916_rdata));
  assign f916_clk = clk;
  assign f916_rst = rst;
  // Bindings to f916

  // f918
  logic [0:0] f918_wen;
  logic [31:0] f918_wdata;
  logic [0:0] f918_clk;
  logic [0:0] f918_rst;
  logic [31:0] f918_rdata;
  sr_buffer_32_1 f918(.wen(f918_wen), .wdata(f918_wdata), .clk(f918_clk), .rst(f918_rst), .rdata(f918_rdata));
  assign f918_clk = clk;
  assign f918_rst = rst;
  // Bindings to f918

  // f920
  logic [0:0] f920_wen;
  logic [31:0] f920_wdata;
  logic [0:0] f920_clk;
  logic [0:0] f920_rst;
  logic [31:0] f920_rdata;
  sr_buffer_32_1 f920(.wen(f920_wen), .wdata(f920_wdata), .clk(f920_clk), .rst(f920_rst), .rdata(f920_rdata));
  assign f920_clk = clk;
  assign f920_rst = rst;
  // Bindings to f920

  // f922
  logic [0:0] f922_wen;
  logic [31:0] f922_wdata;
  logic [0:0] f922_clk;
  logic [0:0] f922_rst;
  logic [31:0] f922_rdata;
  sr_buffer_32_1 f922(.wen(f922_wen), .wdata(f922_wdata), .clk(f922_clk), .rst(f922_rst), .rdata(f922_rdata));
  assign f922_clk = clk;
  assign f922_rst = rst;
  // Bindings to f922

  // f924
  logic [0:0] f924_wen;
  logic [31:0] f924_wdata;
  logic [0:0] f924_clk;
  logic [0:0] f924_rst;
  logic [31:0] f924_rdata;
  sr_buffer_32_1 f924(.wen(f924_wen), .wdata(f924_wdata), .clk(f924_clk), .rst(f924_rst), .rdata(f924_rdata));
  assign f924_clk = clk;
  assign f924_rst = rst;
  // Bindings to f924

  // f926
  logic [0:0] f926_wen;
  logic [31:0] f926_wdata;
  logic [0:0] f926_clk;
  logic [0:0] f926_rst;
  logic [31:0] f926_rdata;
  sr_buffer_32_1 f926(.wen(f926_wen), .wdata(f926_wdata), .clk(f926_clk), .rst(f926_rst), .rdata(f926_rdata));
  assign f926_clk = clk;
  assign f926_rst = rst;
  // Bindings to f926

  // f928
  logic [0:0] f928_wen;
  logic [31:0] f928_wdata;
  logic [0:0] f928_clk;
  logic [0:0] f928_rst;
  logic [31:0] f928_rdata;
  sr_buffer_32_1 f928(.wen(f928_wen), .wdata(f928_wdata), .clk(f928_clk), .rst(f928_rst), .rdata(f928_rdata));
  assign f928_clk = clk;
  assign f928_rst = rst;
  // Bindings to f928

  // f930
  logic [0:0] f930_wen;
  logic [31:0] f930_wdata;
  logic [0:0] f930_clk;
  logic [0:0] f930_rst;
  logic [31:0] f930_rdata;
  sr_buffer_32_1 f930(.wen(f930_wen), .wdata(f930_wdata), .clk(f930_clk), .rst(f930_rst), .rdata(f930_rdata));
  assign f930_clk = clk;
  assign f930_rst = rst;
  // Bindings to f930

  // f932
  logic [0:0] f932_wen;
  logic [31:0] f932_wdata;
  logic [0:0] f932_clk;
  logic [0:0] f932_rst;
  logic [31:0] f932_rdata;
  sr_buffer_32_1 f932(.wen(f932_wen), .wdata(f932_wdata), .clk(f932_clk), .rst(f932_rst), .rdata(f932_rdata));
  assign f932_clk = clk;
  assign f932_rst = rst;
  // Bindings to f932

  // f934
  logic [0:0] f934_wen;
  logic [31:0] f934_wdata;
  logic [0:0] f934_clk;
  logic [0:0] f934_rst;
  logic [31:0] f934_rdata;
  sr_buffer_32_1 f934(.wen(f934_wen), .wdata(f934_wdata), .clk(f934_clk), .rst(f934_rst), .rdata(f934_rdata));
  assign f934_clk = clk;
  assign f934_rst = rst;
  // Bindings to f934

  // f936
  logic [0:0] f936_wen;
  logic [31:0] f936_wdata;
  logic [0:0] f936_clk;
  logic [0:0] f936_rst;
  logic [31:0] f936_rdata;
  sr_buffer_32_1 f936(.wen(f936_wen), .wdata(f936_wdata), .clk(f936_clk), .rst(f936_rst), .rdata(f936_rdata));
  assign f936_clk = clk;
  assign f936_rst = rst;
  // Bindings to f936

  // f938
  logic [0:0] f938_wen;
  logic [31:0] f938_wdata;
  logic [0:0] f938_clk;
  logic [0:0] f938_rst;
  logic [31:0] f938_rdata;
  sr_buffer_32_1 f938(.wen(f938_wen), .wdata(f938_wdata), .clk(f938_clk), .rst(f938_rst), .rdata(f938_rdata));
  assign f938_clk = clk;
  assign f938_rst = rst;
  // Bindings to f938

  // f940
  logic [0:0] f940_wen;
  logic [31:0] f940_wdata;
  logic [0:0] f940_clk;
  logic [0:0] f940_rst;
  logic [31:0] f940_rdata;
  sr_buffer_32_1 f940(.wen(f940_wen), .wdata(f940_wdata), .clk(f940_clk), .rst(f940_rst), .rdata(f940_rdata));
  assign f940_clk = clk;
  assign f940_rst = rst;
  // Bindings to f940

  // f942
  logic [0:0] f942_wen;
  logic [31:0] f942_wdata;
  logic [0:0] f942_clk;
  logic [0:0] f942_rst;
  logic [31:0] f942_rdata;
  sr_buffer_32_1 f942(.wen(f942_wen), .wdata(f942_wdata), .clk(f942_clk), .rst(f942_rst), .rdata(f942_rdata));
  assign f942_clk = clk;
  assign f942_rst = rst;
  // Bindings to f942

  // f944
  logic [0:0] f944_wen;
  logic [31:0] f944_wdata;
  logic [0:0] f944_clk;
  logic [0:0] f944_rst;
  logic [31:0] f944_rdata;
  sr_buffer_32_1 f944(.wen(f944_wen), .wdata(f944_wdata), .clk(f944_clk), .rst(f944_rst), .rdata(f944_rdata));
  assign f944_clk = clk;
  assign f944_rst = rst;
  // Bindings to f944

  // f946
  logic [0:0] f946_wen;
  logic [31:0] f946_wdata;
  logic [0:0] f946_clk;
  logic [0:0] f946_rst;
  logic [31:0] f946_rdata;
  sr_buffer_32_1 f946(.wen(f946_wen), .wdata(f946_wdata), .clk(f946_clk), .rst(f946_rst), .rdata(f946_rdata));
  assign f946_clk = clk;
  assign f946_rst = rst;
  // Bindings to f946

  // f948
  logic [0:0] f948_wen;
  logic [31:0] f948_wdata;
  logic [0:0] f948_clk;
  logic [0:0] f948_rst;
  logic [31:0] f948_rdata;
  sr_buffer_32_1 f948(.wen(f948_wen), .wdata(f948_wdata), .clk(f948_clk), .rst(f948_rst), .rdata(f948_rdata));
  assign f948_clk = clk;
  assign f948_rst = rst;
  // Bindings to f948

  // f950
  logic [0:0] f950_wen;
  logic [31:0] f950_wdata;
  logic [0:0] f950_clk;
  logic [0:0] f950_rst;
  logic [31:0] f950_rdata;
  sr_buffer_32_1 f950(.wen(f950_wen), .wdata(f950_wdata), .clk(f950_clk), .rst(f950_rst), .rdata(f950_rdata));
  assign f950_clk = clk;
  assign f950_rst = rst;
  // Bindings to f950

  // f952
  logic [0:0] f952_wen;
  logic [31:0] f952_wdata;
  logic [0:0] f952_clk;
  logic [0:0] f952_rst;
  logic [31:0] f952_rdata;
  sr_buffer_32_1 f952(.wen(f952_wen), .wdata(f952_wdata), .clk(f952_clk), .rst(f952_rst), .rdata(f952_rdata));
  assign f952_clk = clk;
  assign f952_rst = rst;
  // Bindings to f952

  // f954
  logic [0:0] f954_wen;
  logic [31:0] f954_wdata;
  logic [0:0] f954_clk;
  logic [0:0] f954_rst;
  logic [31:0] f954_rdata;
  sr_buffer_32_1 f954(.wen(f954_wen), .wdata(f954_wdata), .clk(f954_clk), .rst(f954_rst), .rdata(f954_rdata));
  assign f954_clk = clk;
  assign f954_rst = rst;
  // Bindings to f954

  // f956
  logic [0:0] f956_wen;
  logic [31:0] f956_wdata;
  logic [0:0] f956_clk;
  logic [0:0] f956_rst;
  logic [31:0] f956_rdata;
  sr_buffer_32_1 f956(.wen(f956_wen), .wdata(f956_wdata), .clk(f956_clk), .rst(f956_rst), .rdata(f956_rdata));
  assign f956_clk = clk;
  assign f956_rst = rst;
  // Bindings to f956

  // f958
  logic [0:0] f958_wen;
  logic [31:0] f958_wdata;
  logic [0:0] f958_clk;
  logic [0:0] f958_rst;
  logic [31:0] f958_rdata;
  sr_buffer_32_1 f958(.wen(f958_wen), .wdata(f958_wdata), .clk(f958_clk), .rst(f958_rst), .rdata(f958_rdata));
  assign f958_clk = clk;
  assign f958_rst = rst;
  // Bindings to f958

  // f960
  logic [0:0] f960_wen;
  logic [31:0] f960_wdata;
  logic [0:0] f960_clk;
  logic [0:0] f960_rst;
  logic [31:0] f960_rdata;
  sr_buffer_32_1 f960(.wen(f960_wen), .wdata(f960_wdata), .clk(f960_clk), .rst(f960_rst), .rdata(f960_rdata));
  assign f960_clk = clk;
  assign f960_rst = rst;
  // Bindings to f960

  // f962
  logic [0:0] f962_wen;
  logic [31:0] f962_wdata;
  logic [0:0] f962_clk;
  logic [0:0] f962_rst;
  logic [31:0] f962_rdata;
  sr_buffer_32_1 f962(.wen(f962_wen), .wdata(f962_wdata), .clk(f962_clk), .rst(f962_rst), .rdata(f962_rdata));
  assign f962_clk = clk;
  assign f962_rst = rst;
  // Bindings to f962

  // f964
  logic [0:0] f964_wen;
  logic [31:0] f964_wdata;
  logic [0:0] f964_clk;
  logic [0:0] f964_rst;
  logic [31:0] f964_rdata;
  sr_buffer_32_1 f964(.wen(f964_wen), .wdata(f964_wdata), .clk(f964_clk), .rst(f964_rst), .rdata(f964_rdata));
  assign f964_clk = clk;
  assign f964_rst = rst;
  // Bindings to f964

  // f966
  logic [0:0] f966_wen;
  logic [31:0] f966_wdata;
  logic [0:0] f966_clk;
  logic [0:0] f966_rst;
  logic [31:0] f966_rdata;
  sr_buffer_32_1 f966(.wen(f966_wen), .wdata(f966_wdata), .clk(f966_clk), .rst(f966_rst), .rdata(f966_rdata));
  assign f966_clk = clk;
  assign f966_rst = rst;
  // Bindings to f966

  // f968
  logic [0:0] f968_wen;
  logic [31:0] f968_wdata;
  logic [0:0] f968_clk;
  logic [0:0] f968_rst;
  logic [31:0] f968_rdata;
  sr_buffer_32_1 f968(.wen(f968_wen), .wdata(f968_wdata), .clk(f968_clk), .rst(f968_rst), .rdata(f968_rdata));
  assign f968_clk = clk;
  assign f968_rst = rst;
  // Bindings to f968

  // f970
  logic [0:0] f970_wen;
  logic [31:0] f970_wdata;
  logic [0:0] f970_clk;
  logic [0:0] f970_rst;
  logic [31:0] f970_rdata;
  sr_buffer_32_1 f970(.wen(f970_wen), .wdata(f970_wdata), .clk(f970_clk), .rst(f970_rst), .rdata(f970_rdata));
  assign f970_clk = clk;
  assign f970_rst = rst;
  // Bindings to f970

  // f972
  logic [0:0] f972_wen;
  logic [31:0] f972_wdata;
  logic [0:0] f972_clk;
  logic [0:0] f972_rst;
  logic [31:0] f972_rdata;
  sr_buffer_32_1 f972(.wen(f972_wen), .wdata(f972_wdata), .clk(f972_clk), .rst(f972_rst), .rdata(f972_rdata));
  assign f972_clk = clk;
  assign f972_rst = rst;
  // Bindings to f972

  // f974
  logic [0:0] f974_wen;
  logic [31:0] f974_wdata;
  logic [0:0] f974_clk;
  logic [0:0] f974_rst;
  logic [31:0] f974_rdata;
  sr_buffer_32_1 f974(.wen(f974_wen), .wdata(f974_wdata), .clk(f974_clk), .rst(f974_rst), .rdata(f974_rdata));
  assign f974_clk = clk;
  assign f974_rst = rst;
  // Bindings to f974

  // f976
  logic [0:0] f976_wen;
  logic [31:0] f976_wdata;
  logic [0:0] f976_clk;
  logic [0:0] f976_rst;
  logic [31:0] f976_rdata;
  sr_buffer_32_1 f976(.wen(f976_wen), .wdata(f976_wdata), .clk(f976_clk), .rst(f976_rst), .rdata(f976_rdata));
  assign f976_clk = clk;
  assign f976_rst = rst;
  // Bindings to f976

  // f978
  logic [0:0] f978_wen;
  logic [31:0] f978_wdata;
  logic [0:0] f978_clk;
  logic [0:0] f978_rst;
  logic [31:0] f978_rdata;
  sr_buffer_32_1 f978(.wen(f978_wen), .wdata(f978_wdata), .clk(f978_clk), .rst(f978_rst), .rdata(f978_rdata));
  assign f978_clk = clk;
  assign f978_rst = rst;
  // Bindings to f978

  // f980
  logic [0:0] f980_wen;
  logic [31:0] f980_wdata;
  logic [0:0] f980_clk;
  logic [0:0] f980_rst;
  logic [31:0] f980_rdata;
  sr_buffer_32_1 f980(.wen(f980_wen), .wdata(f980_wdata), .clk(f980_clk), .rst(f980_rst), .rdata(f980_rdata));
  assign f980_clk = clk;
  assign f980_rst = rst;
  // Bindings to f980

  // f982
  logic [0:0] f982_wen;
  logic [31:0] f982_wdata;
  logic [0:0] f982_clk;
  logic [0:0] f982_rst;
  logic [31:0] f982_rdata;
  sr_buffer_32_1 f982(.wen(f982_wen), .wdata(f982_wdata), .clk(f982_clk), .rst(f982_rst), .rdata(f982_rdata));
  assign f982_clk = clk;
  assign f982_rst = rst;
  // Bindings to f982

  // f984
  logic [0:0] f984_wen;
  logic [31:0] f984_wdata;
  logic [0:0] f984_clk;
  logic [0:0] f984_rst;
  logic [31:0] f984_rdata;
  sr_buffer_32_1 f984(.wen(f984_wen), .wdata(f984_wdata), .clk(f984_clk), .rst(f984_rst), .rdata(f984_rdata));
  assign f984_clk = clk;
  assign f984_rst = rst;
  // Bindings to f984

  // f986
  logic [0:0] f986_wen;
  logic [31:0] f986_wdata;
  logic [0:0] f986_clk;
  logic [0:0] f986_rst;
  logic [31:0] f986_rdata;
  sr_buffer_32_1 f986(.wen(f986_wen), .wdata(f986_wdata), .clk(f986_clk), .rst(f986_rst), .rdata(f986_rdata));
  assign f986_clk = clk;
  assign f986_rst = rst;
  // Bindings to f986

  // f988
  logic [0:0] f988_wen;
  logic [31:0] f988_wdata;
  logic [0:0] f988_clk;
  logic [0:0] f988_rst;
  logic [31:0] f988_rdata;
  sr_buffer_32_1 f988(.wen(f988_wen), .wdata(f988_wdata), .clk(f988_clk), .rst(f988_rst), .rdata(f988_rdata));
  assign f988_clk = clk;
  assign f988_rst = rst;
  // Bindings to f988

  // f990
  logic [0:0] f990_wen;
  logic [31:0] f990_wdata;
  logic [0:0] f990_clk;
  logic [0:0] f990_rst;
  logic [31:0] f990_rdata;
  sr_buffer_32_1 f990(.wen(f990_wen), .wdata(f990_wdata), .clk(f990_clk), .rst(f990_rst), .rdata(f990_rdata));
  assign f990_clk = clk;
  assign f990_rst = rst;
  // Bindings to f990

  // f992
  logic [0:0] f992_wen;
  logic [31:0] f992_wdata;
  logic [0:0] f992_clk;
  logic [0:0] f992_rst;
  logic [31:0] f992_rdata;
  sr_buffer_32_1 f992(.wen(f992_wen), .wdata(f992_wdata), .clk(f992_clk), .rst(f992_rst), .rdata(f992_rdata));
  assign f992_clk = clk;
  assign f992_rst = rst;
  // Bindings to f992

  // f994
  logic [0:0] f994_wen;
  logic [31:0] f994_wdata;
  logic [0:0] f994_clk;
  logic [0:0] f994_rst;
  logic [31:0] f994_rdata;
  sr_buffer_32_1 f994(.wen(f994_wen), .wdata(f994_wdata), .clk(f994_clk), .rst(f994_rst), .rdata(f994_rdata));
  assign f994_clk = clk;
  assign f994_rst = rst;
  // Bindings to f994

  // f996
  logic [0:0] f996_wen;
  logic [31:0] f996_wdata;
  logic [0:0] f996_clk;
  logic [0:0] f996_rst;
  logic [31:0] f996_rdata;
  sr_buffer_32_1 f996(.wen(f996_wen), .wdata(f996_wdata), .clk(f996_clk), .rst(f996_rst), .rdata(f996_rdata));
  assign f996_clk = clk;
  assign f996_rst = rst;
  // Bindings to f996

  // f998
  logic [0:0] f998_wen;
  logic [31:0] f998_wdata;
  logic [0:0] f998_clk;
  logic [0:0] f998_rst;
  logic [31:0] f998_rdata;
  sr_buffer_32_1 f998(.wen(f998_wen), .wdata(f998_wdata), .clk(f998_clk), .rst(f998_rst), .rdata(f998_rdata));
  assign f998_clk = clk;
  assign f998_rst = rst;
  // Bindings to f998

  // f1000
  logic [0:0] f1000_wen;
  logic [31:0] f1000_wdata;
  logic [0:0] f1000_clk;
  logic [0:0] f1000_rst;
  logic [31:0] f1000_rdata;
  sr_buffer_32_1 f1000(.wen(f1000_wen), .wdata(f1000_wdata), .clk(f1000_clk), .rst(f1000_rst), .rdata(f1000_rdata));
  assign f1000_clk = clk;
  assign f1000_rst = rst;
  // Bindings to f1000

  // f1002
  logic [0:0] f1002_wen;
  logic [31:0] f1002_wdata;
  logic [0:0] f1002_clk;
  logic [0:0] f1002_rst;
  logic [31:0] f1002_rdata;
  sr_buffer_32_1 f1002(.wen(f1002_wen), .wdata(f1002_wdata), .clk(f1002_clk), .rst(f1002_rst), .rdata(f1002_rdata));
  assign f1002_clk = clk;
  assign f1002_rst = rst;
  // Bindings to f1002

  // f1004
  logic [0:0] f1004_wen;
  logic [31:0] f1004_wdata;
  logic [0:0] f1004_clk;
  logic [0:0] f1004_rst;
  logic [31:0] f1004_rdata;
  sr_buffer_32_1 f1004(.wen(f1004_wen), .wdata(f1004_wdata), .clk(f1004_clk), .rst(f1004_rst), .rdata(f1004_rdata));
  assign f1004_clk = clk;
  assign f1004_rst = rst;
  // Bindings to f1004

  // f1006
  logic [0:0] f1006_wen;
  logic [31:0] f1006_wdata;
  logic [0:0] f1006_clk;
  logic [0:0] f1006_rst;
  logic [31:0] f1006_rdata;
  sr_buffer_32_1 f1006(.wen(f1006_wen), .wdata(f1006_wdata), .clk(f1006_clk), .rst(f1006_rst), .rdata(f1006_rdata));
  assign f1006_clk = clk;
  assign f1006_rst = rst;
  // Bindings to f1006

  // f1008
  logic [0:0] f1008_wen;
  logic [31:0] f1008_wdata;
  logic [0:0] f1008_clk;
  logic [0:0] f1008_rst;
  logic [31:0] f1008_rdata;
  sr_buffer_32_1 f1008(.wen(f1008_wen), .wdata(f1008_wdata), .clk(f1008_clk), .rst(f1008_rst), .rdata(f1008_rdata));
  assign f1008_clk = clk;
  assign f1008_rst = rst;
  // Bindings to f1008

  // f1010
  logic [0:0] f1010_wen;
  logic [31:0] f1010_wdata;
  logic [0:0] f1010_clk;
  logic [0:0] f1010_rst;
  logic [31:0] f1010_rdata;
  sr_buffer_32_1 f1010(.wen(f1010_wen), .wdata(f1010_wdata), .clk(f1010_clk), .rst(f1010_rst), .rdata(f1010_rdata));
  assign f1010_clk = clk;
  assign f1010_rst = rst;
  // Bindings to f1010

  // f1012
  logic [0:0] f1012_wen;
  logic [31:0] f1012_wdata;
  logic [0:0] f1012_clk;
  logic [0:0] f1012_rst;
  logic [31:0] f1012_rdata;
  sr_buffer_32_1 f1012(.wen(f1012_wen), .wdata(f1012_wdata), .clk(f1012_clk), .rst(f1012_rst), .rdata(f1012_rdata));
  assign f1012_clk = clk;
  assign f1012_rst = rst;
  // Bindings to f1012

  // f1014
  logic [0:0] f1014_wen;
  logic [31:0] f1014_wdata;
  logic [0:0] f1014_clk;
  logic [0:0] f1014_rst;
  logic [31:0] f1014_rdata;
  sr_buffer_32_1 f1014(.wen(f1014_wen), .wdata(f1014_wdata), .clk(f1014_clk), .rst(f1014_rst), .rdata(f1014_rdata));
  assign f1014_clk = clk;
  assign f1014_rst = rst;
  // Bindings to f1014

  // f1016
  logic [0:0] f1016_wen;
  logic [31:0] f1016_wdata;
  logic [0:0] f1016_clk;
  logic [0:0] f1016_rst;
  logic [31:0] f1016_rdata;
  sr_buffer_32_1 f1016(.wen(f1016_wen), .wdata(f1016_wdata), .clk(f1016_clk), .rst(f1016_rst), .rdata(f1016_rdata));
  assign f1016_clk = clk;
  assign f1016_rst = rst;
  // Bindings to f1016

  // f1018
  logic [0:0] f1018_wen;
  logic [31:0] f1018_wdata;
  logic [0:0] f1018_clk;
  logic [0:0] f1018_rst;
  logic [31:0] f1018_rdata;
  sr_buffer_32_1 f1018(.wen(f1018_wen), .wdata(f1018_wdata), .clk(f1018_clk), .rst(f1018_rst), .rdata(f1018_rdata));
  assign f1018_clk = clk;
  assign f1018_rst = rst;
  // Bindings to f1018

  // f1020
  logic [0:0] f1020_wen;
  logic [31:0] f1020_wdata;
  logic [0:0] f1020_clk;
  logic [0:0] f1020_rst;
  logic [31:0] f1020_rdata;
  sr_buffer_32_1 f1020(.wen(f1020_wen), .wdata(f1020_wdata), .clk(f1020_clk), .rst(f1020_rst), .rdata(f1020_rdata));
  assign f1020_clk = clk;
  assign f1020_rst = rst;
  // Bindings to f1020

  // f1022
  logic [0:0] f1022_wen;
  logic [31:0] f1022_wdata;
  logic [0:0] f1022_clk;
  logic [0:0] f1022_rst;
  logic [31:0] f1022_rdata;
  sr_buffer_32_1 f1022(.wen(f1022_wen), .wdata(f1022_wdata), .clk(f1022_clk), .rst(f1022_rst), .rdata(f1022_rdata));
  assign f1022_clk = clk;
  assign f1022_rst = rst;
  // Bindings to f1022

  // f1024
  logic [0:0] f1024_wen;
  logic [31:0] f1024_wdata;
  logic [0:0] f1024_clk;
  logic [0:0] f1024_rst;
  logic [31:0] f1024_rdata;
  sr_buffer_32_1 f1024(.wen(f1024_wen), .wdata(f1024_wdata), .clk(f1024_clk), .rst(f1024_rst), .rdata(f1024_rdata));
  assign f1024_clk = clk;
  assign f1024_rst = rst;
  // Bindings to f1024

  // f1026
  logic [0:0] f1026_wen;
  logic [31:0] f1026_wdata;
  logic [0:0] f1026_clk;
  logic [0:0] f1026_rst;
  logic [31:0] f1026_rdata;
  sr_buffer_32_1 f1026(.wen(f1026_wen), .wdata(f1026_wdata), .clk(f1026_clk), .rst(f1026_rst), .rdata(f1026_rdata));
  assign f1026_clk = clk;
  assign f1026_rst = rst;
  // Bindings to f1026

  // f1028
  logic [0:0] f1028_wen;
  logic [31:0] f1028_wdata;
  logic [0:0] f1028_clk;
  logic [0:0] f1028_rst;
  logic [31:0] f1028_rdata;
  sr_buffer_32_1 f1028(.wen(f1028_wen), .wdata(f1028_wdata), .clk(f1028_clk), .rst(f1028_rst), .rdata(f1028_rdata));
  assign f1028_clk = clk;
  assign f1028_rst = rst;
  // Bindings to f1028

  // f1030
  logic [0:0] f1030_wen;
  logic [31:0] f1030_wdata;
  logic [0:0] f1030_clk;
  logic [0:0] f1030_rst;
  logic [31:0] f1030_rdata;
  sr_buffer_32_1 f1030(.wen(f1030_wen), .wdata(f1030_wdata), .clk(f1030_clk), .rst(f1030_rst), .rdata(f1030_rdata));
  assign f1030_clk = clk;
  assign f1030_rst = rst;
  // Bindings to f1030

  // f1032
  logic [0:0] f1032_wen;
  logic [31:0] f1032_wdata;
  logic [0:0] f1032_clk;
  logic [0:0] f1032_rst;
  logic [31:0] f1032_rdata;
  sr_buffer_32_1 f1032(.wen(f1032_wen), .wdata(f1032_wdata), .clk(f1032_clk), .rst(f1032_rst), .rdata(f1032_rdata));
  assign f1032_clk = clk;
  assign f1032_rst = rst;
  // Bindings to f1032

  // f1034
  logic [0:0] f1034_wen;
  logic [31:0] f1034_wdata;
  logic [0:0] f1034_clk;
  logic [0:0] f1034_rst;
  logic [31:0] f1034_rdata;
  sr_buffer_32_1 f1034(.wen(f1034_wen), .wdata(f1034_wdata), .clk(f1034_clk), .rst(f1034_rst), .rdata(f1034_rdata));
  assign f1034_clk = clk;
  assign f1034_rst = rst;
  // Bindings to f1034

  // f1036
  logic [0:0] f1036_wen;
  logic [31:0] f1036_wdata;
  logic [0:0] f1036_clk;
  logic [0:0] f1036_rst;
  logic [31:0] f1036_rdata;
  sr_buffer_32_1 f1036(.wen(f1036_wen), .wdata(f1036_wdata), .clk(f1036_clk), .rst(f1036_rst), .rdata(f1036_rdata));
  assign f1036_clk = clk;
  assign f1036_rst = rst;
  // Bindings to f1036

  // f1038
  logic [0:0] f1038_wen;
  logic [31:0] f1038_wdata;
  logic [0:0] f1038_clk;
  logic [0:0] f1038_rst;
  logic [31:0] f1038_rdata;
  sr_buffer_32_1 f1038(.wen(f1038_wen), .wdata(f1038_wdata), .clk(f1038_clk), .rst(f1038_rst), .rdata(f1038_rdata));
  assign f1038_clk = clk;
  assign f1038_rst = rst;
  // Bindings to f1038

  // f1040
  logic [0:0] f1040_wen;
  logic [31:0] f1040_wdata;
  logic [0:0] f1040_clk;
  logic [0:0] f1040_rst;
  logic [31:0] f1040_rdata;
  sr_buffer_32_1 f1040(.wen(f1040_wen), .wdata(f1040_wdata), .clk(f1040_clk), .rst(f1040_rst), .rdata(f1040_rdata));
  assign f1040_clk = clk;
  assign f1040_rst = rst;
  // Bindings to f1040

  // f1042
  logic [0:0] f1042_wen;
  logic [31:0] f1042_wdata;
  logic [0:0] f1042_clk;
  logic [0:0] f1042_rst;
  logic [31:0] f1042_rdata;
  sr_buffer_32_1 f1042(.wen(f1042_wen), .wdata(f1042_wdata), .clk(f1042_clk), .rst(f1042_rst), .rdata(f1042_rdata));
  assign f1042_clk = clk;
  assign f1042_rst = rst;
  // Bindings to f1042

  // f1044
  logic [0:0] f1044_wen;
  logic [31:0] f1044_wdata;
  logic [0:0] f1044_clk;
  logic [0:0] f1044_rst;
  logic [31:0] f1044_rdata;
  sr_buffer_32_1 f1044(.wen(f1044_wen), .wdata(f1044_wdata), .clk(f1044_clk), .rst(f1044_rst), .rdata(f1044_rdata));
  assign f1044_clk = clk;
  assign f1044_rst = rst;
  // Bindings to f1044

  // f1046
  logic [0:0] f1046_wen;
  logic [31:0] f1046_wdata;
  logic [0:0] f1046_clk;
  logic [0:0] f1046_rst;
  logic [31:0] f1046_rdata;
  sr_buffer_32_1 f1046(.wen(f1046_wen), .wdata(f1046_wdata), .clk(f1046_clk), .rst(f1046_rst), .rdata(f1046_rdata));
  assign f1046_clk = clk;
  assign f1046_rst = rst;
  // Bindings to f1046

  // f1048
  logic [0:0] f1048_wen;
  logic [31:0] f1048_wdata;
  logic [0:0] f1048_clk;
  logic [0:0] f1048_rst;
  logic [31:0] f1048_rdata;
  sr_buffer_32_1 f1048(.wen(f1048_wen), .wdata(f1048_wdata), .clk(f1048_clk), .rst(f1048_rst), .rdata(f1048_rdata));
  assign f1048_clk = clk;
  assign f1048_rst = rst;
  // Bindings to f1048

  // f1050
  logic [0:0] f1050_wen;
  logic [31:0] f1050_wdata;
  logic [0:0] f1050_clk;
  logic [0:0] f1050_rst;
  logic [31:0] f1050_rdata;
  sr_buffer_32_1 f1050(.wen(f1050_wen), .wdata(f1050_wdata), .clk(f1050_clk), .rst(f1050_rst), .rdata(f1050_rdata));
  assign f1050_clk = clk;
  assign f1050_rst = rst;
  // Bindings to f1050

  // f1052
  logic [0:0] f1052_wen;
  logic [31:0] f1052_wdata;
  logic [0:0] f1052_clk;
  logic [0:0] f1052_rst;
  logic [31:0] f1052_rdata;
  sr_buffer_32_1 f1052(.wen(f1052_wen), .wdata(f1052_wdata), .clk(f1052_clk), .rst(f1052_rst), .rdata(f1052_rdata));
  assign f1052_clk = clk;
  assign f1052_rst = rst;
  // Bindings to f1052

  // f1054
  logic [0:0] f1054_wen;
  logic [31:0] f1054_wdata;
  logic [0:0] f1054_clk;
  logic [0:0] f1054_rst;
  logic [31:0] f1054_rdata;
  sr_buffer_32_1 f1054(.wen(f1054_wen), .wdata(f1054_wdata), .clk(f1054_clk), .rst(f1054_rst), .rdata(f1054_rdata));
  assign f1054_clk = clk;
  assign f1054_rst = rst;
  // Bindings to f1054

  // f1056
  logic [0:0] f1056_wen;
  logic [31:0] f1056_wdata;
  logic [0:0] f1056_clk;
  logic [0:0] f1056_rst;
  logic [31:0] f1056_rdata;
  sr_buffer_32_1 f1056(.wen(f1056_wen), .wdata(f1056_wdata), .clk(f1056_clk), .rst(f1056_rst), .rdata(f1056_rdata));
  assign f1056_clk = clk;
  assign f1056_rst = rst;
  // Bindings to f1056

  // f1058
  logic [0:0] f1058_wen;
  logic [31:0] f1058_wdata;
  logic [0:0] f1058_clk;
  logic [0:0] f1058_rst;
  logic [31:0] f1058_rdata;
  sr_buffer_32_1 f1058(.wen(f1058_wen), .wdata(f1058_wdata), .clk(f1058_clk), .rst(f1058_rst), .rdata(f1058_rdata));
  assign f1058_clk = clk;
  assign f1058_rst = rst;
  // Bindings to f1058

  // f1060
  logic [0:0] f1060_wen;
  logic [31:0] f1060_wdata;
  logic [0:0] f1060_clk;
  logic [0:0] f1060_rst;
  logic [31:0] f1060_rdata;
  sr_buffer_32_1 f1060(.wen(f1060_wen), .wdata(f1060_wdata), .clk(f1060_clk), .rst(f1060_rst), .rdata(f1060_rdata));
  assign f1060_clk = clk;
  assign f1060_rst = rst;
  // Bindings to f1060

  // f1062
  logic [0:0] f1062_wen;
  logic [31:0] f1062_wdata;
  logic [0:0] f1062_clk;
  logic [0:0] f1062_rst;
  logic [31:0] f1062_rdata;
  sr_buffer_32_1 f1062(.wen(f1062_wen), .wdata(f1062_wdata), .clk(f1062_clk), .rst(f1062_rst), .rdata(f1062_rdata));
  assign f1062_clk = clk;
  assign f1062_rst = rst;
  // Bindings to f1062

  // f1064
  logic [0:0] f1064_wen;
  logic [31:0] f1064_wdata;
  logic [0:0] f1064_clk;
  logic [0:0] f1064_rst;
  logic [31:0] f1064_rdata;
  sr_buffer_32_1 f1064(.wen(f1064_wen), .wdata(f1064_wdata), .clk(f1064_clk), .rst(f1064_rst), .rdata(f1064_rdata));
  assign f1064_clk = clk;
  assign f1064_rst = rst;
  // Bindings to f1064

  // f1066
  logic [0:0] f1066_wen;
  logic [31:0] f1066_wdata;
  logic [0:0] f1066_clk;
  logic [0:0] f1066_rst;
  logic [31:0] f1066_rdata;
  sr_buffer_32_1 f1066(.wen(f1066_wen), .wdata(f1066_wdata), .clk(f1066_clk), .rst(f1066_rst), .rdata(f1066_rdata));
  assign f1066_clk = clk;
  assign f1066_rst = rst;
  // Bindings to f1066

  // f1068
  logic [0:0] f1068_wen;
  logic [31:0] f1068_wdata;
  logic [0:0] f1068_clk;
  logic [0:0] f1068_rst;
  logic [31:0] f1068_rdata;
  sr_buffer_32_1 f1068(.wen(f1068_wen), .wdata(f1068_wdata), .clk(f1068_clk), .rst(f1068_rst), .rdata(f1068_rdata));
  assign f1068_clk = clk;
  assign f1068_rst = rst;
  // Bindings to f1068

  // f1070
  logic [0:0] f1070_wen;
  logic [31:0] f1070_wdata;
  logic [0:0] f1070_clk;
  logic [0:0] f1070_rst;
  logic [31:0] f1070_rdata;
  sr_buffer_32_1 f1070(.wen(f1070_wen), .wdata(f1070_wdata), .clk(f1070_clk), .rst(f1070_rst), .rdata(f1070_rdata));
  assign f1070_clk = clk;
  assign f1070_rst = rst;
  // Bindings to f1070

  // f1072
  logic [0:0] f1072_wen;
  logic [31:0] f1072_wdata;
  logic [0:0] f1072_clk;
  logic [0:0] f1072_rst;
  logic [31:0] f1072_rdata;
  sr_buffer_32_1 f1072(.wen(f1072_wen), .wdata(f1072_wdata), .clk(f1072_clk), .rst(f1072_rst), .rdata(f1072_rdata));
  assign f1072_clk = clk;
  assign f1072_rst = rst;
  // Bindings to f1072

  // f1074
  logic [0:0] f1074_wen;
  logic [31:0] f1074_wdata;
  logic [0:0] f1074_clk;
  logic [0:0] f1074_rst;
  logic [31:0] f1074_rdata;
  sr_buffer_32_1 f1074(.wen(f1074_wen), .wdata(f1074_wdata), .clk(f1074_clk), .rst(f1074_rst), .rdata(f1074_rdata));
  assign f1074_clk = clk;
  assign f1074_rst = rst;
  // Bindings to f1074

  // f1076
  logic [0:0] f1076_wen;
  logic [31:0] f1076_wdata;
  logic [0:0] f1076_clk;
  logic [0:0] f1076_rst;
  logic [31:0] f1076_rdata;
  sr_buffer_32_1 f1076(.wen(f1076_wen), .wdata(f1076_wdata), .clk(f1076_clk), .rst(f1076_rst), .rdata(f1076_rdata));
  assign f1076_clk = clk;
  assign f1076_rst = rst;
  // Bindings to f1076

  // f1078
  logic [0:0] f1078_wen;
  logic [31:0] f1078_wdata;
  logic [0:0] f1078_clk;
  logic [0:0] f1078_rst;
  logic [31:0] f1078_rdata;
  sr_buffer_32_1 f1078(.wen(f1078_wen), .wdata(f1078_wdata), .clk(f1078_clk), .rst(f1078_rst), .rdata(f1078_rdata));
  assign f1078_clk = clk;
  assign f1078_rst = rst;
  // Bindings to f1078

  // f1080
  logic [0:0] f1080_wen;
  logic [31:0] f1080_wdata;
  logic [0:0] f1080_clk;
  logic [0:0] f1080_rst;
  logic [31:0] f1080_rdata;
  sr_buffer_32_1 f1080(.wen(f1080_wen), .wdata(f1080_wdata), .clk(f1080_clk), .rst(f1080_rst), .rdata(f1080_rdata));
  assign f1080_clk = clk;
  assign f1080_rst = rst;
  // Bindings to f1080

  // f1082
  logic [0:0] f1082_wen;
  logic [31:0] f1082_wdata;
  logic [0:0] f1082_clk;
  logic [0:0] f1082_rst;
  logic [31:0] f1082_rdata;
  sr_buffer_32_1 f1082(.wen(f1082_wen), .wdata(f1082_wdata), .clk(f1082_clk), .rst(f1082_rst), .rdata(f1082_rdata));
  assign f1082_clk = clk;
  assign f1082_rst = rst;
  // Bindings to f1082

  // f1084
  logic [0:0] f1084_wen;
  logic [31:0] f1084_wdata;
  logic [0:0] f1084_clk;
  logic [0:0] f1084_rst;
  logic [31:0] f1084_rdata;
  sr_buffer_32_1 f1084(.wen(f1084_wen), .wdata(f1084_wdata), .clk(f1084_clk), .rst(f1084_rst), .rdata(f1084_rdata));
  assign f1084_clk = clk;
  assign f1084_rst = rst;
  // Bindings to f1084

  // f1086
  logic [0:0] f1086_wen;
  logic [31:0] f1086_wdata;
  logic [0:0] f1086_clk;
  logic [0:0] f1086_rst;
  logic [31:0] f1086_rdata;
  sr_buffer_32_1 f1086(.wen(f1086_wen), .wdata(f1086_wdata), .clk(f1086_clk), .rst(f1086_rst), .rdata(f1086_rdata));
  assign f1086_clk = clk;
  assign f1086_rst = rst;
  // Bindings to f1086

  // f1088
  logic [0:0] f1088_wen;
  logic [31:0] f1088_wdata;
  logic [0:0] f1088_clk;
  logic [0:0] f1088_rst;
  logic [31:0] f1088_rdata;
  sr_buffer_32_1 f1088(.wen(f1088_wen), .wdata(f1088_wdata), .clk(f1088_clk), .rst(f1088_rst), .rdata(f1088_rdata));
  assign f1088_clk = clk;
  assign f1088_rst = rst;
  // Bindings to f1088

  // f1090
  logic [0:0] f1090_wen;
  logic [31:0] f1090_wdata;
  logic [0:0] f1090_clk;
  logic [0:0] f1090_rst;
  logic [31:0] f1090_rdata;
  sr_buffer_32_1 f1090(.wen(f1090_wen), .wdata(f1090_wdata), .clk(f1090_clk), .rst(f1090_rst), .rdata(f1090_rdata));
  assign f1090_clk = clk;
  assign f1090_rst = rst;
  // Bindings to f1090

  // f1092
  logic [0:0] f1092_wen;
  logic [31:0] f1092_wdata;
  logic [0:0] f1092_clk;
  logic [0:0] f1092_rst;
  logic [31:0] f1092_rdata;
  sr_buffer_32_1 f1092(.wen(f1092_wen), .wdata(f1092_wdata), .clk(f1092_clk), .rst(f1092_rst), .rdata(f1092_rdata));
  assign f1092_clk = clk;
  assign f1092_rst = rst;
  // Bindings to f1092

  // f1094
  logic [0:0] f1094_wen;
  logic [31:0] f1094_wdata;
  logic [0:0] f1094_clk;
  logic [0:0] f1094_rst;
  logic [31:0] f1094_rdata;
  sr_buffer_32_1 f1094(.wen(f1094_wen), .wdata(f1094_wdata), .clk(f1094_clk), .rst(f1094_rst), .rdata(f1094_rdata));
  assign f1094_clk = clk;
  assign f1094_rst = rst;
  // Bindings to f1094

  // f1096
  logic [0:0] f1096_wen;
  logic [31:0] f1096_wdata;
  logic [0:0] f1096_clk;
  logic [0:0] f1096_rst;
  logic [31:0] f1096_rdata;
  sr_buffer_32_1 f1096(.wen(f1096_wen), .wdata(f1096_wdata), .clk(f1096_clk), .rst(f1096_rst), .rdata(f1096_rdata));
  assign f1096_clk = clk;
  assign f1096_rst = rst;
  // Bindings to f1096

  // f1098
  logic [0:0] f1098_wen;
  logic [31:0] f1098_wdata;
  logic [0:0] f1098_clk;
  logic [0:0] f1098_rst;
  logic [31:0] f1098_rdata;
  sr_buffer_32_1 f1098(.wen(f1098_wen), .wdata(f1098_wdata), .clk(f1098_clk), .rst(f1098_rst), .rdata(f1098_rdata));
  assign f1098_clk = clk;
  assign f1098_rst = rst;
  // Bindings to f1098

  // f1100
  logic [0:0] f1100_wen;
  logic [31:0] f1100_wdata;
  logic [0:0] f1100_clk;
  logic [0:0] f1100_rst;
  logic [31:0] f1100_rdata;
  sr_buffer_32_1 f1100(.wen(f1100_wen), .wdata(f1100_wdata), .clk(f1100_clk), .rst(f1100_rst), .rdata(f1100_rdata));
  assign f1100_clk = clk;
  assign f1100_rst = rst;
  // Bindings to f1100

  // f1102
  logic [0:0] f1102_wen;
  logic [31:0] f1102_wdata;
  logic [0:0] f1102_clk;
  logic [0:0] f1102_rst;
  logic [31:0] f1102_rdata;
  sr_buffer_32_1 f1102(.wen(f1102_wen), .wdata(f1102_wdata), .clk(f1102_clk), .rst(f1102_rst), .rdata(f1102_rdata));
  assign f1102_clk = clk;
  assign f1102_rst = rst;
  // Bindings to f1102

  // f1104
  logic [0:0] f1104_wen;
  logic [31:0] f1104_wdata;
  logic [0:0] f1104_clk;
  logic [0:0] f1104_rst;
  logic [31:0] f1104_rdata;
  sr_buffer_32_1 f1104(.wen(f1104_wen), .wdata(f1104_wdata), .clk(f1104_clk), .rst(f1104_rst), .rdata(f1104_rdata));
  assign f1104_clk = clk;
  assign f1104_rst = rst;
  // Bindings to f1104

  // f1106
  logic [0:0] f1106_wen;
  logic [31:0] f1106_wdata;
  logic [0:0] f1106_clk;
  logic [0:0] f1106_rst;
  logic [31:0] f1106_rdata;
  sr_buffer_32_1 f1106(.wen(f1106_wen), .wdata(f1106_wdata), .clk(f1106_clk), .rst(f1106_rst), .rdata(f1106_rdata));
  assign f1106_clk = clk;
  assign f1106_rst = rst;
  // Bindings to f1106

  // f1108
  logic [0:0] f1108_wen;
  logic [31:0] f1108_wdata;
  logic [0:0] f1108_clk;
  logic [0:0] f1108_rst;
  logic [31:0] f1108_rdata;
  sr_buffer_32_1 f1108(.wen(f1108_wen), .wdata(f1108_wdata), .clk(f1108_clk), .rst(f1108_rst), .rdata(f1108_rdata));
  assign f1108_clk = clk;
  assign f1108_rst = rst;
  // Bindings to f1108

  // f1110
  logic [0:0] f1110_wen;
  logic [31:0] f1110_wdata;
  logic [0:0] f1110_clk;
  logic [0:0] f1110_rst;
  logic [31:0] f1110_rdata;
  sr_buffer_32_1 f1110(.wen(f1110_wen), .wdata(f1110_wdata), .clk(f1110_clk), .rst(f1110_rst), .rdata(f1110_rdata));
  assign f1110_clk = clk;
  assign f1110_rst = rst;
  // Bindings to f1110

  // f1112
  logic [0:0] f1112_wen;
  logic [31:0] f1112_wdata;
  logic [0:0] f1112_clk;
  logic [0:0] f1112_rst;
  logic [31:0] f1112_rdata;
  sr_buffer_32_1 f1112(.wen(f1112_wen), .wdata(f1112_wdata), .clk(f1112_clk), .rst(f1112_rst), .rdata(f1112_rdata));
  assign f1112_clk = clk;
  assign f1112_rst = rst;
  // Bindings to f1112

  // f1114
  logic [0:0] f1114_wen;
  logic [31:0] f1114_wdata;
  logic [0:0] f1114_clk;
  logic [0:0] f1114_rst;
  logic [31:0] f1114_rdata;
  sr_buffer_32_1 f1114(.wen(f1114_wen), .wdata(f1114_wdata), .clk(f1114_clk), .rst(f1114_rst), .rdata(f1114_rdata));
  assign f1114_clk = clk;
  assign f1114_rst = rst;
  // Bindings to f1114

  // f1116
  logic [0:0] f1116_wen;
  logic [31:0] f1116_wdata;
  logic [0:0] f1116_clk;
  logic [0:0] f1116_rst;
  logic [31:0] f1116_rdata;
  sr_buffer_32_1 f1116(.wen(f1116_wen), .wdata(f1116_wdata), .clk(f1116_clk), .rst(f1116_rst), .rdata(f1116_rdata));
  assign f1116_clk = clk;
  assign f1116_rst = rst;
  // Bindings to f1116

  // f1118
  logic [0:0] f1118_wen;
  logic [31:0] f1118_wdata;
  logic [0:0] f1118_clk;
  logic [0:0] f1118_rst;
  logic [31:0] f1118_rdata;
  sr_buffer_32_1 f1118(.wen(f1118_wen), .wdata(f1118_wdata), .clk(f1118_clk), .rst(f1118_rst), .rdata(f1118_rdata));
  assign f1118_clk = clk;
  assign f1118_rst = rst;
  // Bindings to f1118

  // f1120
  logic [0:0] f1120_wen;
  logic [31:0] f1120_wdata;
  logic [0:0] f1120_clk;
  logic [0:0] f1120_rst;
  logic [31:0] f1120_rdata;
  sr_buffer_32_1 f1120(.wen(f1120_wen), .wdata(f1120_wdata), .clk(f1120_clk), .rst(f1120_rst), .rdata(f1120_rdata));
  assign f1120_clk = clk;
  assign f1120_rst = rst;
  // Bindings to f1120

  // f1122
  logic [0:0] f1122_wen;
  logic [31:0] f1122_wdata;
  logic [0:0] f1122_clk;
  logic [0:0] f1122_rst;
  logic [31:0] f1122_rdata;
  sr_buffer_32_1 f1122(.wen(f1122_wen), .wdata(f1122_wdata), .clk(f1122_clk), .rst(f1122_rst), .rdata(f1122_rdata));
  assign f1122_clk = clk;
  assign f1122_rst = rst;
  // Bindings to f1122

  // f1124
  logic [0:0] f1124_wen;
  logic [31:0] f1124_wdata;
  logic [0:0] f1124_clk;
  logic [0:0] f1124_rst;
  logic [31:0] f1124_rdata;
  sr_buffer_32_1 f1124(.wen(f1124_wen), .wdata(f1124_wdata), .clk(f1124_clk), .rst(f1124_rst), .rdata(f1124_rdata));
  assign f1124_clk = clk;
  assign f1124_rst = rst;
  // Bindings to f1124

  // f1126
  logic [0:0] f1126_wen;
  logic [31:0] f1126_wdata;
  logic [0:0] f1126_clk;
  logic [0:0] f1126_rst;
  logic [31:0] f1126_rdata;
  sr_buffer_32_1 f1126(.wen(f1126_wen), .wdata(f1126_wdata), .clk(f1126_clk), .rst(f1126_rst), .rdata(f1126_rdata));
  assign f1126_clk = clk;
  assign f1126_rst = rst;
  // Bindings to f1126

  // f1128
  logic [0:0] f1128_wen;
  logic [31:0] f1128_wdata;
  logic [0:0] f1128_clk;
  logic [0:0] f1128_rst;
  logic [31:0] f1128_rdata;
  sr_buffer_32_1 f1128(.wen(f1128_wen), .wdata(f1128_wdata), .clk(f1128_clk), .rst(f1128_rst), .rdata(f1128_rdata));
  assign f1128_clk = clk;
  assign f1128_rst = rst;
  // Bindings to f1128

  // f1130
  logic [0:0] f1130_wen;
  logic [31:0] f1130_wdata;
  logic [0:0] f1130_clk;
  logic [0:0] f1130_rst;
  logic [31:0] f1130_rdata;
  sr_buffer_32_1 f1130(.wen(f1130_wen), .wdata(f1130_wdata), .clk(f1130_clk), .rst(f1130_rst), .rdata(f1130_rdata));
  assign f1130_clk = clk;
  assign f1130_rst = rst;
  // Bindings to f1130

  // f1132
  logic [0:0] f1132_wen;
  logic [31:0] f1132_wdata;
  logic [0:0] f1132_clk;
  logic [0:0] f1132_rst;
  logic [31:0] f1132_rdata;
  sr_buffer_32_1 f1132(.wen(f1132_wen), .wdata(f1132_wdata), .clk(f1132_clk), .rst(f1132_rst), .rdata(f1132_rdata));
  assign f1132_clk = clk;
  assign f1132_rst = rst;
  // Bindings to f1132

  // f1134
  logic [0:0] f1134_wen;
  logic [31:0] f1134_wdata;
  logic [0:0] f1134_clk;
  logic [0:0] f1134_rst;
  logic [31:0] f1134_rdata;
  sr_buffer_32_1 f1134(.wen(f1134_wen), .wdata(f1134_wdata), .clk(f1134_clk), .rst(f1134_rst), .rdata(f1134_rdata));
  assign f1134_clk = clk;
  assign f1134_rst = rst;
  // Bindings to f1134

  // f1136
  logic [0:0] f1136_wen;
  logic [31:0] f1136_wdata;
  logic [0:0] f1136_clk;
  logic [0:0] f1136_rst;
  logic [31:0] f1136_rdata;
  sr_buffer_32_1 f1136(.wen(f1136_wen), .wdata(f1136_wdata), .clk(f1136_clk), .rst(f1136_rst), .rdata(f1136_rdata));
  assign f1136_clk = clk;
  assign f1136_rst = rst;
  // Bindings to f1136

  // f1138
  logic [0:0] f1138_wen;
  logic [31:0] f1138_wdata;
  logic [0:0] f1138_clk;
  logic [0:0] f1138_rst;
  logic [31:0] f1138_rdata;
  sr_buffer_32_1 f1138(.wen(f1138_wen), .wdata(f1138_wdata), .clk(f1138_clk), .rst(f1138_rst), .rdata(f1138_rdata));
  assign f1138_clk = clk;
  assign f1138_rst = rst;
  // Bindings to f1138

  // f1140
  logic [0:0] f1140_wen;
  logic [31:0] f1140_wdata;
  logic [0:0] f1140_clk;
  logic [0:0] f1140_rst;
  logic [31:0] f1140_rdata;
  sr_buffer_32_1 f1140(.wen(f1140_wen), .wdata(f1140_wdata), .clk(f1140_clk), .rst(f1140_rst), .rdata(f1140_rdata));
  assign f1140_clk = clk;
  assign f1140_rst = rst;
  // Bindings to f1140

  // f1142
  logic [0:0] f1142_wen;
  logic [31:0] f1142_wdata;
  logic [0:0] f1142_clk;
  logic [0:0] f1142_rst;
  logic [31:0] f1142_rdata;
  sr_buffer_32_1 f1142(.wen(f1142_wen), .wdata(f1142_wdata), .clk(f1142_clk), .rst(f1142_rst), .rdata(f1142_rdata));
  assign f1142_clk = clk;
  assign f1142_rst = rst;
  // Bindings to f1142

  // f1144
  logic [0:0] f1144_wen;
  logic [31:0] f1144_wdata;
  logic [0:0] f1144_clk;
  logic [0:0] f1144_rst;
  logic [31:0] f1144_rdata;
  sr_buffer_32_1 f1144(.wen(f1144_wen), .wdata(f1144_wdata), .clk(f1144_clk), .rst(f1144_rst), .rdata(f1144_rdata));
  assign f1144_clk = clk;
  assign f1144_rst = rst;
  // Bindings to f1144

  // f1146
  logic [0:0] f1146_wen;
  logic [31:0] f1146_wdata;
  logic [0:0] f1146_clk;
  logic [0:0] f1146_rst;
  logic [31:0] f1146_rdata;
  sr_buffer_32_1 f1146(.wen(f1146_wen), .wdata(f1146_wdata), .clk(f1146_clk), .rst(f1146_rst), .rdata(f1146_rdata));
  assign f1146_clk = clk;
  assign f1146_rst = rst;
  // Bindings to f1146

  // f1148
  logic [0:0] f1148_wen;
  logic [31:0] f1148_wdata;
  logic [0:0] f1148_clk;
  logic [0:0] f1148_rst;
  logic [31:0] f1148_rdata;
  sr_buffer_32_1 f1148(.wen(f1148_wen), .wdata(f1148_wdata), .clk(f1148_clk), .rst(f1148_rst), .rdata(f1148_rdata));
  assign f1148_clk = clk;
  assign f1148_rst = rst;
  // Bindings to f1148

  // f1150
  logic [0:0] f1150_wen;
  logic [31:0] f1150_wdata;
  logic [0:0] f1150_clk;
  logic [0:0] f1150_rst;
  logic [31:0] f1150_rdata;
  sr_buffer_32_1 f1150(.wen(f1150_wen), .wdata(f1150_wdata), .clk(f1150_clk), .rst(f1150_rst), .rdata(f1150_rdata));
  assign f1150_clk = clk;
  assign f1150_rst = rst;
  // Bindings to f1150

  // f1152
  logic [0:0] f1152_wen;
  logic [31:0] f1152_wdata;
  logic [0:0] f1152_clk;
  logic [0:0] f1152_rst;
  logic [31:0] f1152_rdata;
  sr_buffer_32_1 f1152(.wen(f1152_wen), .wdata(f1152_wdata), .clk(f1152_clk), .rst(f1152_rst), .rdata(f1152_rdata));
  assign f1152_clk = clk;
  assign f1152_rst = rst;
  // Bindings to f1152

  // f1154
  logic [0:0] f1154_wen;
  logic [31:0] f1154_wdata;
  logic [0:0] f1154_clk;
  logic [0:0] f1154_rst;
  logic [31:0] f1154_rdata;
  sr_buffer_32_1 f1154(.wen(f1154_wen), .wdata(f1154_wdata), .clk(f1154_clk), .rst(f1154_rst), .rdata(f1154_rdata));
  assign f1154_clk = clk;
  assign f1154_rst = rst;
  // Bindings to f1154

  // f1156
  logic [0:0] f1156_wen;
  logic [31:0] f1156_wdata;
  logic [0:0] f1156_clk;
  logic [0:0] f1156_rst;
  logic [31:0] f1156_rdata;
  sr_buffer_32_1 f1156(.wen(f1156_wen), .wdata(f1156_wdata), .clk(f1156_clk), .rst(f1156_rst), .rdata(f1156_rdata));
  assign f1156_clk = clk;
  assign f1156_rst = rst;
  // Bindings to f1156

  // f1158
  logic [0:0] f1158_wen;
  logic [31:0] f1158_wdata;
  logic [0:0] f1158_clk;
  logic [0:0] f1158_rst;
  logic [31:0] f1158_rdata;
  sr_buffer_32_1 f1158(.wen(f1158_wen), .wdata(f1158_wdata), .clk(f1158_clk), .rst(f1158_rst), .rdata(f1158_rdata));
  assign f1158_clk = clk;
  assign f1158_rst = rst;
  // Bindings to f1158

  // f1160
  logic [0:0] f1160_wen;
  logic [31:0] f1160_wdata;
  logic [0:0] f1160_clk;
  logic [0:0] f1160_rst;
  logic [31:0] f1160_rdata;
  sr_buffer_32_1 f1160(.wen(f1160_wen), .wdata(f1160_wdata), .clk(f1160_clk), .rst(f1160_rst), .rdata(f1160_rdata));
  assign f1160_clk = clk;
  assign f1160_rst = rst;
  // Bindings to f1160

  // f1162
  logic [0:0] f1162_wen;
  logic [31:0] f1162_wdata;
  logic [0:0] f1162_clk;
  logic [0:0] f1162_rst;
  logic [31:0] f1162_rdata;
  sr_buffer_32_1 f1162(.wen(f1162_wen), .wdata(f1162_wdata), .clk(f1162_clk), .rst(f1162_rst), .rdata(f1162_rdata));
  assign f1162_clk = clk;
  assign f1162_rst = rst;
  // Bindings to f1162

  // f1164
  logic [0:0] f1164_wen;
  logic [31:0] f1164_wdata;
  logic [0:0] f1164_clk;
  logic [0:0] f1164_rst;
  logic [31:0] f1164_rdata;
  sr_buffer_32_1 f1164(.wen(f1164_wen), .wdata(f1164_wdata), .clk(f1164_clk), .rst(f1164_rst), .rdata(f1164_rdata));
  assign f1164_clk = clk;
  assign f1164_rst = rst;
  // Bindings to f1164

  // f1166
  logic [0:0] f1166_wen;
  logic [31:0] f1166_wdata;
  logic [0:0] f1166_clk;
  logic [0:0] f1166_rst;
  logic [31:0] f1166_rdata;
  sr_buffer_32_1 f1166(.wen(f1166_wen), .wdata(f1166_wdata), .clk(f1166_clk), .rst(f1166_rst), .rdata(f1166_rdata));
  assign f1166_clk = clk;
  assign f1166_rst = rst;
  // Bindings to f1166

  // f1168
  logic [0:0] f1168_wen;
  logic [31:0] f1168_wdata;
  logic [0:0] f1168_clk;
  logic [0:0] f1168_rst;
  logic [31:0] f1168_rdata;
  sr_buffer_32_1 f1168(.wen(f1168_wen), .wdata(f1168_wdata), .clk(f1168_clk), .rst(f1168_rst), .rdata(f1168_rdata));
  assign f1168_clk = clk;
  assign f1168_rst = rst;
  // Bindings to f1168

  // f1170
  logic [0:0] f1170_wen;
  logic [31:0] f1170_wdata;
  logic [0:0] f1170_clk;
  logic [0:0] f1170_rst;
  logic [31:0] f1170_rdata;
  sr_buffer_32_1 f1170(.wen(f1170_wen), .wdata(f1170_wdata), .clk(f1170_clk), .rst(f1170_rst), .rdata(f1170_rdata));
  assign f1170_clk = clk;
  assign f1170_rst = rst;
  // Bindings to f1170

  // f1172
  logic [0:0] f1172_wen;
  logic [31:0] f1172_wdata;
  logic [0:0] f1172_clk;
  logic [0:0] f1172_rst;
  logic [31:0] f1172_rdata;
  sr_buffer_32_1 f1172(.wen(f1172_wen), .wdata(f1172_wdata), .clk(f1172_clk), .rst(f1172_rst), .rdata(f1172_rdata));
  assign f1172_clk = clk;
  assign f1172_rst = rst;
  // Bindings to f1172

  // f1174
  logic [0:0] f1174_wen;
  logic [31:0] f1174_wdata;
  logic [0:0] f1174_clk;
  logic [0:0] f1174_rst;
  logic [31:0] f1174_rdata;
  sr_buffer_32_1 f1174(.wen(f1174_wen), .wdata(f1174_wdata), .clk(f1174_clk), .rst(f1174_rst), .rdata(f1174_rdata));
  assign f1174_clk = clk;
  assign f1174_rst = rst;
  // Bindings to f1174

  // f1176
  logic [0:0] f1176_wen;
  logic [31:0] f1176_wdata;
  logic [0:0] f1176_clk;
  logic [0:0] f1176_rst;
  logic [31:0] f1176_rdata;
  sr_buffer_32_1 f1176(.wen(f1176_wen), .wdata(f1176_wdata), .clk(f1176_clk), .rst(f1176_rst), .rdata(f1176_rdata));
  assign f1176_clk = clk;
  assign f1176_rst = rst;
  // Bindings to f1176

  // f1178
  logic [0:0] f1178_wen;
  logic [31:0] f1178_wdata;
  logic [0:0] f1178_clk;
  logic [0:0] f1178_rst;
  logic [31:0] f1178_rdata;
  sr_buffer_32_1 f1178(.wen(f1178_wen), .wdata(f1178_wdata), .clk(f1178_clk), .rst(f1178_rst), .rdata(f1178_rdata));
  assign f1178_clk = clk;
  assign f1178_rst = rst;
  // Bindings to f1178

  // f1180
  logic [0:0] f1180_wen;
  logic [31:0] f1180_wdata;
  logic [0:0] f1180_clk;
  logic [0:0] f1180_rst;
  logic [31:0] f1180_rdata;
  sr_buffer_32_1 f1180(.wen(f1180_wen), .wdata(f1180_wdata), .clk(f1180_clk), .rst(f1180_rst), .rdata(f1180_rdata));
  assign f1180_clk = clk;
  assign f1180_rst = rst;
  // Bindings to f1180

  // f1182
  logic [0:0] f1182_wen;
  logic [31:0] f1182_wdata;
  logic [0:0] f1182_clk;
  logic [0:0] f1182_rst;
  logic [31:0] f1182_rdata;
  sr_buffer_32_1 f1182(.wen(f1182_wen), .wdata(f1182_wdata), .clk(f1182_clk), .rst(f1182_rst), .rdata(f1182_rdata));
  assign f1182_clk = clk;
  assign f1182_rst = rst;
  // Bindings to f1182

  // f1184
  logic [0:0] f1184_wen;
  logic [31:0] f1184_wdata;
  logic [0:0] f1184_clk;
  logic [0:0] f1184_rst;
  logic [31:0] f1184_rdata;
  sr_buffer_32_1 f1184(.wen(f1184_wen), .wdata(f1184_wdata), .clk(f1184_clk), .rst(f1184_rst), .rdata(f1184_rdata));
  assign f1184_clk = clk;
  assign f1184_rst = rst;
  // Bindings to f1184

  // f1186
  logic [0:0] f1186_wen;
  logic [31:0] f1186_wdata;
  logic [0:0] f1186_clk;
  logic [0:0] f1186_rst;
  logic [31:0] f1186_rdata;
  sr_buffer_32_1 f1186(.wen(f1186_wen), .wdata(f1186_wdata), .clk(f1186_clk), .rst(f1186_rst), .rdata(f1186_rdata));
  assign f1186_clk = clk;
  assign f1186_rst = rst;
  // Bindings to f1186

  // f1188
  logic [0:0] f1188_wen;
  logic [31:0] f1188_wdata;
  logic [0:0] f1188_clk;
  logic [0:0] f1188_rst;
  logic [31:0] f1188_rdata;
  sr_buffer_32_1 f1188(.wen(f1188_wen), .wdata(f1188_wdata), .clk(f1188_clk), .rst(f1188_rst), .rdata(f1188_rdata));
  assign f1188_clk = clk;
  assign f1188_rst = rst;
  // Bindings to f1188

  // f1190
  logic [0:0] f1190_wen;
  logic [31:0] f1190_wdata;
  logic [0:0] f1190_clk;
  logic [0:0] f1190_rst;
  logic [31:0] f1190_rdata;
  sr_buffer_32_1 f1190(.wen(f1190_wen), .wdata(f1190_wdata), .clk(f1190_clk), .rst(f1190_rst), .rdata(f1190_rdata));
  assign f1190_clk = clk;
  assign f1190_rst = rst;
  // Bindings to f1190

  // f1192
  logic [0:0] f1192_wen;
  logic [31:0] f1192_wdata;
  logic [0:0] f1192_clk;
  logic [0:0] f1192_rst;
  logic [31:0] f1192_rdata;
  sr_buffer_32_1 f1192(.wen(f1192_wen), .wdata(f1192_wdata), .clk(f1192_clk), .rst(f1192_rst), .rdata(f1192_rdata));
  assign f1192_clk = clk;
  assign f1192_rst = rst;
  // Bindings to f1192

  // f1194
  logic [0:0] f1194_wen;
  logic [31:0] f1194_wdata;
  logic [0:0] f1194_clk;
  logic [0:0] f1194_rst;
  logic [31:0] f1194_rdata;
  sr_buffer_32_1 f1194(.wen(f1194_wen), .wdata(f1194_wdata), .clk(f1194_clk), .rst(f1194_rst), .rdata(f1194_rdata));
  assign f1194_clk = clk;
  assign f1194_rst = rst;
  // Bindings to f1194

  // f1196
  logic [0:0] f1196_wen;
  logic [31:0] f1196_wdata;
  logic [0:0] f1196_clk;
  logic [0:0] f1196_rst;
  logic [31:0] f1196_rdata;
  sr_buffer_32_1 f1196(.wen(f1196_wen), .wdata(f1196_wdata), .clk(f1196_clk), .rst(f1196_rst), .rdata(f1196_rdata));
  assign f1196_clk = clk;
  assign f1196_rst = rst;
  // Bindings to f1196

  // f1198
  logic [0:0] f1198_wen;
  logic [31:0] f1198_wdata;
  logic [0:0] f1198_clk;
  logic [0:0] f1198_rst;
  logic [31:0] f1198_rdata;
  sr_buffer_32_1 f1198(.wen(f1198_wen), .wdata(f1198_wdata), .clk(f1198_clk), .rst(f1198_rst), .rdata(f1198_rdata));
  assign f1198_clk = clk;
  assign f1198_rst = rst;
  // Bindings to f1198

  // f1200
  logic [0:0] f1200_wen;
  logic [31:0] f1200_wdata;
  logic [0:0] f1200_clk;
  logic [0:0] f1200_rst;
  logic [31:0] f1200_rdata;
  sr_buffer_32_1 f1200(.wen(f1200_wen), .wdata(f1200_wdata), .clk(f1200_clk), .rst(f1200_rst), .rdata(f1200_rdata));
  assign f1200_clk = clk;
  assign f1200_rst = rst;
  // Bindings to f1200

  // f1202
  logic [0:0] f1202_wen;
  logic [31:0] f1202_wdata;
  logic [0:0] f1202_clk;
  logic [0:0] f1202_rst;
  logic [31:0] f1202_rdata;
  sr_buffer_32_1 f1202(.wen(f1202_wen), .wdata(f1202_wdata), .clk(f1202_clk), .rst(f1202_rst), .rdata(f1202_rdata));
  assign f1202_clk = clk;
  assign f1202_rst = rst;
  // Bindings to f1202

  // f1204
  logic [0:0] f1204_wen;
  logic [31:0] f1204_wdata;
  logic [0:0] f1204_clk;
  logic [0:0] f1204_rst;
  logic [31:0] f1204_rdata;
  sr_buffer_32_1 f1204(.wen(f1204_wen), .wdata(f1204_wdata), .clk(f1204_clk), .rst(f1204_rst), .rdata(f1204_rdata));
  assign f1204_clk = clk;
  assign f1204_rst = rst;
  // Bindings to f1204

  // f1206
  logic [0:0] f1206_wen;
  logic [31:0] f1206_wdata;
  logic [0:0] f1206_clk;
  logic [0:0] f1206_rst;
  logic [31:0] f1206_rdata;
  sr_buffer_32_1 f1206(.wen(f1206_wen), .wdata(f1206_wdata), .clk(f1206_clk), .rst(f1206_rst), .rdata(f1206_rdata));
  assign f1206_clk = clk;
  assign f1206_rst = rst;
  // Bindings to f1206

  // f1208
  logic [0:0] f1208_wen;
  logic [31:0] f1208_wdata;
  logic [0:0] f1208_clk;
  logic [0:0] f1208_rst;
  logic [31:0] f1208_rdata;
  sr_buffer_32_1 f1208(.wen(f1208_wen), .wdata(f1208_wdata), .clk(f1208_clk), .rst(f1208_rst), .rdata(f1208_rdata));
  assign f1208_clk = clk;
  assign f1208_rst = rst;
  // Bindings to f1208

  // f1210
  logic [0:0] f1210_wen;
  logic [31:0] f1210_wdata;
  logic [0:0] f1210_clk;
  logic [0:0] f1210_rst;
  logic [31:0] f1210_rdata;
  sr_buffer_32_1 f1210(.wen(f1210_wen), .wdata(f1210_wdata), .clk(f1210_clk), .rst(f1210_rst), .rdata(f1210_rdata));
  assign f1210_clk = clk;
  assign f1210_rst = rst;
  // Bindings to f1210

  // f1212
  logic [0:0] f1212_wen;
  logic [31:0] f1212_wdata;
  logic [0:0] f1212_clk;
  logic [0:0] f1212_rst;
  logic [31:0] f1212_rdata;
  sr_buffer_32_1 f1212(.wen(f1212_wen), .wdata(f1212_wdata), .clk(f1212_clk), .rst(f1212_rst), .rdata(f1212_rdata));
  assign f1212_clk = clk;
  assign f1212_rst = rst;
  // Bindings to f1212

  // f1214
  logic [0:0] f1214_wen;
  logic [31:0] f1214_wdata;
  logic [0:0] f1214_clk;
  logic [0:0] f1214_rst;
  logic [31:0] f1214_rdata;
  sr_buffer_32_1 f1214(.wen(f1214_wen), .wdata(f1214_wdata), .clk(f1214_clk), .rst(f1214_rst), .rdata(f1214_rdata));
  assign f1214_clk = clk;
  assign f1214_rst = rst;
  // Bindings to f1214

  // f1216
  logic [0:0] f1216_wen;
  logic [31:0] f1216_wdata;
  logic [0:0] f1216_clk;
  logic [0:0] f1216_rst;
  logic [31:0] f1216_rdata;
  sr_buffer_32_1 f1216(.wen(f1216_wen), .wdata(f1216_wdata), .clk(f1216_clk), .rst(f1216_rst), .rdata(f1216_rdata));
  assign f1216_clk = clk;
  assign f1216_rst = rst;
  // Bindings to f1216

  // f1218
  logic [0:0] f1218_wen;
  logic [31:0] f1218_wdata;
  logic [0:0] f1218_clk;
  logic [0:0] f1218_rst;
  logic [31:0] f1218_rdata;
  sr_buffer_32_1 f1218(.wen(f1218_wen), .wdata(f1218_wdata), .clk(f1218_clk), .rst(f1218_rst), .rdata(f1218_rdata));
  assign f1218_clk = clk;
  assign f1218_rst = rst;
  // Bindings to f1218

  // f1220
  logic [0:0] f1220_wen;
  logic [31:0] f1220_wdata;
  logic [0:0] f1220_clk;
  logic [0:0] f1220_rst;
  logic [31:0] f1220_rdata;
  sr_buffer_32_1 f1220(.wen(f1220_wen), .wdata(f1220_wdata), .clk(f1220_clk), .rst(f1220_rst), .rdata(f1220_rdata));
  assign f1220_clk = clk;
  assign f1220_rst = rst;
  // Bindings to f1220

  // f1222
  logic [0:0] f1222_wen;
  logic [31:0] f1222_wdata;
  logic [0:0] f1222_clk;
  logic [0:0] f1222_rst;
  logic [31:0] f1222_rdata;
  sr_buffer_32_1 f1222(.wen(f1222_wen), .wdata(f1222_wdata), .clk(f1222_clk), .rst(f1222_rst), .rdata(f1222_rdata));
  assign f1222_clk = clk;
  assign f1222_rst = rst;
  // Bindings to f1222

  // f1224
  logic [0:0] f1224_wen;
  logic [31:0] f1224_wdata;
  logic [0:0] f1224_clk;
  logic [0:0] f1224_rst;
  logic [31:0] f1224_rdata;
  sr_buffer_32_1 f1224(.wen(f1224_wen), .wdata(f1224_wdata), .clk(f1224_clk), .rst(f1224_rst), .rdata(f1224_rdata));
  assign f1224_clk = clk;
  assign f1224_rst = rst;
  // Bindings to f1224

  // f1226
  logic [0:0] f1226_wen;
  logic [31:0] f1226_wdata;
  logic [0:0] f1226_clk;
  logic [0:0] f1226_rst;
  logic [31:0] f1226_rdata;
  sr_buffer_32_1 f1226(.wen(f1226_wen), .wdata(f1226_wdata), .clk(f1226_clk), .rst(f1226_rst), .rdata(f1226_rdata));
  assign f1226_clk = clk;
  assign f1226_rst = rst;
  // Bindings to f1226

  // f1228
  logic [0:0] f1228_wen;
  logic [31:0] f1228_wdata;
  logic [0:0] f1228_clk;
  logic [0:0] f1228_rst;
  logic [31:0] f1228_rdata;
  sr_buffer_32_1 f1228(.wen(f1228_wen), .wdata(f1228_wdata), .clk(f1228_clk), .rst(f1228_rst), .rdata(f1228_rdata));
  assign f1228_clk = clk;
  assign f1228_rst = rst;
  // Bindings to f1228

  // f1230
  logic [0:0] f1230_wen;
  logic [31:0] f1230_wdata;
  logic [0:0] f1230_clk;
  logic [0:0] f1230_rst;
  logic [31:0] f1230_rdata;
  sr_buffer_32_1 f1230(.wen(f1230_wen), .wdata(f1230_wdata), .clk(f1230_clk), .rst(f1230_rst), .rdata(f1230_rdata));
  assign f1230_clk = clk;
  assign f1230_rst = rst;
  // Bindings to f1230

  // f1232
  logic [0:0] f1232_wen;
  logic [31:0] f1232_wdata;
  logic [0:0] f1232_clk;
  logic [0:0] f1232_rst;
  logic [31:0] f1232_rdata;
  sr_buffer_32_1 f1232(.wen(f1232_wen), .wdata(f1232_wdata), .clk(f1232_clk), .rst(f1232_rst), .rdata(f1232_rdata));
  assign f1232_clk = clk;
  assign f1232_rst = rst;
  // Bindings to f1232

  // f1234
  logic [0:0] f1234_wen;
  logic [31:0] f1234_wdata;
  logic [0:0] f1234_clk;
  logic [0:0] f1234_rst;
  logic [31:0] f1234_rdata;
  sr_buffer_32_1 f1234(.wen(f1234_wen), .wdata(f1234_wdata), .clk(f1234_clk), .rst(f1234_rst), .rdata(f1234_rdata));
  assign f1234_clk = clk;
  assign f1234_rst = rst;
  // Bindings to f1234

  // f1236
  logic [0:0] f1236_wen;
  logic [31:0] f1236_wdata;
  logic [0:0] f1236_clk;
  logic [0:0] f1236_rst;
  logic [31:0] f1236_rdata;
  sr_buffer_32_1 f1236(.wen(f1236_wen), .wdata(f1236_wdata), .clk(f1236_clk), .rst(f1236_rst), .rdata(f1236_rdata));
  assign f1236_clk = clk;
  assign f1236_rst = rst;
  // Bindings to f1236

  // f1238
  logic [0:0] f1238_wen;
  logic [31:0] f1238_wdata;
  logic [0:0] f1238_clk;
  logic [0:0] f1238_rst;
  logic [31:0] f1238_rdata;
  sr_buffer_32_1 f1238(.wen(f1238_wen), .wdata(f1238_wdata), .clk(f1238_clk), .rst(f1238_rst), .rdata(f1238_rdata));
  assign f1238_clk = clk;
  assign f1238_rst = rst;
  // Bindings to f1238

  // f1240
  logic [0:0] f1240_wen;
  logic [31:0] f1240_wdata;
  logic [0:0] f1240_clk;
  logic [0:0] f1240_rst;
  logic [31:0] f1240_rdata;
  sr_buffer_32_1 f1240(.wen(f1240_wen), .wdata(f1240_wdata), .clk(f1240_clk), .rst(f1240_rst), .rdata(f1240_rdata));
  assign f1240_clk = clk;
  assign f1240_rst = rst;
  // Bindings to f1240

  // f1242
  logic [0:0] f1242_wen;
  logic [31:0] f1242_wdata;
  logic [0:0] f1242_clk;
  logic [0:0] f1242_rst;
  logic [31:0] f1242_rdata;
  sr_buffer_32_1 f1242(.wen(f1242_wen), .wdata(f1242_wdata), .clk(f1242_clk), .rst(f1242_rst), .rdata(f1242_rdata));
  assign f1242_clk = clk;
  assign f1242_rst = rst;
  // Bindings to f1242

  // f1244
  logic [0:0] f1244_wen;
  logic [31:0] f1244_wdata;
  logic [0:0] f1244_clk;
  logic [0:0] f1244_rst;
  logic [31:0] f1244_rdata;
  sr_buffer_32_1 f1244(.wen(f1244_wen), .wdata(f1244_wdata), .clk(f1244_clk), .rst(f1244_rst), .rdata(f1244_rdata));
  assign f1244_clk = clk;
  assign f1244_rst = rst;
  // Bindings to f1244

  // f1246
  logic [0:0] f1246_wen;
  logic [31:0] f1246_wdata;
  logic [0:0] f1246_clk;
  logic [0:0] f1246_rst;
  logic [31:0] f1246_rdata;
  sr_buffer_32_1 f1246(.wen(f1246_wen), .wdata(f1246_wdata), .clk(f1246_clk), .rst(f1246_rst), .rdata(f1246_rdata));
  assign f1246_clk = clk;
  assign f1246_rst = rst;
  // Bindings to f1246

  // f1248
  logic [0:0] f1248_wen;
  logic [31:0] f1248_wdata;
  logic [0:0] f1248_clk;
  logic [0:0] f1248_rst;
  logic [31:0] f1248_rdata;
  sr_buffer_32_1 f1248(.wen(f1248_wen), .wdata(f1248_wdata), .clk(f1248_clk), .rst(f1248_rst), .rdata(f1248_rdata));
  assign f1248_clk = clk;
  assign f1248_rst = rst;
  // Bindings to f1248

  // f1250
  logic [0:0] f1250_wen;
  logic [31:0] f1250_wdata;
  logic [0:0] f1250_clk;
  logic [0:0] f1250_rst;
  logic [31:0] f1250_rdata;
  sr_buffer_32_1 f1250(.wen(f1250_wen), .wdata(f1250_wdata), .clk(f1250_clk), .rst(f1250_rst), .rdata(f1250_rdata));
  assign f1250_clk = clk;
  assign f1250_rst = rst;
  // Bindings to f1250

  // f1252
  logic [0:0] f1252_wen;
  logic [31:0] f1252_wdata;
  logic [0:0] f1252_clk;
  logic [0:0] f1252_rst;
  logic [31:0] f1252_rdata;
  sr_buffer_32_1 f1252(.wen(f1252_wen), .wdata(f1252_wdata), .clk(f1252_clk), .rst(f1252_rst), .rdata(f1252_rdata));
  assign f1252_clk = clk;
  assign f1252_rst = rst;
  // Bindings to f1252

  // f1254
  logic [0:0] f1254_wen;
  logic [31:0] f1254_wdata;
  logic [0:0] f1254_clk;
  logic [0:0] f1254_rst;
  logic [31:0] f1254_rdata;
  sr_buffer_32_1 f1254(.wen(f1254_wen), .wdata(f1254_wdata), .clk(f1254_clk), .rst(f1254_rst), .rdata(f1254_rdata));
  assign f1254_clk = clk;
  assign f1254_rst = rst;
  // Bindings to f1254

  // f1256
  logic [0:0] f1256_wen;
  logic [31:0] f1256_wdata;
  logic [0:0] f1256_clk;
  logic [0:0] f1256_rst;
  logic [31:0] f1256_rdata;
  sr_buffer_32_1 f1256(.wen(f1256_wen), .wdata(f1256_wdata), .clk(f1256_clk), .rst(f1256_rst), .rdata(f1256_rdata));
  assign f1256_clk = clk;
  assign f1256_rst = rst;
  // Bindings to f1256

  // f1258
  logic [0:0] f1258_wen;
  logic [31:0] f1258_wdata;
  logic [0:0] f1258_clk;
  logic [0:0] f1258_rst;
  logic [31:0] f1258_rdata;
  sr_buffer_32_1 f1258(.wen(f1258_wen), .wdata(f1258_wdata), .clk(f1258_clk), .rst(f1258_rst), .rdata(f1258_rdata));
  assign f1258_clk = clk;
  assign f1258_rst = rst;
  // Bindings to f1258

  // f1260
  logic [0:0] f1260_wen;
  logic [31:0] f1260_wdata;
  logic [0:0] f1260_clk;
  logic [0:0] f1260_rst;
  logic [31:0] f1260_rdata;
  sr_buffer_32_1 f1260(.wen(f1260_wen), .wdata(f1260_wdata), .clk(f1260_clk), .rst(f1260_rst), .rdata(f1260_rdata));
  assign f1260_clk = clk;
  assign f1260_rst = rst;
  // Bindings to f1260

  // f1262
  logic [0:0] f1262_wen;
  logic [31:0] f1262_wdata;
  logic [0:0] f1262_clk;
  logic [0:0] f1262_rst;
  logic [31:0] f1262_rdata;
  sr_buffer_32_1 f1262(.wen(f1262_wen), .wdata(f1262_wdata), .clk(f1262_clk), .rst(f1262_rst), .rdata(f1262_rdata));
  assign f1262_clk = clk;
  assign f1262_rst = rst;
  // Bindings to f1262

  // f1264
  logic [0:0] f1264_wen;
  logic [31:0] f1264_wdata;
  logic [0:0] f1264_clk;
  logic [0:0] f1264_rst;
  logic [31:0] f1264_rdata;
  sr_buffer_32_1 f1264(.wen(f1264_wen), .wdata(f1264_wdata), .clk(f1264_clk), .rst(f1264_rst), .rdata(f1264_rdata));
  assign f1264_clk = clk;
  assign f1264_rst = rst;
  // Bindings to f1264

  // f1266
  logic [0:0] f1266_wen;
  logic [31:0] f1266_wdata;
  logic [0:0] f1266_clk;
  logic [0:0] f1266_rst;
  logic [31:0] f1266_rdata;
  sr_buffer_32_1 f1266(.wen(f1266_wen), .wdata(f1266_wdata), .clk(f1266_clk), .rst(f1266_rst), .rdata(f1266_rdata));
  assign f1266_clk = clk;
  assign f1266_rst = rst;
  // Bindings to f1266

  // f1268
  logic [0:0] f1268_wen;
  logic [31:0] f1268_wdata;
  logic [0:0] f1268_clk;
  logic [0:0] f1268_rst;
  logic [31:0] f1268_rdata;
  sr_buffer_32_1 f1268(.wen(f1268_wen), .wdata(f1268_wdata), .clk(f1268_clk), .rst(f1268_rst), .rdata(f1268_rdata));
  assign f1268_clk = clk;
  assign f1268_rst = rst;
  // Bindings to f1268

  // f1270
  logic [0:0] f1270_wen;
  logic [31:0] f1270_wdata;
  logic [0:0] f1270_clk;
  logic [0:0] f1270_rst;
  logic [31:0] f1270_rdata;
  sr_buffer_32_1 f1270(.wen(f1270_wen), .wdata(f1270_wdata), .clk(f1270_clk), .rst(f1270_rst), .rdata(f1270_rdata));
  assign f1270_clk = clk;
  assign f1270_rst = rst;
  // Bindings to f1270

  // f1272
  logic [0:0] f1272_wen;
  logic [31:0] f1272_wdata;
  logic [0:0] f1272_clk;
  logic [0:0] f1272_rst;
  logic [31:0] f1272_rdata;
  sr_buffer_32_1 f1272(.wen(f1272_wen), .wdata(f1272_wdata), .clk(f1272_clk), .rst(f1272_rst), .rdata(f1272_rdata));
  assign f1272_clk = clk;
  assign f1272_rst = rst;
  // Bindings to f1272

  // f1274
  logic [0:0] f1274_wen;
  logic [31:0] f1274_wdata;
  logic [0:0] f1274_clk;
  logic [0:0] f1274_rst;
  logic [31:0] f1274_rdata;
  sr_buffer_32_1 f1274(.wen(f1274_wen), .wdata(f1274_wdata), .clk(f1274_clk), .rst(f1274_rst), .rdata(f1274_rdata));
  assign f1274_clk = clk;
  assign f1274_rst = rst;
  // Bindings to f1274

  // f1276
  logic [0:0] f1276_wen;
  logic [31:0] f1276_wdata;
  logic [0:0] f1276_clk;
  logic [0:0] f1276_rst;
  logic [31:0] f1276_rdata;
  sr_buffer_32_1 f1276(.wen(f1276_wen), .wdata(f1276_wdata), .clk(f1276_clk), .rst(f1276_rst), .rdata(f1276_rdata));
  assign f1276_clk = clk;
  assign f1276_rst = rst;
  // Bindings to f1276

  // f1278
  logic [0:0] f1278_wen;
  logic [31:0] f1278_wdata;
  logic [0:0] f1278_clk;
  logic [0:0] f1278_rst;
  logic [31:0] f1278_rdata;
  sr_buffer_32_1 f1278(.wen(f1278_wen), .wdata(f1278_wdata), .clk(f1278_clk), .rst(f1278_rst), .rdata(f1278_rdata));
  assign f1278_clk = clk;
  assign f1278_rst = rst;
  // Bindings to f1278

  // f1280
  logic [0:0] f1280_wen;
  logic [31:0] f1280_wdata;
  logic [0:0] f1280_clk;
  logic [0:0] f1280_rst;
  logic [31:0] f1280_rdata;
  sr_buffer_32_1 f1280(.wen(f1280_wen), .wdata(f1280_wdata), .clk(f1280_clk), .rst(f1280_rst), .rdata(f1280_rdata));
  assign f1280_clk = clk;
  assign f1280_rst = rst;
  // Bindings to f1280

  // f1282
  logic [0:0] f1282_wen;
  logic [31:0] f1282_wdata;
  logic [0:0] f1282_clk;
  logic [0:0] f1282_rst;
  logic [31:0] f1282_rdata;
  sr_buffer_32_1 f1282(.wen(f1282_wen), .wdata(f1282_wdata), .clk(f1282_clk), .rst(f1282_rst), .rdata(f1282_rdata));
  assign f1282_clk = clk;
  assign f1282_rst = rst;
  // Bindings to f1282

  // f1284
  logic [0:0] f1284_wen;
  logic [31:0] f1284_wdata;
  logic [0:0] f1284_clk;
  logic [0:0] f1284_rst;
  logic [31:0] f1284_rdata;
  sr_buffer_32_1 f1284(.wen(f1284_wen), .wdata(f1284_wdata), .clk(f1284_clk), .rst(f1284_rst), .rdata(f1284_rdata));
  assign f1284_clk = clk;
  assign f1284_rst = rst;
  // Bindings to f1284

  // f1286
  logic [0:0] f1286_wen;
  logic [31:0] f1286_wdata;
  logic [0:0] f1286_clk;
  logic [0:0] f1286_rst;
  logic [31:0] f1286_rdata;
  sr_buffer_32_1 f1286(.wen(f1286_wen), .wdata(f1286_wdata), .clk(f1286_clk), .rst(f1286_rst), .rdata(f1286_rdata));
  assign f1286_clk = clk;
  assign f1286_rst = rst;
  // Bindings to f1286

  // f1288
  logic [0:0] f1288_wen;
  logic [31:0] f1288_wdata;
  logic [0:0] f1288_clk;
  logic [0:0] f1288_rst;
  logic [31:0] f1288_rdata;
  sr_buffer_32_1 f1288(.wen(f1288_wen), .wdata(f1288_wdata), .clk(f1288_clk), .rst(f1288_rst), .rdata(f1288_rdata));
  assign f1288_clk = clk;
  assign f1288_rst = rst;
  // Bindings to f1288

  // f1290
  logic [0:0] f1290_wen;
  logic [31:0] f1290_wdata;
  logic [0:0] f1290_clk;
  logic [0:0] f1290_rst;
  logic [31:0] f1290_rdata;
  sr_buffer_32_1 f1290(.wen(f1290_wen), .wdata(f1290_wdata), .clk(f1290_clk), .rst(f1290_rst), .rdata(f1290_rdata));
  assign f1290_clk = clk;
  assign f1290_rst = rst;
  // Bindings to f1290

  // f1292
  logic [0:0] f1292_wen;
  logic [31:0] f1292_wdata;
  logic [0:0] f1292_clk;
  logic [0:0] f1292_rst;
  logic [31:0] f1292_rdata;
  sr_buffer_32_1 f1292(.wen(f1292_wen), .wdata(f1292_wdata), .clk(f1292_clk), .rst(f1292_rst), .rdata(f1292_rdata));
  assign f1292_clk = clk;
  assign f1292_rst = rst;
  // Bindings to f1292

  // f1294
  logic [0:0] f1294_wen;
  logic [31:0] f1294_wdata;
  logic [0:0] f1294_clk;
  logic [0:0] f1294_rst;
  logic [31:0] f1294_rdata;
  sr_buffer_32_1 f1294(.wen(f1294_wen), .wdata(f1294_wdata), .clk(f1294_clk), .rst(f1294_rst), .rdata(f1294_rdata));
  assign f1294_clk = clk;
  assign f1294_rst = rst;
  // Bindings to f1294

  // f1296
  logic [0:0] f1296_wen;
  logic [31:0] f1296_wdata;
  logic [0:0] f1296_clk;
  logic [0:0] f1296_rst;
  logic [31:0] f1296_rdata;
  sr_buffer_32_1 f1296(.wen(f1296_wen), .wdata(f1296_wdata), .clk(f1296_clk), .rst(f1296_rst), .rdata(f1296_rdata));
  assign f1296_clk = clk;
  assign f1296_rst = rst;
  // Bindings to f1296

  // f1298
  logic [0:0] f1298_wen;
  logic [31:0] f1298_wdata;
  logic [0:0] f1298_clk;
  logic [0:0] f1298_rst;
  logic [31:0] f1298_rdata;
  sr_buffer_32_1 f1298(.wen(f1298_wen), .wdata(f1298_wdata), .clk(f1298_clk), .rst(f1298_rst), .rdata(f1298_rdata));
  assign f1298_clk = clk;
  assign f1298_rst = rst;
  // Bindings to f1298

  // f1300
  logic [0:0] f1300_wen;
  logic [31:0] f1300_wdata;
  logic [0:0] f1300_clk;
  logic [0:0] f1300_rst;
  logic [31:0] f1300_rdata;
  sr_buffer_32_1 f1300(.wen(f1300_wen), .wdata(f1300_wdata), .clk(f1300_clk), .rst(f1300_rst), .rdata(f1300_rdata));
  assign f1300_clk = clk;
  assign f1300_rst = rst;
  // Bindings to f1300

  // f1302
  logic [0:0] f1302_wen;
  logic [31:0] f1302_wdata;
  logic [0:0] f1302_clk;
  logic [0:0] f1302_rst;
  logic [31:0] f1302_rdata;
  sr_buffer_32_1 f1302(.wen(f1302_wen), .wdata(f1302_wdata), .clk(f1302_clk), .rst(f1302_rst), .rdata(f1302_rdata));
  assign f1302_clk = clk;
  assign f1302_rst = rst;
  // Bindings to f1302

  // f1304
  logic [0:0] f1304_wen;
  logic [31:0] f1304_wdata;
  logic [0:0] f1304_clk;
  logic [0:0] f1304_rst;
  logic [31:0] f1304_rdata;
  sr_buffer_32_1 f1304(.wen(f1304_wen), .wdata(f1304_wdata), .clk(f1304_clk), .rst(f1304_rst), .rdata(f1304_rdata));
  assign f1304_clk = clk;
  assign f1304_rst = rst;
  // Bindings to f1304

  // f1306
  logic [0:0] f1306_wen;
  logic [31:0] f1306_wdata;
  logic [0:0] f1306_clk;
  logic [0:0] f1306_rst;
  logic [31:0] f1306_rdata;
  sr_buffer_32_1 f1306(.wen(f1306_wen), .wdata(f1306_wdata), .clk(f1306_clk), .rst(f1306_rst), .rdata(f1306_rdata));
  assign f1306_clk = clk;
  assign f1306_rst = rst;
  // Bindings to f1306

  // f1308
  logic [0:0] f1308_wen;
  logic [31:0] f1308_wdata;
  logic [0:0] f1308_clk;
  logic [0:0] f1308_rst;
  logic [31:0] f1308_rdata;
  sr_buffer_32_1 f1308(.wen(f1308_wen), .wdata(f1308_wdata), .clk(f1308_clk), .rst(f1308_rst), .rdata(f1308_rdata));
  assign f1308_clk = clk;
  assign f1308_rst = rst;
  // Bindings to f1308

  // f1310
  logic [0:0] f1310_wen;
  logic [31:0] f1310_wdata;
  logic [0:0] f1310_clk;
  logic [0:0] f1310_rst;
  logic [31:0] f1310_rdata;
  sr_buffer_32_1 f1310(.wen(f1310_wen), .wdata(f1310_wdata), .clk(f1310_clk), .rst(f1310_rst), .rdata(f1310_rdata));
  assign f1310_clk = clk;
  assign f1310_rst = rst;
  // Bindings to f1310

  // f1312
  logic [0:0] f1312_wen;
  logic [31:0] f1312_wdata;
  logic [0:0] f1312_clk;
  logic [0:0] f1312_rst;
  logic [31:0] f1312_rdata;
  sr_buffer_32_1 f1312(.wen(f1312_wen), .wdata(f1312_wdata), .clk(f1312_clk), .rst(f1312_rst), .rdata(f1312_rdata));
  assign f1312_clk = clk;
  assign f1312_rst = rst;
  // Bindings to f1312

  // f1314
  logic [0:0] f1314_wen;
  logic [31:0] f1314_wdata;
  logic [0:0] f1314_clk;
  logic [0:0] f1314_rst;
  logic [31:0] f1314_rdata;
  sr_buffer_32_1 f1314(.wen(f1314_wen), .wdata(f1314_wdata), .clk(f1314_clk), .rst(f1314_rst), .rdata(f1314_rdata));
  assign f1314_clk = clk;
  assign f1314_rst = rst;
  // Bindings to f1314

  // f1316
  logic [0:0] f1316_wen;
  logic [31:0] f1316_wdata;
  logic [0:0] f1316_clk;
  logic [0:0] f1316_rst;
  logic [31:0] f1316_rdata;
  sr_buffer_32_1 f1316(.wen(f1316_wen), .wdata(f1316_wdata), .clk(f1316_clk), .rst(f1316_rst), .rdata(f1316_rdata));
  assign f1316_clk = clk;
  assign f1316_rst = rst;
  // Bindings to f1316

  // f1318
  logic [0:0] f1318_wen;
  logic [31:0] f1318_wdata;
  logic [0:0] f1318_clk;
  logic [0:0] f1318_rst;
  logic [31:0] f1318_rdata;
  sr_buffer_32_1 f1318(.wen(f1318_wen), .wdata(f1318_wdata), .clk(f1318_clk), .rst(f1318_rst), .rdata(f1318_rdata));
  assign f1318_clk = clk;
  assign f1318_rst = rst;
  // Bindings to f1318

  // f1320
  logic [0:0] f1320_wen;
  logic [31:0] f1320_wdata;
  logic [0:0] f1320_clk;
  logic [0:0] f1320_rst;
  logic [31:0] f1320_rdata;
  sr_buffer_32_1 f1320(.wen(f1320_wen), .wdata(f1320_wdata), .clk(f1320_clk), .rst(f1320_rst), .rdata(f1320_rdata));
  assign f1320_clk = clk;
  assign f1320_rst = rst;
  // Bindings to f1320

  // f1322
  logic [0:0] f1322_wen;
  logic [31:0] f1322_wdata;
  logic [0:0] f1322_clk;
  logic [0:0] f1322_rst;
  logic [31:0] f1322_rdata;
  sr_buffer_32_1 f1322(.wen(f1322_wen), .wdata(f1322_wdata), .clk(f1322_clk), .rst(f1322_rst), .rdata(f1322_rdata));
  assign f1322_clk = clk;
  assign f1322_rst = rst;
  // Bindings to f1322

  // f1324
  logic [0:0] f1324_wen;
  logic [31:0] f1324_wdata;
  logic [0:0] f1324_clk;
  logic [0:0] f1324_rst;
  logic [31:0] f1324_rdata;
  sr_buffer_32_1 f1324(.wen(f1324_wen), .wdata(f1324_wdata), .clk(f1324_clk), .rst(f1324_rst), .rdata(f1324_rdata));
  assign f1324_clk = clk;
  assign f1324_rst = rst;
  // Bindings to f1324

  // f1326
  logic [0:0] f1326_wen;
  logic [31:0] f1326_wdata;
  logic [0:0] f1326_clk;
  logic [0:0] f1326_rst;
  logic [31:0] f1326_rdata;
  sr_buffer_32_1 f1326(.wen(f1326_wen), .wdata(f1326_wdata), .clk(f1326_clk), .rst(f1326_rst), .rdata(f1326_rdata));
  assign f1326_clk = clk;
  assign f1326_rst = rst;
  // Bindings to f1326

  // f1328
  logic [0:0] f1328_wen;
  logic [31:0] f1328_wdata;
  logic [0:0] f1328_clk;
  logic [0:0] f1328_rst;
  logic [31:0] f1328_rdata;
  sr_buffer_32_1 f1328(.wen(f1328_wen), .wdata(f1328_wdata), .clk(f1328_clk), .rst(f1328_rst), .rdata(f1328_rdata));
  assign f1328_clk = clk;
  assign f1328_rst = rst;
  // Bindings to f1328

  // f1330
  logic [0:0] f1330_wen;
  logic [31:0] f1330_wdata;
  logic [0:0] f1330_clk;
  logic [0:0] f1330_rst;
  logic [31:0] f1330_rdata;
  sr_buffer_32_1 f1330(.wen(f1330_wen), .wdata(f1330_wdata), .clk(f1330_clk), .rst(f1330_rst), .rdata(f1330_rdata));
  assign f1330_clk = clk;
  assign f1330_rst = rst;
  // Bindings to f1330

  // f1332
  logic [0:0] f1332_wen;
  logic [31:0] f1332_wdata;
  logic [0:0] f1332_clk;
  logic [0:0] f1332_rst;
  logic [31:0] f1332_rdata;
  sr_buffer_32_1 f1332(.wen(f1332_wen), .wdata(f1332_wdata), .clk(f1332_clk), .rst(f1332_rst), .rdata(f1332_rdata));
  assign f1332_clk = clk;
  assign f1332_rst = rst;
  // Bindings to f1332

  // f1334
  logic [0:0] f1334_wen;
  logic [31:0] f1334_wdata;
  logic [0:0] f1334_clk;
  logic [0:0] f1334_rst;
  logic [31:0] f1334_rdata;
  sr_buffer_32_1 f1334(.wen(f1334_wen), .wdata(f1334_wdata), .clk(f1334_clk), .rst(f1334_rst), .rdata(f1334_rdata));
  assign f1334_clk = clk;
  assign f1334_rst = rst;
  // Bindings to f1334

  // f1336
  logic [0:0] f1336_wen;
  logic [31:0] f1336_wdata;
  logic [0:0] f1336_clk;
  logic [0:0] f1336_rst;
  logic [31:0] f1336_rdata;
  sr_buffer_32_1 f1336(.wen(f1336_wen), .wdata(f1336_wdata), .clk(f1336_clk), .rst(f1336_rst), .rdata(f1336_rdata));
  assign f1336_clk = clk;
  assign f1336_rst = rst;
  // Bindings to f1336

  // f1338
  logic [0:0] f1338_wen;
  logic [31:0] f1338_wdata;
  logic [0:0] f1338_clk;
  logic [0:0] f1338_rst;
  logic [31:0] f1338_rdata;
  sr_buffer_32_1 f1338(.wen(f1338_wen), .wdata(f1338_wdata), .clk(f1338_clk), .rst(f1338_rst), .rdata(f1338_rdata));
  assign f1338_clk = clk;
  assign f1338_rst = rst;
  // Bindings to f1338

  // f1340
  logic [0:0] f1340_wen;
  logic [31:0] f1340_wdata;
  logic [0:0] f1340_clk;
  logic [0:0] f1340_rst;
  logic [31:0] f1340_rdata;
  sr_buffer_32_1 f1340(.wen(f1340_wen), .wdata(f1340_wdata), .clk(f1340_clk), .rst(f1340_rst), .rdata(f1340_rdata));
  assign f1340_clk = clk;
  assign f1340_rst = rst;
  // Bindings to f1340

  // f1342
  logic [0:0] f1342_wen;
  logic [31:0] f1342_wdata;
  logic [0:0] f1342_clk;
  logic [0:0] f1342_rst;
  logic [31:0] f1342_rdata;
  sr_buffer_32_1 f1342(.wen(f1342_wen), .wdata(f1342_wdata), .clk(f1342_clk), .rst(f1342_rst), .rdata(f1342_rdata));
  assign f1342_clk = clk;
  assign f1342_rst = rst;
  // Bindings to f1342

  // f1344
  logic [0:0] f1344_wen;
  logic [31:0] f1344_wdata;
  logic [0:0] f1344_clk;
  logic [0:0] f1344_rst;
  logic [31:0] f1344_rdata;
  sr_buffer_32_1 f1344(.wen(f1344_wen), .wdata(f1344_wdata), .clk(f1344_clk), .rst(f1344_rst), .rdata(f1344_rdata));
  assign f1344_clk = clk;
  assign f1344_rst = rst;
  // Bindings to f1344

  // f1346
  logic [0:0] f1346_wen;
  logic [31:0] f1346_wdata;
  logic [0:0] f1346_clk;
  logic [0:0] f1346_rst;
  logic [31:0] f1346_rdata;
  sr_buffer_32_1 f1346(.wen(f1346_wen), .wdata(f1346_wdata), .clk(f1346_clk), .rst(f1346_rst), .rdata(f1346_rdata));
  assign f1346_clk = clk;
  assign f1346_rst = rst;
  // Bindings to f1346

  // f1348
  logic [0:0] f1348_wen;
  logic [31:0] f1348_wdata;
  logic [0:0] f1348_clk;
  logic [0:0] f1348_rst;
  logic [31:0] f1348_rdata;
  sr_buffer_32_1 f1348(.wen(f1348_wen), .wdata(f1348_wdata), .clk(f1348_clk), .rst(f1348_rst), .rdata(f1348_rdata));
  assign f1348_clk = clk;
  assign f1348_rst = rst;
  // Bindings to f1348

  // f1350
  logic [0:0] f1350_wen;
  logic [31:0] f1350_wdata;
  logic [0:0] f1350_clk;
  logic [0:0] f1350_rst;
  logic [31:0] f1350_rdata;
  sr_buffer_32_1 f1350(.wen(f1350_wen), .wdata(f1350_wdata), .clk(f1350_clk), .rst(f1350_rst), .rdata(f1350_rdata));
  assign f1350_clk = clk;
  assign f1350_rst = rst;
  // Bindings to f1350

  // f1352
  logic [0:0] f1352_wen;
  logic [31:0] f1352_wdata;
  logic [0:0] f1352_clk;
  logic [0:0] f1352_rst;
  logic [31:0] f1352_rdata;
  sr_buffer_32_1 f1352(.wen(f1352_wen), .wdata(f1352_wdata), .clk(f1352_clk), .rst(f1352_rst), .rdata(f1352_rdata));
  assign f1352_clk = clk;
  assign f1352_rst = rst;
  // Bindings to f1352

  // f1354
  logic [0:0] f1354_wen;
  logic [31:0] f1354_wdata;
  logic [0:0] f1354_clk;
  logic [0:0] f1354_rst;
  logic [31:0] f1354_rdata;
  sr_buffer_32_1 f1354(.wen(f1354_wen), .wdata(f1354_wdata), .clk(f1354_clk), .rst(f1354_rst), .rdata(f1354_rdata));
  assign f1354_clk = clk;
  assign f1354_rst = rst;
  // Bindings to f1354

  // f1356
  logic [0:0] f1356_wen;
  logic [31:0] f1356_wdata;
  logic [0:0] f1356_clk;
  logic [0:0] f1356_rst;
  logic [31:0] f1356_rdata;
  sr_buffer_32_1 f1356(.wen(f1356_wen), .wdata(f1356_wdata), .clk(f1356_clk), .rst(f1356_rst), .rdata(f1356_rdata));
  assign f1356_clk = clk;
  assign f1356_rst = rst;
  // Bindings to f1356

  // f1358
  logic [0:0] f1358_wen;
  logic [31:0] f1358_wdata;
  logic [0:0] f1358_clk;
  logic [0:0] f1358_rst;
  logic [31:0] f1358_rdata;
  sr_buffer_32_1 f1358(.wen(f1358_wen), .wdata(f1358_wdata), .clk(f1358_clk), .rst(f1358_rst), .rdata(f1358_rdata));
  assign f1358_clk = clk;
  assign f1358_rst = rst;
  // Bindings to f1358

  // f1360
  logic [0:0] f1360_wen;
  logic [31:0] f1360_wdata;
  logic [0:0] f1360_clk;
  logic [0:0] f1360_rst;
  logic [31:0] f1360_rdata;
  sr_buffer_32_1 f1360(.wen(f1360_wen), .wdata(f1360_wdata), .clk(f1360_clk), .rst(f1360_rst), .rdata(f1360_rdata));
  assign f1360_clk = clk;
  assign f1360_rst = rst;
  // Bindings to f1360

  // f1362
  logic [0:0] f1362_wen;
  logic [31:0] f1362_wdata;
  logic [0:0] f1362_clk;
  logic [0:0] f1362_rst;
  logic [31:0] f1362_rdata;
  sr_buffer_32_1 f1362(.wen(f1362_wen), .wdata(f1362_wdata), .clk(f1362_clk), .rst(f1362_rst), .rdata(f1362_rdata));
  assign f1362_clk = clk;
  assign f1362_rst = rst;
  // Bindings to f1362

  // f1364
  logic [0:0] f1364_wen;
  logic [31:0] f1364_wdata;
  logic [0:0] f1364_clk;
  logic [0:0] f1364_rst;
  logic [31:0] f1364_rdata;
  sr_buffer_32_1 f1364(.wen(f1364_wen), .wdata(f1364_wdata), .clk(f1364_clk), .rst(f1364_rst), .rdata(f1364_rdata));
  assign f1364_clk = clk;
  assign f1364_rst = rst;
  // Bindings to f1364

  // f1366
  logic [0:0] f1366_wen;
  logic [31:0] f1366_wdata;
  logic [0:0] f1366_clk;
  logic [0:0] f1366_rst;
  logic [31:0] f1366_rdata;
  sr_buffer_32_1 f1366(.wen(f1366_wen), .wdata(f1366_wdata), .clk(f1366_clk), .rst(f1366_rst), .rdata(f1366_rdata));
  assign f1366_clk = clk;
  assign f1366_rst = rst;
  // Bindings to f1366

  // f1368
  logic [0:0] f1368_wen;
  logic [31:0] f1368_wdata;
  logic [0:0] f1368_clk;
  logic [0:0] f1368_rst;
  logic [31:0] f1368_rdata;
  sr_buffer_32_1 f1368(.wen(f1368_wen), .wdata(f1368_wdata), .clk(f1368_clk), .rst(f1368_rst), .rdata(f1368_rdata));
  assign f1368_clk = clk;
  assign f1368_rst = rst;
  // Bindings to f1368

  // f1370
  logic [0:0] f1370_wen;
  logic [31:0] f1370_wdata;
  logic [0:0] f1370_clk;
  logic [0:0] f1370_rst;
  logic [31:0] f1370_rdata;
  sr_buffer_32_1 f1370(.wen(f1370_wen), .wdata(f1370_wdata), .clk(f1370_clk), .rst(f1370_rst), .rdata(f1370_rdata));
  assign f1370_clk = clk;
  assign f1370_rst = rst;
  // Bindings to f1370

  // f1372
  logic [0:0] f1372_wen;
  logic [31:0] f1372_wdata;
  logic [0:0] f1372_clk;
  logic [0:0] f1372_rst;
  logic [31:0] f1372_rdata;
  sr_buffer_32_1 f1372(.wen(f1372_wen), .wdata(f1372_wdata), .clk(f1372_clk), .rst(f1372_rst), .rdata(f1372_rdata));
  assign f1372_clk = clk;
  assign f1372_rst = rst;
  // Bindings to f1372

  // f1374
  logic [0:0] f1374_wen;
  logic [31:0] f1374_wdata;
  logic [0:0] f1374_clk;
  logic [0:0] f1374_rst;
  logic [31:0] f1374_rdata;
  sr_buffer_32_1 f1374(.wen(f1374_wen), .wdata(f1374_wdata), .clk(f1374_clk), .rst(f1374_rst), .rdata(f1374_rdata));
  assign f1374_clk = clk;
  assign f1374_rst = rst;
  // Bindings to f1374

  // f1376
  logic [0:0] f1376_wen;
  logic [31:0] f1376_wdata;
  logic [0:0] f1376_clk;
  logic [0:0] f1376_rst;
  logic [31:0] f1376_rdata;
  sr_buffer_32_1 f1376(.wen(f1376_wen), .wdata(f1376_wdata), .clk(f1376_clk), .rst(f1376_rst), .rdata(f1376_rdata));
  assign f1376_clk = clk;
  assign f1376_rst = rst;
  // Bindings to f1376

  // f1378
  logic [0:0] f1378_wen;
  logic [31:0] f1378_wdata;
  logic [0:0] f1378_clk;
  logic [0:0] f1378_rst;
  logic [31:0] f1378_rdata;
  sr_buffer_32_1 f1378(.wen(f1378_wen), .wdata(f1378_wdata), .clk(f1378_clk), .rst(f1378_rst), .rdata(f1378_rdata));
  assign f1378_clk = clk;
  assign f1378_rst = rst;
  // Bindings to f1378

  // f1380
  logic [0:0] f1380_wen;
  logic [31:0] f1380_wdata;
  logic [0:0] f1380_clk;
  logic [0:0] f1380_rst;
  logic [31:0] f1380_rdata;
  sr_buffer_32_1 f1380(.wen(f1380_wen), .wdata(f1380_wdata), .clk(f1380_clk), .rst(f1380_rst), .rdata(f1380_rdata));
  assign f1380_clk = clk;
  assign f1380_rst = rst;
  // Bindings to f1380

  // f1382
  logic [0:0] f1382_wen;
  logic [31:0] f1382_wdata;
  logic [0:0] f1382_clk;
  logic [0:0] f1382_rst;
  logic [31:0] f1382_rdata;
  sr_buffer_32_1 f1382(.wen(f1382_wen), .wdata(f1382_wdata), .clk(f1382_clk), .rst(f1382_rst), .rdata(f1382_rdata));
  assign f1382_clk = clk;
  assign f1382_rst = rst;
  // Bindings to f1382

  // f1384
  logic [0:0] f1384_wen;
  logic [31:0] f1384_wdata;
  logic [0:0] f1384_clk;
  logic [0:0] f1384_rst;
  logic [31:0] f1384_rdata;
  sr_buffer_32_1 f1384(.wen(f1384_wen), .wdata(f1384_wdata), .clk(f1384_clk), .rst(f1384_rst), .rdata(f1384_rdata));
  assign f1384_clk = clk;
  assign f1384_rst = rst;
  // Bindings to f1384

  // f1386
  logic [0:0] f1386_wen;
  logic [31:0] f1386_wdata;
  logic [0:0] f1386_clk;
  logic [0:0] f1386_rst;
  logic [31:0] f1386_rdata;
  sr_buffer_32_1 f1386(.wen(f1386_wen), .wdata(f1386_wdata), .clk(f1386_clk), .rst(f1386_rst), .rdata(f1386_rdata));
  assign f1386_clk = clk;
  assign f1386_rst = rst;
  // Bindings to f1386

  // f1388
  logic [0:0] f1388_wen;
  logic [31:0] f1388_wdata;
  logic [0:0] f1388_clk;
  logic [0:0] f1388_rst;
  logic [31:0] f1388_rdata;
  sr_buffer_32_1 f1388(.wen(f1388_wen), .wdata(f1388_wdata), .clk(f1388_clk), .rst(f1388_rst), .rdata(f1388_rdata));
  assign f1388_clk = clk;
  assign f1388_rst = rst;
  // Bindings to f1388

  // f1390
  logic [0:0] f1390_wen;
  logic [31:0] f1390_wdata;
  logic [0:0] f1390_clk;
  logic [0:0] f1390_rst;
  logic [31:0] f1390_rdata;
  sr_buffer_32_1 f1390(.wen(f1390_wen), .wdata(f1390_wdata), .clk(f1390_clk), .rst(f1390_rst), .rdata(f1390_rdata));
  assign f1390_clk = clk;
  assign f1390_rst = rst;
  // Bindings to f1390

  // f1392
  logic [0:0] f1392_wen;
  logic [31:0] f1392_wdata;
  logic [0:0] f1392_clk;
  logic [0:0] f1392_rst;
  logic [31:0] f1392_rdata;
  sr_buffer_32_1 f1392(.wen(f1392_wen), .wdata(f1392_wdata), .clk(f1392_clk), .rst(f1392_rst), .rdata(f1392_rdata));
  assign f1392_clk = clk;
  assign f1392_rst = rst;
  // Bindings to f1392

  // f1394
  logic [0:0] f1394_wen;
  logic [31:0] f1394_wdata;
  logic [0:0] f1394_clk;
  logic [0:0] f1394_rst;
  logic [31:0] f1394_rdata;
  sr_buffer_32_1 f1394(.wen(f1394_wen), .wdata(f1394_wdata), .clk(f1394_clk), .rst(f1394_rst), .rdata(f1394_rdata));
  assign f1394_clk = clk;
  assign f1394_rst = rst;
  // Bindings to f1394

  // f1396
  logic [0:0] f1396_wen;
  logic [31:0] f1396_wdata;
  logic [0:0] f1396_clk;
  logic [0:0] f1396_rst;
  logic [31:0] f1396_rdata;
  sr_buffer_32_1 f1396(.wen(f1396_wen), .wdata(f1396_wdata), .clk(f1396_clk), .rst(f1396_rst), .rdata(f1396_rdata));
  assign f1396_clk = clk;
  assign f1396_rst = rst;
  // Bindings to f1396

  // f1398
  logic [0:0] f1398_wen;
  logic [31:0] f1398_wdata;
  logic [0:0] f1398_clk;
  logic [0:0] f1398_rst;
  logic [31:0] f1398_rdata;
  sr_buffer_32_1 f1398(.wen(f1398_wen), .wdata(f1398_wdata), .clk(f1398_clk), .rst(f1398_rst), .rdata(f1398_rdata));
  assign f1398_clk = clk;
  assign f1398_rst = rst;
  // Bindings to f1398

  // f1400
  logic [0:0] f1400_wen;
  logic [31:0] f1400_wdata;
  logic [0:0] f1400_clk;
  logic [0:0] f1400_rst;
  logic [31:0] f1400_rdata;
  sr_buffer_32_1 f1400(.wen(f1400_wen), .wdata(f1400_wdata), .clk(f1400_clk), .rst(f1400_rst), .rdata(f1400_rdata));
  assign f1400_clk = clk;
  assign f1400_rst = rst;
  // Bindings to f1400

  // f1402
  logic [0:0] f1402_wen;
  logic [31:0] f1402_wdata;
  logic [0:0] f1402_clk;
  logic [0:0] f1402_rst;
  logic [31:0] f1402_rdata;
  sr_buffer_32_1 f1402(.wen(f1402_wen), .wdata(f1402_wdata), .clk(f1402_clk), .rst(f1402_rst), .rdata(f1402_rdata));
  assign f1402_clk = clk;
  assign f1402_rst = rst;
  // Bindings to f1402

  // f1404
  logic [0:0] f1404_wen;
  logic [31:0] f1404_wdata;
  logic [0:0] f1404_clk;
  logic [0:0] f1404_rst;
  logic [31:0] f1404_rdata;
  sr_buffer_32_1 f1404(.wen(f1404_wen), .wdata(f1404_wdata), .clk(f1404_clk), .rst(f1404_rst), .rdata(f1404_rdata));
  assign f1404_clk = clk;
  assign f1404_rst = rst;
  // Bindings to f1404

  // f1406
  logic [0:0] f1406_wen;
  logic [31:0] f1406_wdata;
  logic [0:0] f1406_clk;
  logic [0:0] f1406_rst;
  logic [31:0] f1406_rdata;
  sr_buffer_32_1 f1406(.wen(f1406_wen), .wdata(f1406_wdata), .clk(f1406_clk), .rst(f1406_rst), .rdata(f1406_rdata));
  assign f1406_clk = clk;
  assign f1406_rst = rst;
  // Bindings to f1406

  // f1408
  logic [0:0] f1408_wen;
  logic [31:0] f1408_wdata;
  logic [0:0] f1408_clk;
  logic [0:0] f1408_rst;
  logic [31:0] f1408_rdata;
  sr_buffer_32_1 f1408(.wen(f1408_wen), .wdata(f1408_wdata), .clk(f1408_clk), .rst(f1408_rst), .rdata(f1408_rdata));
  assign f1408_clk = clk;
  assign f1408_rst = rst;
  // Bindings to f1408

  // f1410
  logic [0:0] f1410_wen;
  logic [31:0] f1410_wdata;
  logic [0:0] f1410_clk;
  logic [0:0] f1410_rst;
  logic [31:0] f1410_rdata;
  sr_buffer_32_1 f1410(.wen(f1410_wen), .wdata(f1410_wdata), .clk(f1410_clk), .rst(f1410_rst), .rdata(f1410_rdata));
  assign f1410_clk = clk;
  assign f1410_rst = rst;
  // Bindings to f1410

  // f1412
  logic [0:0] f1412_wen;
  logic [31:0] f1412_wdata;
  logic [0:0] f1412_clk;
  logic [0:0] f1412_rst;
  logic [31:0] f1412_rdata;
  sr_buffer_32_1 f1412(.wen(f1412_wen), .wdata(f1412_wdata), .clk(f1412_clk), .rst(f1412_rst), .rdata(f1412_rdata));
  assign f1412_clk = clk;
  assign f1412_rst = rst;
  // Bindings to f1412

  // f1414
  logic [0:0] f1414_wen;
  logic [31:0] f1414_wdata;
  logic [0:0] f1414_clk;
  logic [0:0] f1414_rst;
  logic [31:0] f1414_rdata;
  sr_buffer_32_1 f1414(.wen(f1414_wen), .wdata(f1414_wdata), .clk(f1414_clk), .rst(f1414_rst), .rdata(f1414_rdata));
  assign f1414_clk = clk;
  assign f1414_rst = rst;
  // Bindings to f1414

  // f1416
  logic [0:0] f1416_wen;
  logic [31:0] f1416_wdata;
  logic [0:0] f1416_clk;
  logic [0:0] f1416_rst;
  logic [31:0] f1416_rdata;
  sr_buffer_32_1 f1416(.wen(f1416_wen), .wdata(f1416_wdata), .clk(f1416_clk), .rst(f1416_rst), .rdata(f1416_rdata));
  assign f1416_clk = clk;
  assign f1416_rst = rst;
  // Bindings to f1416

  // f1418
  logic [0:0] f1418_wen;
  logic [31:0] f1418_wdata;
  logic [0:0] f1418_clk;
  logic [0:0] f1418_rst;
  logic [31:0] f1418_rdata;
  sr_buffer_32_1 f1418(.wen(f1418_wen), .wdata(f1418_wdata), .clk(f1418_clk), .rst(f1418_rst), .rdata(f1418_rdata));
  assign f1418_clk = clk;
  assign f1418_rst = rst;
  // Bindings to f1418

  // f1420
  logic [0:0] f1420_wen;
  logic [31:0] f1420_wdata;
  logic [0:0] f1420_clk;
  logic [0:0] f1420_rst;
  logic [31:0] f1420_rdata;
  sr_buffer_32_1 f1420(.wen(f1420_wen), .wdata(f1420_wdata), .clk(f1420_clk), .rst(f1420_rst), .rdata(f1420_rdata));
  assign f1420_clk = clk;
  assign f1420_rst = rst;
  // Bindings to f1420

  // f1422
  logic [0:0] f1422_wen;
  logic [31:0] f1422_wdata;
  logic [0:0] f1422_clk;
  logic [0:0] f1422_rst;
  logic [31:0] f1422_rdata;
  sr_buffer_32_1 f1422(.wen(f1422_wen), .wdata(f1422_wdata), .clk(f1422_clk), .rst(f1422_rst), .rdata(f1422_rdata));
  assign f1422_clk = clk;
  assign f1422_rst = rst;
  // Bindings to f1422

  // f1424
  logic [0:0] f1424_wen;
  logic [31:0] f1424_wdata;
  logic [0:0] f1424_clk;
  logic [0:0] f1424_rst;
  logic [31:0] f1424_rdata;
  sr_buffer_32_1 f1424(.wen(f1424_wen), .wdata(f1424_wdata), .clk(f1424_clk), .rst(f1424_rst), .rdata(f1424_rdata));
  assign f1424_clk = clk;
  assign f1424_rst = rst;
  // Bindings to f1424

  // f1426
  logic [0:0] f1426_wen;
  logic [31:0] f1426_wdata;
  logic [0:0] f1426_clk;
  logic [0:0] f1426_rst;
  logic [31:0] f1426_rdata;
  sr_buffer_32_1 f1426(.wen(f1426_wen), .wdata(f1426_wdata), .clk(f1426_clk), .rst(f1426_rst), .rdata(f1426_rdata));
  assign f1426_clk = clk;
  assign f1426_rst = rst;
  // Bindings to f1426

  // f1428
  logic [0:0] f1428_wen;
  logic [31:0] f1428_wdata;
  logic [0:0] f1428_clk;
  logic [0:0] f1428_rst;
  logic [31:0] f1428_rdata;
  sr_buffer_32_1 f1428(.wen(f1428_wen), .wdata(f1428_wdata), .clk(f1428_clk), .rst(f1428_rst), .rdata(f1428_rdata));
  assign f1428_clk = clk;
  assign f1428_rst = rst;
  // Bindings to f1428

  // f1430
  logic [0:0] f1430_wen;
  logic [31:0] f1430_wdata;
  logic [0:0] f1430_clk;
  logic [0:0] f1430_rst;
  logic [31:0] f1430_rdata;
  sr_buffer_32_1 f1430(.wen(f1430_wen), .wdata(f1430_wdata), .clk(f1430_clk), .rst(f1430_rst), .rdata(f1430_rdata));
  assign f1430_clk = clk;
  assign f1430_rst = rst;
  // Bindings to f1430

  // f1432
  logic [0:0] f1432_wen;
  logic [31:0] f1432_wdata;
  logic [0:0] f1432_clk;
  logic [0:0] f1432_rst;
  logic [31:0] f1432_rdata;
  sr_buffer_32_1 f1432(.wen(f1432_wen), .wdata(f1432_wdata), .clk(f1432_clk), .rst(f1432_rst), .rdata(f1432_rdata));
  assign f1432_clk = clk;
  assign f1432_rst = rst;
  // Bindings to f1432

  // f1434
  logic [0:0] f1434_wen;
  logic [31:0] f1434_wdata;
  logic [0:0] f1434_clk;
  logic [0:0] f1434_rst;
  logic [31:0] f1434_rdata;
  sr_buffer_32_1 f1434(.wen(f1434_wen), .wdata(f1434_wdata), .clk(f1434_clk), .rst(f1434_rst), .rdata(f1434_rdata));
  assign f1434_clk = clk;
  assign f1434_rst = rst;
  // Bindings to f1434

  // f1436
  logic [0:0] f1436_wen;
  logic [31:0] f1436_wdata;
  logic [0:0] f1436_clk;
  logic [0:0] f1436_rst;
  logic [31:0] f1436_rdata;
  sr_buffer_32_1 f1436(.wen(f1436_wen), .wdata(f1436_wdata), .clk(f1436_clk), .rst(f1436_rst), .rdata(f1436_rdata));
  assign f1436_clk = clk;
  assign f1436_rst = rst;
  // Bindings to f1436

  // f1438
  logic [0:0] f1438_wen;
  logic [31:0] f1438_wdata;
  logic [0:0] f1438_clk;
  logic [0:0] f1438_rst;
  logic [31:0] f1438_rdata;
  sr_buffer_32_1 f1438(.wen(f1438_wen), .wdata(f1438_wdata), .clk(f1438_clk), .rst(f1438_rst), .rdata(f1438_rdata));
  assign f1438_clk = clk;
  assign f1438_rst = rst;
  // Bindings to f1438

  // f1440
  logic [0:0] f1440_wen;
  logic [31:0] f1440_wdata;
  logic [0:0] f1440_clk;
  logic [0:0] f1440_rst;
  logic [31:0] f1440_rdata;
  sr_buffer_32_1 f1440(.wen(f1440_wen), .wdata(f1440_wdata), .clk(f1440_clk), .rst(f1440_rst), .rdata(f1440_rdata));
  assign f1440_clk = clk;
  assign f1440_rst = rst;
  // Bindings to f1440

  // f1442
  logic [0:0] f1442_wen;
  logic [31:0] f1442_wdata;
  logic [0:0] f1442_clk;
  logic [0:0] f1442_rst;
  logic [31:0] f1442_rdata;
  sr_buffer_32_1 f1442(.wen(f1442_wen), .wdata(f1442_wdata), .clk(f1442_clk), .rst(f1442_rst), .rdata(f1442_rdata));
  assign f1442_clk = clk;
  assign f1442_rst = rst;
  // Bindings to f1442

  // f1444
  logic [0:0] f1444_wen;
  logic [31:0] f1444_wdata;
  logic [0:0] f1444_clk;
  logic [0:0] f1444_rst;
  logic [31:0] f1444_rdata;
  sr_buffer_32_1 f1444(.wen(f1444_wen), .wdata(f1444_wdata), .clk(f1444_clk), .rst(f1444_rst), .rdata(f1444_rdata));
  assign f1444_clk = clk;
  assign f1444_rst = rst;
  // Bindings to f1444

  // f1446
  logic [0:0] f1446_wen;
  logic [31:0] f1446_wdata;
  logic [0:0] f1446_clk;
  logic [0:0] f1446_rst;
  logic [31:0] f1446_rdata;
  sr_buffer_32_1 f1446(.wen(f1446_wen), .wdata(f1446_wdata), .clk(f1446_clk), .rst(f1446_rst), .rdata(f1446_rdata));
  assign f1446_clk = clk;
  assign f1446_rst = rst;
  // Bindings to f1446

  // f1448
  logic [0:0] f1448_wen;
  logic [31:0] f1448_wdata;
  logic [0:0] f1448_clk;
  logic [0:0] f1448_rst;
  logic [31:0] f1448_rdata;
  sr_buffer_32_1 f1448(.wen(f1448_wen), .wdata(f1448_wdata), .clk(f1448_clk), .rst(f1448_rst), .rdata(f1448_rdata));
  assign f1448_clk = clk;
  assign f1448_rst = rst;
  // Bindings to f1448

  // f1450
  logic [0:0] f1450_wen;
  logic [31:0] f1450_wdata;
  logic [0:0] f1450_clk;
  logic [0:0] f1450_rst;
  logic [31:0] f1450_rdata;
  sr_buffer_32_1 f1450(.wen(f1450_wen), .wdata(f1450_wdata), .clk(f1450_clk), .rst(f1450_rst), .rdata(f1450_rdata));
  assign f1450_clk = clk;
  assign f1450_rst = rst;
  // Bindings to f1450

  // f1452
  logic [0:0] f1452_wen;
  logic [31:0] f1452_wdata;
  logic [0:0] f1452_clk;
  logic [0:0] f1452_rst;
  logic [31:0] f1452_rdata;
  sr_buffer_32_1 f1452(.wen(f1452_wen), .wdata(f1452_wdata), .clk(f1452_clk), .rst(f1452_rst), .rdata(f1452_rdata));
  assign f1452_clk = clk;
  assign f1452_rst = rst;
  // Bindings to f1452

  // f1454
  logic [0:0] f1454_wen;
  logic [31:0] f1454_wdata;
  logic [0:0] f1454_clk;
  logic [0:0] f1454_rst;
  logic [31:0] f1454_rdata;
  sr_buffer_32_1 f1454(.wen(f1454_wen), .wdata(f1454_wdata), .clk(f1454_clk), .rst(f1454_rst), .rdata(f1454_rdata));
  assign f1454_clk = clk;
  assign f1454_rst = rst;
  // Bindings to f1454

  // f1456
  logic [0:0] f1456_wen;
  logic [31:0] f1456_wdata;
  logic [0:0] f1456_clk;
  logic [0:0] f1456_rst;
  logic [31:0] f1456_rdata;
  sr_buffer_32_1 f1456(.wen(f1456_wen), .wdata(f1456_wdata), .clk(f1456_clk), .rst(f1456_rst), .rdata(f1456_rdata));
  assign f1456_clk = clk;
  assign f1456_rst = rst;
  // Bindings to f1456

  // f1458
  logic [0:0] f1458_wen;
  logic [31:0] f1458_wdata;
  logic [0:0] f1458_clk;
  logic [0:0] f1458_rst;
  logic [31:0] f1458_rdata;
  sr_buffer_32_1 f1458(.wen(f1458_wen), .wdata(f1458_wdata), .clk(f1458_clk), .rst(f1458_rst), .rdata(f1458_rdata));
  assign f1458_clk = clk;
  assign f1458_rst = rst;
  // Bindings to f1458

  // f1460
  logic [0:0] f1460_wen;
  logic [31:0] f1460_wdata;
  logic [0:0] f1460_clk;
  logic [0:0] f1460_rst;
  logic [31:0] f1460_rdata;
  sr_buffer_32_1 f1460(.wen(f1460_wen), .wdata(f1460_wdata), .clk(f1460_clk), .rst(f1460_rst), .rdata(f1460_rdata));
  assign f1460_clk = clk;
  assign f1460_rst = rst;
  // Bindings to f1460

  // f1462
  logic [0:0] f1462_wen;
  logic [31:0] f1462_wdata;
  logic [0:0] f1462_clk;
  logic [0:0] f1462_rst;
  logic [31:0] f1462_rdata;
  sr_buffer_32_1 f1462(.wen(f1462_wen), .wdata(f1462_wdata), .clk(f1462_clk), .rst(f1462_rst), .rdata(f1462_rdata));
  assign f1462_clk = clk;
  assign f1462_rst = rst;
  // Bindings to f1462

  // f1464
  logic [0:0] f1464_wen;
  logic [31:0] f1464_wdata;
  logic [0:0] f1464_clk;
  logic [0:0] f1464_rst;
  logic [31:0] f1464_rdata;
  sr_buffer_32_1 f1464(.wen(f1464_wen), .wdata(f1464_wdata), .clk(f1464_clk), .rst(f1464_rst), .rdata(f1464_rdata));
  assign f1464_clk = clk;
  assign f1464_rst = rst;
  // Bindings to f1464

  // f1466
  logic [0:0] f1466_wen;
  logic [31:0] f1466_wdata;
  logic [0:0] f1466_clk;
  logic [0:0] f1466_rst;
  logic [31:0] f1466_rdata;
  sr_buffer_32_1 f1466(.wen(f1466_wen), .wdata(f1466_wdata), .clk(f1466_clk), .rst(f1466_rst), .rdata(f1466_rdata));
  assign f1466_clk = clk;
  assign f1466_rst = rst;
  // Bindings to f1466

  // f1468
  logic [0:0] f1468_wen;
  logic [31:0] f1468_wdata;
  logic [0:0] f1468_clk;
  logic [0:0] f1468_rst;
  logic [31:0] f1468_rdata;
  sr_buffer_32_1 f1468(.wen(f1468_wen), .wdata(f1468_wdata), .clk(f1468_clk), .rst(f1468_rst), .rdata(f1468_rdata));
  assign f1468_clk = clk;
  assign f1468_rst = rst;
  // Bindings to f1468

  // f1470
  logic [0:0] f1470_wen;
  logic [31:0] f1470_wdata;
  logic [0:0] f1470_clk;
  logic [0:0] f1470_rst;
  logic [31:0] f1470_rdata;
  sr_buffer_32_1 f1470(.wen(f1470_wen), .wdata(f1470_wdata), .clk(f1470_clk), .rst(f1470_rst), .rdata(f1470_rdata));
  assign f1470_clk = clk;
  assign f1470_rst = rst;
  // Bindings to f1470

  // f1472
  logic [0:0] f1472_wen;
  logic [31:0] f1472_wdata;
  logic [0:0] f1472_clk;
  logic [0:0] f1472_rst;
  logic [31:0] f1472_rdata;
  sr_buffer_32_1 f1472(.wen(f1472_wen), .wdata(f1472_wdata), .clk(f1472_clk), .rst(f1472_rst), .rdata(f1472_rdata));
  assign f1472_clk = clk;
  assign f1472_rst = rst;
  // Bindings to f1472

  // f1474
  logic [0:0] f1474_wen;
  logic [31:0] f1474_wdata;
  logic [0:0] f1474_clk;
  logic [0:0] f1474_rst;
  logic [31:0] f1474_rdata;
  sr_buffer_32_1 f1474(.wen(f1474_wen), .wdata(f1474_wdata), .clk(f1474_clk), .rst(f1474_rst), .rdata(f1474_rdata));
  assign f1474_clk = clk;
  assign f1474_rst = rst;
  // Bindings to f1474

  // f1476
  logic [0:0] f1476_wen;
  logic [31:0] f1476_wdata;
  logic [0:0] f1476_clk;
  logic [0:0] f1476_rst;
  logic [31:0] f1476_rdata;
  sr_buffer_32_1 f1476(.wen(f1476_wen), .wdata(f1476_wdata), .clk(f1476_clk), .rst(f1476_rst), .rdata(f1476_rdata));
  assign f1476_clk = clk;
  assign f1476_rst = rst;
  // Bindings to f1476

  // f1478
  logic [0:0] f1478_wen;
  logic [31:0] f1478_wdata;
  logic [0:0] f1478_clk;
  logic [0:0] f1478_rst;
  logic [31:0] f1478_rdata;
  sr_buffer_32_1 f1478(.wen(f1478_wen), .wdata(f1478_wdata), .clk(f1478_clk), .rst(f1478_rst), .rdata(f1478_rdata));
  assign f1478_clk = clk;
  assign f1478_rst = rst;
  // Bindings to f1478

  // f1480
  logic [0:0] f1480_wen;
  logic [31:0] f1480_wdata;
  logic [0:0] f1480_clk;
  logic [0:0] f1480_rst;
  logic [31:0] f1480_rdata;
  sr_buffer_32_1 f1480(.wen(f1480_wen), .wdata(f1480_wdata), .clk(f1480_clk), .rst(f1480_rst), .rdata(f1480_rdata));
  assign f1480_clk = clk;
  assign f1480_rst = rst;
  // Bindings to f1480

  // f1482
  logic [0:0] f1482_wen;
  logic [31:0] f1482_wdata;
  logic [0:0] f1482_clk;
  logic [0:0] f1482_rst;
  logic [31:0] f1482_rdata;
  sr_buffer_32_1 f1482(.wen(f1482_wen), .wdata(f1482_wdata), .clk(f1482_clk), .rst(f1482_rst), .rdata(f1482_rdata));
  assign f1482_clk = clk;
  assign f1482_rst = rst;
  // Bindings to f1482

  // f1484
  logic [0:0] f1484_wen;
  logic [31:0] f1484_wdata;
  logic [0:0] f1484_clk;
  logic [0:0] f1484_rst;
  logic [31:0] f1484_rdata;
  sr_buffer_32_1 f1484(.wen(f1484_wen), .wdata(f1484_wdata), .clk(f1484_clk), .rst(f1484_rst), .rdata(f1484_rdata));
  assign f1484_clk = clk;
  assign f1484_rst = rst;
  // Bindings to f1484

  // f1486
  logic [0:0] f1486_wen;
  logic [31:0] f1486_wdata;
  logic [0:0] f1486_clk;
  logic [0:0] f1486_rst;
  logic [31:0] f1486_rdata;
  sr_buffer_32_1 f1486(.wen(f1486_wen), .wdata(f1486_wdata), .clk(f1486_clk), .rst(f1486_rst), .rdata(f1486_rdata));
  assign f1486_clk = clk;
  assign f1486_rst = rst;
  // Bindings to f1486

  // f1488
  logic [0:0] f1488_wen;
  logic [31:0] f1488_wdata;
  logic [0:0] f1488_clk;
  logic [0:0] f1488_rst;
  logic [31:0] f1488_rdata;
  sr_buffer_32_1 f1488(.wen(f1488_wen), .wdata(f1488_wdata), .clk(f1488_clk), .rst(f1488_rst), .rdata(f1488_rdata));
  assign f1488_clk = clk;
  assign f1488_rst = rst;
  // Bindings to f1488

  // f1490
  logic [0:0] f1490_wen;
  logic [31:0] f1490_wdata;
  logic [0:0] f1490_clk;
  logic [0:0] f1490_rst;
  logic [31:0] f1490_rdata;
  sr_buffer_32_1 f1490(.wen(f1490_wen), .wdata(f1490_wdata), .clk(f1490_clk), .rst(f1490_rst), .rdata(f1490_rdata));
  assign f1490_clk = clk;
  assign f1490_rst = rst;
  // Bindings to f1490

  // f1492
  logic [0:0] f1492_wen;
  logic [31:0] f1492_wdata;
  logic [0:0] f1492_clk;
  logic [0:0] f1492_rst;
  logic [31:0] f1492_rdata;
  sr_buffer_32_1 f1492(.wen(f1492_wen), .wdata(f1492_wdata), .clk(f1492_clk), .rst(f1492_rst), .rdata(f1492_rdata));
  assign f1492_clk = clk;
  assign f1492_rst = rst;
  // Bindings to f1492

  // f1494
  logic [0:0] f1494_wen;
  logic [31:0] f1494_wdata;
  logic [0:0] f1494_clk;
  logic [0:0] f1494_rst;
  logic [31:0] f1494_rdata;
  sr_buffer_32_1 f1494(.wen(f1494_wen), .wdata(f1494_wdata), .clk(f1494_clk), .rst(f1494_rst), .rdata(f1494_rdata));
  assign f1494_clk = clk;
  assign f1494_rst = rst;
  // Bindings to f1494

  // f1496
  logic [0:0] f1496_wen;
  logic [31:0] f1496_wdata;
  logic [0:0] f1496_clk;
  logic [0:0] f1496_rst;
  logic [31:0] f1496_rdata;
  sr_buffer_32_1 f1496(.wen(f1496_wen), .wdata(f1496_wdata), .clk(f1496_clk), .rst(f1496_rst), .rdata(f1496_rdata));
  assign f1496_clk = clk;
  assign f1496_rst = rst;
  // Bindings to f1496

  // f1498
  logic [0:0] f1498_wen;
  logic [31:0] f1498_wdata;
  logic [0:0] f1498_clk;
  logic [0:0] f1498_rst;
  logic [31:0] f1498_rdata;
  sr_buffer_32_1 f1498(.wen(f1498_wen), .wdata(f1498_wdata), .clk(f1498_clk), .rst(f1498_rst), .rdata(f1498_rdata));
  assign f1498_clk = clk;
  assign f1498_rst = rst;
  // Bindings to f1498

  // f1500
  logic [0:0] f1500_wen;
  logic [31:0] f1500_wdata;
  logic [0:0] f1500_clk;
  logic [0:0] f1500_rst;
  logic [31:0] f1500_rdata;
  sr_buffer_32_1 f1500(.wen(f1500_wen), .wdata(f1500_wdata), .clk(f1500_clk), .rst(f1500_rst), .rdata(f1500_rdata));
  assign f1500_clk = clk;
  assign f1500_rst = rst;
  // Bindings to f1500

  // f1502
  logic [0:0] f1502_wen;
  logic [31:0] f1502_wdata;
  logic [0:0] f1502_clk;
  logic [0:0] f1502_rst;
  logic [31:0] f1502_rdata;
  sr_buffer_32_1 f1502(.wen(f1502_wen), .wdata(f1502_wdata), .clk(f1502_clk), .rst(f1502_rst), .rdata(f1502_rdata));
  assign f1502_clk = clk;
  assign f1502_rst = rst;
  // Bindings to f1502

  // f1504
  logic [0:0] f1504_wen;
  logic [31:0] f1504_wdata;
  logic [0:0] f1504_clk;
  logic [0:0] f1504_rst;
  logic [31:0] f1504_rdata;
  sr_buffer_32_1 f1504(.wen(f1504_wen), .wdata(f1504_wdata), .clk(f1504_clk), .rst(f1504_rst), .rdata(f1504_rdata));
  assign f1504_clk = clk;
  assign f1504_rst = rst;
  // Bindings to f1504

  // f1506
  logic [0:0] f1506_wen;
  logic [31:0] f1506_wdata;
  logic [0:0] f1506_clk;
  logic [0:0] f1506_rst;
  logic [31:0] f1506_rdata;
  sr_buffer_32_1 f1506(.wen(f1506_wen), .wdata(f1506_wdata), .clk(f1506_clk), .rst(f1506_rst), .rdata(f1506_rdata));
  assign f1506_clk = clk;
  assign f1506_rst = rst;
  // Bindings to f1506

  // f1508
  logic [0:0] f1508_wen;
  logic [31:0] f1508_wdata;
  logic [0:0] f1508_clk;
  logic [0:0] f1508_rst;
  logic [31:0] f1508_rdata;
  sr_buffer_32_1 f1508(.wen(f1508_wen), .wdata(f1508_wdata), .clk(f1508_clk), .rst(f1508_rst), .rdata(f1508_rdata));
  assign f1508_clk = clk;
  assign f1508_rst = rst;
  // Bindings to f1508

  // f1510
  logic [0:0] f1510_wen;
  logic [31:0] f1510_wdata;
  logic [0:0] f1510_clk;
  logic [0:0] f1510_rst;
  logic [31:0] f1510_rdata;
  sr_buffer_32_1 f1510(.wen(f1510_wen), .wdata(f1510_wdata), .clk(f1510_clk), .rst(f1510_rst), .rdata(f1510_rdata));
  assign f1510_clk = clk;
  assign f1510_rst = rst;
  // Bindings to f1510

  // f1512
  logic [0:0] f1512_wen;
  logic [31:0] f1512_wdata;
  logic [0:0] f1512_clk;
  logic [0:0] f1512_rst;
  logic [31:0] f1512_rdata;
  sr_buffer_32_1 f1512(.wen(f1512_wen), .wdata(f1512_wdata), .clk(f1512_clk), .rst(f1512_rst), .rdata(f1512_rdata));
  assign f1512_clk = clk;
  assign f1512_rst = rst;
  // Bindings to f1512

  // f1514
  logic [0:0] f1514_wen;
  logic [31:0] f1514_wdata;
  logic [0:0] f1514_clk;
  logic [0:0] f1514_rst;
  logic [31:0] f1514_rdata;
  sr_buffer_32_1 f1514(.wen(f1514_wen), .wdata(f1514_wdata), .clk(f1514_clk), .rst(f1514_rst), .rdata(f1514_rdata));
  assign f1514_clk = clk;
  assign f1514_rst = rst;
  // Bindings to f1514

  // f1516
  logic [0:0] f1516_wen;
  logic [31:0] f1516_wdata;
  logic [0:0] f1516_clk;
  logic [0:0] f1516_rst;
  logic [31:0] f1516_rdata;
  sr_buffer_32_1 f1516(.wen(f1516_wen), .wdata(f1516_wdata), .clk(f1516_clk), .rst(f1516_rst), .rdata(f1516_rdata));
  assign f1516_clk = clk;
  assign f1516_rst = rst;
  // Bindings to f1516

  // f1518
  logic [0:0] f1518_wen;
  logic [31:0] f1518_wdata;
  logic [0:0] f1518_clk;
  logic [0:0] f1518_rst;
  logic [31:0] f1518_rdata;
  sr_buffer_32_1 f1518(.wen(f1518_wen), .wdata(f1518_wdata), .clk(f1518_clk), .rst(f1518_rst), .rdata(f1518_rdata));
  assign f1518_clk = clk;
  assign f1518_rst = rst;
  // Bindings to f1518

  // f1520
  logic [0:0] f1520_wen;
  logic [31:0] f1520_wdata;
  logic [0:0] f1520_clk;
  logic [0:0] f1520_rst;
  logic [31:0] f1520_rdata;
  sr_buffer_32_1 f1520(.wen(f1520_wen), .wdata(f1520_wdata), .clk(f1520_clk), .rst(f1520_rst), .rdata(f1520_rdata));
  assign f1520_clk = clk;
  assign f1520_rst = rst;
  // Bindings to f1520

  // f1522
  logic [0:0] f1522_wen;
  logic [31:0] f1522_wdata;
  logic [0:0] f1522_clk;
  logic [0:0] f1522_rst;
  logic [31:0] f1522_rdata;
  sr_buffer_32_1 f1522(.wen(f1522_wen), .wdata(f1522_wdata), .clk(f1522_clk), .rst(f1522_rst), .rdata(f1522_rdata));
  assign f1522_clk = clk;
  assign f1522_rst = rst;
  // Bindings to f1522

  // f1524
  logic [0:0] f1524_wen;
  logic [31:0] f1524_wdata;
  logic [0:0] f1524_clk;
  logic [0:0] f1524_rst;
  logic [31:0] f1524_rdata;
  sr_buffer_32_1 f1524(.wen(f1524_wen), .wdata(f1524_wdata), .clk(f1524_clk), .rst(f1524_rst), .rdata(f1524_rdata));
  assign f1524_clk = clk;
  assign f1524_rst = rst;
  // Bindings to f1524

  // f1526
  logic [0:0] f1526_wen;
  logic [31:0] f1526_wdata;
  logic [0:0] f1526_clk;
  logic [0:0] f1526_rst;
  logic [31:0] f1526_rdata;
  sr_buffer_32_1 f1526(.wen(f1526_wen), .wdata(f1526_wdata), .clk(f1526_clk), .rst(f1526_rst), .rdata(f1526_rdata));
  assign f1526_clk = clk;
  assign f1526_rst = rst;
  // Bindings to f1526

  // f1528
  logic [0:0] f1528_wen;
  logic [31:0] f1528_wdata;
  logic [0:0] f1528_clk;
  logic [0:0] f1528_rst;
  logic [31:0] f1528_rdata;
  sr_buffer_32_1 f1528(.wen(f1528_wen), .wdata(f1528_wdata), .clk(f1528_clk), .rst(f1528_rst), .rdata(f1528_rdata));
  assign f1528_clk = clk;
  assign f1528_rst = rst;
  // Bindings to f1528

  // f1530
  logic [0:0] f1530_wen;
  logic [31:0] f1530_wdata;
  logic [0:0] f1530_clk;
  logic [0:0] f1530_rst;
  logic [31:0] f1530_rdata;
  sr_buffer_32_1 f1530(.wen(f1530_wen), .wdata(f1530_wdata), .clk(f1530_clk), .rst(f1530_rst), .rdata(f1530_rdata));
  assign f1530_clk = clk;
  assign f1530_rst = rst;
  // Bindings to f1530

  // f1532
  logic [0:0] f1532_wen;
  logic [31:0] f1532_wdata;
  logic [0:0] f1532_clk;
  logic [0:0] f1532_rst;
  logic [31:0] f1532_rdata;
  sr_buffer_32_1 f1532(.wen(f1532_wen), .wdata(f1532_wdata), .clk(f1532_clk), .rst(f1532_rst), .rdata(f1532_rdata));
  assign f1532_clk = clk;
  assign f1532_rst = rst;
  // Bindings to f1532

  // f1534
  logic [0:0] f1534_wen;
  logic [31:0] f1534_wdata;
  logic [0:0] f1534_clk;
  logic [0:0] f1534_rst;
  logic [31:0] f1534_rdata;
  sr_buffer_32_1 f1534(.wen(f1534_wen), .wdata(f1534_wdata), .clk(f1534_clk), .rst(f1534_rst), .rdata(f1534_rdata));
  assign f1534_clk = clk;
  assign f1534_rst = rst;
  // Bindings to f1534

  // f1536
  logic [0:0] f1536_wen;
  logic [31:0] f1536_wdata;
  logic [0:0] f1536_clk;
  logic [0:0] f1536_rst;
  logic [31:0] f1536_rdata;
  sr_buffer_32_1 f1536(.wen(f1536_wen), .wdata(f1536_wdata), .clk(f1536_clk), .rst(f1536_rst), .rdata(f1536_rdata));
  assign f1536_clk = clk;
  assign f1536_rst = rst;
  // Bindings to f1536

  // f1538
  logic [0:0] f1538_wen;
  logic [31:0] f1538_wdata;
  logic [0:0] f1538_clk;
  logic [0:0] f1538_rst;
  logic [31:0] f1538_rdata;
  sr_buffer_32_1 f1538(.wen(f1538_wen), .wdata(f1538_wdata), .clk(f1538_clk), .rst(f1538_rst), .rdata(f1538_rdata));
  assign f1538_clk = clk;
  assign f1538_rst = rst;
  // Bindings to f1538

  // f1540
  logic [0:0] f1540_wen;
  logic [31:0] f1540_wdata;
  logic [0:0] f1540_clk;
  logic [0:0] f1540_rst;
  logic [31:0] f1540_rdata;
  sr_buffer_32_1 f1540(.wen(f1540_wen), .wdata(f1540_wdata), .clk(f1540_clk), .rst(f1540_rst), .rdata(f1540_rdata));
  assign f1540_clk = clk;
  assign f1540_rst = rst;
  // Bindings to f1540

  // f1542
  logic [0:0] f1542_wen;
  logic [31:0] f1542_wdata;
  logic [0:0] f1542_clk;
  logic [0:0] f1542_rst;
  logic [31:0] f1542_rdata;
  sr_buffer_32_1 f1542(.wen(f1542_wen), .wdata(f1542_wdata), .clk(f1542_clk), .rst(f1542_rst), .rdata(f1542_rdata));
  assign f1542_clk = clk;
  assign f1542_rst = rst;
  // Bindings to f1542

  // f1544
  logic [0:0] f1544_wen;
  logic [31:0] f1544_wdata;
  logic [0:0] f1544_clk;
  logic [0:0] f1544_rst;
  logic [31:0] f1544_rdata;
  sr_buffer_32_1 f1544(.wen(f1544_wen), .wdata(f1544_wdata), .clk(f1544_clk), .rst(f1544_rst), .rdata(f1544_rdata));
  assign f1544_clk = clk;
  assign f1544_rst = rst;
  // Bindings to f1544

  // f1546
  logic [0:0] f1546_wen;
  logic [31:0] f1546_wdata;
  logic [0:0] f1546_clk;
  logic [0:0] f1546_rst;
  logic [31:0] f1546_rdata;
  sr_buffer_32_1 f1546(.wen(f1546_wen), .wdata(f1546_wdata), .clk(f1546_clk), .rst(f1546_rst), .rdata(f1546_rdata));
  assign f1546_clk = clk;
  assign f1546_rst = rst;
  // Bindings to f1546

  // f1548
  logic [0:0] f1548_wen;
  logic [31:0] f1548_wdata;
  logic [0:0] f1548_clk;
  logic [0:0] f1548_rst;
  logic [31:0] f1548_rdata;
  sr_buffer_32_1 f1548(.wen(f1548_wen), .wdata(f1548_wdata), .clk(f1548_clk), .rst(f1548_rst), .rdata(f1548_rdata));
  assign f1548_clk = clk;
  assign f1548_rst = rst;
  // Bindings to f1548

  // f1550
  logic [0:0] f1550_wen;
  logic [31:0] f1550_wdata;
  logic [0:0] f1550_clk;
  logic [0:0] f1550_rst;
  logic [31:0] f1550_rdata;
  sr_buffer_32_1 f1550(.wen(f1550_wen), .wdata(f1550_wdata), .clk(f1550_clk), .rst(f1550_rst), .rdata(f1550_rdata));
  assign f1550_clk = clk;
  assign f1550_rst = rst;
  // Bindings to f1550

  // f1552
  logic [0:0] f1552_wen;
  logic [31:0] f1552_wdata;
  logic [0:0] f1552_clk;
  logic [0:0] f1552_rst;
  logic [31:0] f1552_rdata;
  sr_buffer_32_1 f1552(.wen(f1552_wen), .wdata(f1552_wdata), .clk(f1552_clk), .rst(f1552_rst), .rdata(f1552_rdata));
  assign f1552_clk = clk;
  assign f1552_rst = rst;
  // Bindings to f1552

  // f1554
  logic [0:0] f1554_wen;
  logic [31:0] f1554_wdata;
  logic [0:0] f1554_clk;
  logic [0:0] f1554_rst;
  logic [31:0] f1554_rdata;
  sr_buffer_32_1 f1554(.wen(f1554_wen), .wdata(f1554_wdata), .clk(f1554_clk), .rst(f1554_rst), .rdata(f1554_rdata));
  assign f1554_clk = clk;
  assign f1554_rst = rst;
  // Bindings to f1554

  // f1556
  logic [0:0] f1556_wen;
  logic [31:0] f1556_wdata;
  logic [0:0] f1556_clk;
  logic [0:0] f1556_rst;
  logic [31:0] f1556_rdata;
  sr_buffer_32_1 f1556(.wen(f1556_wen), .wdata(f1556_wdata), .clk(f1556_clk), .rst(f1556_rst), .rdata(f1556_rdata));
  assign f1556_clk = clk;
  assign f1556_rst = rst;
  // Bindings to f1556

  // f1558
  logic [0:0] f1558_wen;
  logic [31:0] f1558_wdata;
  logic [0:0] f1558_clk;
  logic [0:0] f1558_rst;
  logic [31:0] f1558_rdata;
  sr_buffer_32_1 f1558(.wen(f1558_wen), .wdata(f1558_wdata), .clk(f1558_clk), .rst(f1558_rst), .rdata(f1558_rdata));
  assign f1558_clk = clk;
  assign f1558_rst = rst;
  // Bindings to f1558

  // f1560
  logic [0:0] f1560_wen;
  logic [31:0] f1560_wdata;
  logic [0:0] f1560_clk;
  logic [0:0] f1560_rst;
  logic [31:0] f1560_rdata;
  sr_buffer_32_1 f1560(.wen(f1560_wen), .wdata(f1560_wdata), .clk(f1560_clk), .rst(f1560_rst), .rdata(f1560_rdata));
  assign f1560_clk = clk;
  assign f1560_rst = rst;
  // Bindings to f1560

  // f1562
  logic [0:0] f1562_wen;
  logic [31:0] f1562_wdata;
  logic [0:0] f1562_clk;
  logic [0:0] f1562_rst;
  logic [31:0] f1562_rdata;
  sr_buffer_32_1 f1562(.wen(f1562_wen), .wdata(f1562_wdata), .clk(f1562_clk), .rst(f1562_rst), .rdata(f1562_rdata));
  assign f1562_clk = clk;
  assign f1562_rst = rst;
  // Bindings to f1562

  // f1564
  logic [0:0] f1564_wen;
  logic [31:0] f1564_wdata;
  logic [0:0] f1564_clk;
  logic [0:0] f1564_rst;
  logic [31:0] f1564_rdata;
  sr_buffer_32_1 f1564(.wen(f1564_wen), .wdata(f1564_wdata), .clk(f1564_clk), .rst(f1564_rst), .rdata(f1564_rdata));
  assign f1564_clk = clk;
  assign f1564_rst = rst;
  // Bindings to f1564

  // f1566
  logic [0:0] f1566_wen;
  logic [31:0] f1566_wdata;
  logic [0:0] f1566_clk;
  logic [0:0] f1566_rst;
  logic [31:0] f1566_rdata;
  sr_buffer_32_1 f1566(.wen(f1566_wen), .wdata(f1566_wdata), .clk(f1566_clk), .rst(f1566_rst), .rdata(f1566_rdata));
  assign f1566_clk = clk;
  assign f1566_rst = rst;
  // Bindings to f1566

  // f1568
  logic [0:0] f1568_wen;
  logic [31:0] f1568_wdata;
  logic [0:0] f1568_clk;
  logic [0:0] f1568_rst;
  logic [31:0] f1568_rdata;
  sr_buffer_32_1 f1568(.wen(f1568_wen), .wdata(f1568_wdata), .clk(f1568_clk), .rst(f1568_rst), .rdata(f1568_rdata));
  assign f1568_clk = clk;
  assign f1568_rst = rst;
  // Bindings to f1568

  // f1570
  logic [0:0] f1570_wen;
  logic [31:0] f1570_wdata;
  logic [0:0] f1570_clk;
  logic [0:0] f1570_rst;
  logic [31:0] f1570_rdata;
  sr_buffer_32_1 f1570(.wen(f1570_wen), .wdata(f1570_wdata), .clk(f1570_clk), .rst(f1570_rst), .rdata(f1570_rdata));
  assign f1570_clk = clk;
  assign f1570_rst = rst;
  // Bindings to f1570

  // f1572
  logic [0:0] f1572_wen;
  logic [31:0] f1572_wdata;
  logic [0:0] f1572_clk;
  logic [0:0] f1572_rst;
  logic [31:0] f1572_rdata;
  sr_buffer_32_1 f1572(.wen(f1572_wen), .wdata(f1572_wdata), .clk(f1572_clk), .rst(f1572_rst), .rdata(f1572_rdata));
  assign f1572_clk = clk;
  assign f1572_rst = rst;
  // Bindings to f1572

  // f1574
  logic [0:0] f1574_wen;
  logic [31:0] f1574_wdata;
  logic [0:0] f1574_clk;
  logic [0:0] f1574_rst;
  logic [31:0] f1574_rdata;
  sr_buffer_32_1 f1574(.wen(f1574_wen), .wdata(f1574_wdata), .clk(f1574_clk), .rst(f1574_rst), .rdata(f1574_rdata));
  assign f1574_clk = clk;
  assign f1574_rst = rst;
  // Bindings to f1574

  // f1576
  logic [0:0] f1576_wen;
  logic [31:0] f1576_wdata;
  logic [0:0] f1576_clk;
  logic [0:0] f1576_rst;
  logic [31:0] f1576_rdata;
  sr_buffer_32_1 f1576(.wen(f1576_wen), .wdata(f1576_wdata), .clk(f1576_clk), .rst(f1576_rst), .rdata(f1576_rdata));
  assign f1576_clk = clk;
  assign f1576_rst = rst;
  // Bindings to f1576

  // f1578
  logic [0:0] f1578_wen;
  logic [31:0] f1578_wdata;
  logic [0:0] f1578_clk;
  logic [0:0] f1578_rst;
  logic [31:0] f1578_rdata;
  sr_buffer_32_1 f1578(.wen(f1578_wen), .wdata(f1578_wdata), .clk(f1578_clk), .rst(f1578_rst), .rdata(f1578_rdata));
  assign f1578_clk = clk;
  assign f1578_rst = rst;
  // Bindings to f1578

  // f1580
  logic [0:0] f1580_wen;
  logic [31:0] f1580_wdata;
  logic [0:0] f1580_clk;
  logic [0:0] f1580_rst;
  logic [31:0] f1580_rdata;
  sr_buffer_32_1 f1580(.wen(f1580_wen), .wdata(f1580_wdata), .clk(f1580_clk), .rst(f1580_rst), .rdata(f1580_rdata));
  assign f1580_clk = clk;
  assign f1580_rst = rst;
  // Bindings to f1580

  // f1582
  logic [0:0] f1582_wen;
  logic [31:0] f1582_wdata;
  logic [0:0] f1582_clk;
  logic [0:0] f1582_rst;
  logic [31:0] f1582_rdata;
  sr_buffer_32_1 f1582(.wen(f1582_wen), .wdata(f1582_wdata), .clk(f1582_clk), .rst(f1582_rst), .rdata(f1582_rdata));
  assign f1582_clk = clk;
  assign f1582_rst = rst;
  // Bindings to f1582

  // f1584
  logic [0:0] f1584_wen;
  logic [31:0] f1584_wdata;
  logic [0:0] f1584_clk;
  logic [0:0] f1584_rst;
  logic [31:0] f1584_rdata;
  sr_buffer_32_1 f1584(.wen(f1584_wen), .wdata(f1584_wdata), .clk(f1584_clk), .rst(f1584_rst), .rdata(f1584_rdata));
  assign f1584_clk = clk;
  assign f1584_rst = rst;
  // Bindings to f1584

  // f1586
  logic [0:0] f1586_wen;
  logic [31:0] f1586_wdata;
  logic [0:0] f1586_clk;
  logic [0:0] f1586_rst;
  logic [31:0] f1586_rdata;
  sr_buffer_32_1 f1586(.wen(f1586_wen), .wdata(f1586_wdata), .clk(f1586_clk), .rst(f1586_rst), .rdata(f1586_rdata));
  assign f1586_clk = clk;
  assign f1586_rst = rst;
  // Bindings to f1586

  // f1588
  logic [0:0] f1588_wen;
  logic [31:0] f1588_wdata;
  logic [0:0] f1588_clk;
  logic [0:0] f1588_rst;
  logic [31:0] f1588_rdata;
  sr_buffer_32_1 f1588(.wen(f1588_wen), .wdata(f1588_wdata), .clk(f1588_clk), .rst(f1588_rst), .rdata(f1588_rdata));
  assign f1588_clk = clk;
  assign f1588_rst = rst;
  // Bindings to f1588

  // f1590
  logic [0:0] f1590_wen;
  logic [31:0] f1590_wdata;
  logic [0:0] f1590_clk;
  logic [0:0] f1590_rst;
  logic [31:0] f1590_rdata;
  sr_buffer_32_1 f1590(.wen(f1590_wen), .wdata(f1590_wdata), .clk(f1590_clk), .rst(f1590_rst), .rdata(f1590_rdata));
  assign f1590_clk = clk;
  assign f1590_rst = rst;
  // Bindings to f1590

  // f1592
  logic [0:0] f1592_wen;
  logic [31:0] f1592_wdata;
  logic [0:0] f1592_clk;
  logic [0:0] f1592_rst;
  logic [31:0] f1592_rdata;
  sr_buffer_32_1 f1592(.wen(f1592_wen), .wdata(f1592_wdata), .clk(f1592_clk), .rst(f1592_rst), .rdata(f1592_rdata));
  assign f1592_clk = clk;
  assign f1592_rst = rst;
  // Bindings to f1592

  // f1594
  logic [0:0] f1594_wen;
  logic [31:0] f1594_wdata;
  logic [0:0] f1594_clk;
  logic [0:0] f1594_rst;
  logic [31:0] f1594_rdata;
  sr_buffer_32_1 f1594(.wen(f1594_wen), .wdata(f1594_wdata), .clk(f1594_clk), .rst(f1594_rst), .rdata(f1594_rdata));
  assign f1594_clk = clk;
  assign f1594_rst = rst;
  // Bindings to f1594

  // f1596
  logic [0:0] f1596_wen;
  logic [31:0] f1596_wdata;
  logic [0:0] f1596_clk;
  logic [0:0] f1596_rst;
  logic [31:0] f1596_rdata;
  sr_buffer_32_1 f1596(.wen(f1596_wen), .wdata(f1596_wdata), .clk(f1596_clk), .rst(f1596_rst), .rdata(f1596_rdata));
  assign f1596_clk = clk;
  assign f1596_rst = rst;
  // Bindings to f1596

  // f1598
  logic [0:0] f1598_wen;
  logic [31:0] f1598_wdata;
  logic [0:0] f1598_clk;
  logic [0:0] f1598_rst;
  logic [31:0] f1598_rdata;
  sr_buffer_32_1 f1598(.wen(f1598_wen), .wdata(f1598_wdata), .clk(f1598_clk), .rst(f1598_rst), .rdata(f1598_rdata));
  assign f1598_clk = clk;
  assign f1598_rst = rst;
  // Bindings to f1598

  // f1600
  logic [0:0] f1600_wen;
  logic [31:0] f1600_wdata;
  logic [0:0] f1600_clk;
  logic [0:0] f1600_rst;
  logic [31:0] f1600_rdata;
  sr_buffer_32_1 f1600(.wen(f1600_wen), .wdata(f1600_wdata), .clk(f1600_clk), .rst(f1600_rst), .rdata(f1600_rdata));
  assign f1600_clk = clk;
  assign f1600_rst = rst;
  // Bindings to f1600

  // f1602
  logic [0:0] f1602_wen;
  logic [31:0] f1602_wdata;
  logic [0:0] f1602_clk;
  logic [0:0] f1602_rst;
  logic [31:0] f1602_rdata;
  sr_buffer_32_1 f1602(.wen(f1602_wen), .wdata(f1602_wdata), .clk(f1602_clk), .rst(f1602_rst), .rdata(f1602_rdata));
  assign f1602_clk = clk;
  assign f1602_rst = rst;
  // Bindings to f1602

  // f1604
  logic [0:0] f1604_wen;
  logic [31:0] f1604_wdata;
  logic [0:0] f1604_clk;
  logic [0:0] f1604_rst;
  logic [31:0] f1604_rdata;
  sr_buffer_32_1 f1604(.wen(f1604_wen), .wdata(f1604_wdata), .clk(f1604_clk), .rst(f1604_rst), .rdata(f1604_rdata));
  assign f1604_clk = clk;
  assign f1604_rst = rst;
  // Bindings to f1604

  // f1606
  logic [0:0] f1606_wen;
  logic [31:0] f1606_wdata;
  logic [0:0] f1606_clk;
  logic [0:0] f1606_rst;
  logic [31:0] f1606_rdata;
  sr_buffer_32_1 f1606(.wen(f1606_wen), .wdata(f1606_wdata), .clk(f1606_clk), .rst(f1606_rst), .rdata(f1606_rdata));
  assign f1606_clk = clk;
  assign f1606_rst = rst;
  // Bindings to f1606

  // f1608
  logic [0:0] f1608_wen;
  logic [31:0] f1608_wdata;
  logic [0:0] f1608_clk;
  logic [0:0] f1608_rst;
  logic [31:0] f1608_rdata;
  sr_buffer_32_1 f1608(.wen(f1608_wen), .wdata(f1608_wdata), .clk(f1608_clk), .rst(f1608_rst), .rdata(f1608_rdata));
  assign f1608_clk = clk;
  assign f1608_rst = rst;
  // Bindings to f1608

  // f1610
  logic [0:0] f1610_wen;
  logic [31:0] f1610_wdata;
  logic [0:0] f1610_clk;
  logic [0:0] f1610_rst;
  logic [31:0] f1610_rdata;
  sr_buffer_32_1 f1610(.wen(f1610_wen), .wdata(f1610_wdata), .clk(f1610_clk), .rst(f1610_rst), .rdata(f1610_rdata));
  assign f1610_clk = clk;
  assign f1610_rst = rst;
  // Bindings to f1610

  // f1612
  logic [0:0] f1612_wen;
  logic [31:0] f1612_wdata;
  logic [0:0] f1612_clk;
  logic [0:0] f1612_rst;
  logic [31:0] f1612_rdata;
  sr_buffer_32_1 f1612(.wen(f1612_wen), .wdata(f1612_wdata), .clk(f1612_clk), .rst(f1612_rst), .rdata(f1612_rdata));
  assign f1612_clk = clk;
  assign f1612_rst = rst;
  // Bindings to f1612

  // f1614
  logic [0:0] f1614_wen;
  logic [31:0] f1614_wdata;
  logic [0:0] f1614_clk;
  logic [0:0] f1614_rst;
  logic [31:0] f1614_rdata;
  sr_buffer_32_1 f1614(.wen(f1614_wen), .wdata(f1614_wdata), .clk(f1614_clk), .rst(f1614_rst), .rdata(f1614_rdata));
  assign f1614_clk = clk;
  assign f1614_rst = rst;
  // Bindings to f1614

  // f1616
  logic [0:0] f1616_wen;
  logic [31:0] f1616_wdata;
  logic [0:0] f1616_clk;
  logic [0:0] f1616_rst;
  logic [31:0] f1616_rdata;
  sr_buffer_32_1 f1616(.wen(f1616_wen), .wdata(f1616_wdata), .clk(f1616_clk), .rst(f1616_rst), .rdata(f1616_rdata));
  assign f1616_clk = clk;
  assign f1616_rst = rst;
  // Bindings to f1616

  // f1618
  logic [0:0] f1618_wen;
  logic [31:0] f1618_wdata;
  logic [0:0] f1618_clk;
  logic [0:0] f1618_rst;
  logic [31:0] f1618_rdata;
  sr_buffer_32_1 f1618(.wen(f1618_wen), .wdata(f1618_wdata), .clk(f1618_clk), .rst(f1618_rst), .rdata(f1618_rdata));
  assign f1618_clk = clk;
  assign f1618_rst = rst;
  // Bindings to f1618

  // f1620
  logic [0:0] f1620_wen;
  logic [31:0] f1620_wdata;
  logic [0:0] f1620_clk;
  logic [0:0] f1620_rst;
  logic [31:0] f1620_rdata;
  sr_buffer_32_1 f1620(.wen(f1620_wen), .wdata(f1620_wdata), .clk(f1620_clk), .rst(f1620_rst), .rdata(f1620_rdata));
  assign f1620_clk = clk;
  assign f1620_rst = rst;
  // Bindings to f1620

  // f1622
  logic [0:0] f1622_wen;
  logic [31:0] f1622_wdata;
  logic [0:0] f1622_clk;
  logic [0:0] f1622_rst;
  logic [31:0] f1622_rdata;
  sr_buffer_32_1 f1622(.wen(f1622_wen), .wdata(f1622_wdata), .clk(f1622_clk), .rst(f1622_rst), .rdata(f1622_rdata));
  assign f1622_clk = clk;
  assign f1622_rst = rst;
  // Bindings to f1622

  // f1624
  logic [0:0] f1624_wen;
  logic [31:0] f1624_wdata;
  logic [0:0] f1624_clk;
  logic [0:0] f1624_rst;
  logic [31:0] f1624_rdata;
  sr_buffer_32_1 f1624(.wen(f1624_wen), .wdata(f1624_wdata), .clk(f1624_clk), .rst(f1624_rst), .rdata(f1624_rdata));
  assign f1624_clk = clk;
  assign f1624_rst = rst;
  // Bindings to f1624

  // f1626
  logic [0:0] f1626_wen;
  logic [31:0] f1626_wdata;
  logic [0:0] f1626_clk;
  logic [0:0] f1626_rst;
  logic [31:0] f1626_rdata;
  sr_buffer_32_1 f1626(.wen(f1626_wen), .wdata(f1626_wdata), .clk(f1626_clk), .rst(f1626_rst), .rdata(f1626_rdata));
  assign f1626_clk = clk;
  assign f1626_rst = rst;
  // Bindings to f1626

  // f1628
  logic [0:0] f1628_wen;
  logic [31:0] f1628_wdata;
  logic [0:0] f1628_clk;
  logic [0:0] f1628_rst;
  logic [31:0] f1628_rdata;
  sr_buffer_32_1 f1628(.wen(f1628_wen), .wdata(f1628_wdata), .clk(f1628_clk), .rst(f1628_rst), .rdata(f1628_rdata));
  assign f1628_clk = clk;
  assign f1628_rst = rst;
  // Bindings to f1628

  // f1630
  logic [0:0] f1630_wen;
  logic [31:0] f1630_wdata;
  logic [0:0] f1630_clk;
  logic [0:0] f1630_rst;
  logic [31:0] f1630_rdata;
  sr_buffer_32_1 f1630(.wen(f1630_wen), .wdata(f1630_wdata), .clk(f1630_clk), .rst(f1630_rst), .rdata(f1630_rdata));
  assign f1630_clk = clk;
  assign f1630_rst = rst;
  // Bindings to f1630

  // f1632
  logic [0:0] f1632_wen;
  logic [31:0] f1632_wdata;
  logic [0:0] f1632_clk;
  logic [0:0] f1632_rst;
  logic [31:0] f1632_rdata;
  sr_buffer_32_1 f1632(.wen(f1632_wen), .wdata(f1632_wdata), .clk(f1632_clk), .rst(f1632_rst), .rdata(f1632_rdata));
  assign f1632_clk = clk;
  assign f1632_rst = rst;
  // Bindings to f1632

  // f1634
  logic [0:0] f1634_wen;
  logic [31:0] f1634_wdata;
  logic [0:0] f1634_clk;
  logic [0:0] f1634_rst;
  logic [31:0] f1634_rdata;
  sr_buffer_32_1 f1634(.wen(f1634_wen), .wdata(f1634_wdata), .clk(f1634_clk), .rst(f1634_rst), .rdata(f1634_rdata));
  assign f1634_clk = clk;
  assign f1634_rst = rst;
  // Bindings to f1634

  // f1636
  logic [0:0] f1636_wen;
  logic [31:0] f1636_wdata;
  logic [0:0] f1636_clk;
  logic [0:0] f1636_rst;
  logic [31:0] f1636_rdata;
  sr_buffer_32_1 f1636(.wen(f1636_wen), .wdata(f1636_wdata), .clk(f1636_clk), .rst(f1636_rst), .rdata(f1636_rdata));
  assign f1636_clk = clk;
  assign f1636_rst = rst;
  // Bindings to f1636

  // f1638
  logic [0:0] f1638_wen;
  logic [31:0] f1638_wdata;
  logic [0:0] f1638_clk;
  logic [0:0] f1638_rst;
  logic [31:0] f1638_rdata;
  sr_buffer_32_1 f1638(.wen(f1638_wen), .wdata(f1638_wdata), .clk(f1638_clk), .rst(f1638_rst), .rdata(f1638_rdata));
  assign f1638_clk = clk;
  assign f1638_rst = rst;
  // Bindings to f1638

  // f1640
  logic [0:0] f1640_wen;
  logic [31:0] f1640_wdata;
  logic [0:0] f1640_clk;
  logic [0:0] f1640_rst;
  logic [31:0] f1640_rdata;
  sr_buffer_32_1 f1640(.wen(f1640_wen), .wdata(f1640_wdata), .clk(f1640_clk), .rst(f1640_rst), .rdata(f1640_rdata));
  assign f1640_clk = clk;
  assign f1640_rst = rst;
  // Bindings to f1640

  // f1642
  logic [0:0] f1642_wen;
  logic [31:0] f1642_wdata;
  logic [0:0] f1642_clk;
  logic [0:0] f1642_rst;
  logic [31:0] f1642_rdata;
  sr_buffer_32_1 f1642(.wen(f1642_wen), .wdata(f1642_wdata), .clk(f1642_clk), .rst(f1642_rst), .rdata(f1642_rdata));
  assign f1642_clk = clk;
  assign f1642_rst = rst;
  // Bindings to f1642

  // f1644
  logic [0:0] f1644_wen;
  logic [31:0] f1644_wdata;
  logic [0:0] f1644_clk;
  logic [0:0] f1644_rst;
  logic [31:0] f1644_rdata;
  sr_buffer_32_1 f1644(.wen(f1644_wen), .wdata(f1644_wdata), .clk(f1644_clk), .rst(f1644_rst), .rdata(f1644_rdata));
  assign f1644_clk = clk;
  assign f1644_rst = rst;
  // Bindings to f1644

  // f1646
  logic [0:0] f1646_wen;
  logic [31:0] f1646_wdata;
  logic [0:0] f1646_clk;
  logic [0:0] f1646_rst;
  logic [31:0] f1646_rdata;
  sr_buffer_32_1 f1646(.wen(f1646_wen), .wdata(f1646_wdata), .clk(f1646_clk), .rst(f1646_rst), .rdata(f1646_rdata));
  assign f1646_clk = clk;
  assign f1646_rst = rst;
  // Bindings to f1646

  // f1648
  logic [0:0] f1648_wen;
  logic [31:0] f1648_wdata;
  logic [0:0] f1648_clk;
  logic [0:0] f1648_rst;
  logic [31:0] f1648_rdata;
  sr_buffer_32_1 f1648(.wen(f1648_wen), .wdata(f1648_wdata), .clk(f1648_clk), .rst(f1648_rst), .rdata(f1648_rdata));
  assign f1648_clk = clk;
  assign f1648_rst = rst;
  // Bindings to f1648

  // f1650
  logic [0:0] f1650_wen;
  logic [31:0] f1650_wdata;
  logic [0:0] f1650_clk;
  logic [0:0] f1650_rst;
  logic [31:0] f1650_rdata;
  sr_buffer_32_1 f1650(.wen(f1650_wen), .wdata(f1650_wdata), .clk(f1650_clk), .rst(f1650_rst), .rdata(f1650_rdata));
  assign f1650_clk = clk;
  assign f1650_rst = rst;
  // Bindings to f1650

  // f1652
  logic [0:0] f1652_wen;
  logic [31:0] f1652_wdata;
  logic [0:0] f1652_clk;
  logic [0:0] f1652_rst;
  logic [31:0] f1652_rdata;
  sr_buffer_32_1 f1652(.wen(f1652_wen), .wdata(f1652_wdata), .clk(f1652_clk), .rst(f1652_rst), .rdata(f1652_rdata));
  assign f1652_clk = clk;
  assign f1652_rst = rst;
  // Bindings to f1652

  // f1654
  logic [0:0] f1654_wen;
  logic [31:0] f1654_wdata;
  logic [0:0] f1654_clk;
  logic [0:0] f1654_rst;
  logic [31:0] f1654_rdata;
  sr_buffer_32_1 f1654(.wen(f1654_wen), .wdata(f1654_wdata), .clk(f1654_clk), .rst(f1654_rst), .rdata(f1654_rdata));
  assign f1654_clk = clk;
  assign f1654_rst = rst;
  // Bindings to f1654

  // f1656
  logic [0:0] f1656_wen;
  logic [31:0] f1656_wdata;
  logic [0:0] f1656_clk;
  logic [0:0] f1656_rst;
  logic [31:0] f1656_rdata;
  sr_buffer_32_1 f1656(.wen(f1656_wen), .wdata(f1656_wdata), .clk(f1656_clk), .rst(f1656_rst), .rdata(f1656_rdata));
  assign f1656_clk = clk;
  assign f1656_rst = rst;
  // Bindings to f1656

  // f1658
  logic [0:0] f1658_wen;
  logic [31:0] f1658_wdata;
  logic [0:0] f1658_clk;
  logic [0:0] f1658_rst;
  logic [31:0] f1658_rdata;
  sr_buffer_32_1 f1658(.wen(f1658_wen), .wdata(f1658_wdata), .clk(f1658_clk), .rst(f1658_rst), .rdata(f1658_rdata));
  assign f1658_clk = clk;
  assign f1658_rst = rst;
  // Bindings to f1658

  // f1660
  logic [0:0] f1660_wen;
  logic [31:0] f1660_wdata;
  logic [0:0] f1660_clk;
  logic [0:0] f1660_rst;
  logic [31:0] f1660_rdata;
  sr_buffer_32_1 f1660(.wen(f1660_wen), .wdata(f1660_wdata), .clk(f1660_clk), .rst(f1660_rst), .rdata(f1660_rdata));
  assign f1660_clk = clk;
  assign f1660_rst = rst;
  // Bindings to f1660

  // f1662
  logic [0:0] f1662_wen;
  logic [31:0] f1662_wdata;
  logic [0:0] f1662_clk;
  logic [0:0] f1662_rst;
  logic [31:0] f1662_rdata;
  sr_buffer_32_1 f1662(.wen(f1662_wen), .wdata(f1662_wdata), .clk(f1662_clk), .rst(f1662_rst), .rdata(f1662_rdata));
  assign f1662_clk = clk;
  assign f1662_rst = rst;
  // Bindings to f1662

  // f1664
  logic [0:0] f1664_wen;
  logic [31:0] f1664_wdata;
  logic [0:0] f1664_clk;
  logic [0:0] f1664_rst;
  logic [31:0] f1664_rdata;
  sr_buffer_32_1 f1664(.wen(f1664_wen), .wdata(f1664_wdata), .clk(f1664_clk), .rst(f1664_rst), .rdata(f1664_rdata));
  assign f1664_clk = clk;
  assign f1664_rst = rst;
  // Bindings to f1664

  // f1666
  logic [0:0] f1666_wen;
  logic [31:0] f1666_wdata;
  logic [0:0] f1666_clk;
  logic [0:0] f1666_rst;
  logic [31:0] f1666_rdata;
  sr_buffer_32_1 f1666(.wen(f1666_wen), .wdata(f1666_wdata), .clk(f1666_clk), .rst(f1666_rst), .rdata(f1666_rdata));
  assign f1666_clk = clk;
  assign f1666_rst = rst;
  // Bindings to f1666

  // f1668
  logic [0:0] f1668_wen;
  logic [31:0] f1668_wdata;
  logic [0:0] f1668_clk;
  logic [0:0] f1668_rst;
  logic [31:0] f1668_rdata;
  sr_buffer_32_1 f1668(.wen(f1668_wen), .wdata(f1668_wdata), .clk(f1668_clk), .rst(f1668_rst), .rdata(f1668_rdata));
  assign f1668_clk = clk;
  assign f1668_rst = rst;
  // Bindings to f1668

  // f1670
  logic [0:0] f1670_wen;
  logic [31:0] f1670_wdata;
  logic [0:0] f1670_clk;
  logic [0:0] f1670_rst;
  logic [31:0] f1670_rdata;
  sr_buffer_32_1 f1670(.wen(f1670_wen), .wdata(f1670_wdata), .clk(f1670_clk), .rst(f1670_rst), .rdata(f1670_rdata));
  assign f1670_clk = clk;
  assign f1670_rst = rst;
  // Bindings to f1670

  // f1672
  logic [0:0] f1672_wen;
  logic [31:0] f1672_wdata;
  logic [0:0] f1672_clk;
  logic [0:0] f1672_rst;
  logic [31:0] f1672_rdata;
  sr_buffer_32_1 f1672(.wen(f1672_wen), .wdata(f1672_wdata), .clk(f1672_clk), .rst(f1672_rst), .rdata(f1672_rdata));
  assign f1672_clk = clk;
  assign f1672_rst = rst;
  // Bindings to f1672

  // f1674
  logic [0:0] f1674_wen;
  logic [31:0] f1674_wdata;
  logic [0:0] f1674_clk;
  logic [0:0] f1674_rst;
  logic [31:0] f1674_rdata;
  sr_buffer_32_1 f1674(.wen(f1674_wen), .wdata(f1674_wdata), .clk(f1674_clk), .rst(f1674_rst), .rdata(f1674_rdata));
  assign f1674_clk = clk;
  assign f1674_rst = rst;
  // Bindings to f1674

  // f1676
  logic [0:0] f1676_wen;
  logic [31:0] f1676_wdata;
  logic [0:0] f1676_clk;
  logic [0:0] f1676_rst;
  logic [31:0] f1676_rdata;
  sr_buffer_32_1 f1676(.wen(f1676_wen), .wdata(f1676_wdata), .clk(f1676_clk), .rst(f1676_rst), .rdata(f1676_rdata));
  assign f1676_clk = clk;
  assign f1676_rst = rst;
  // Bindings to f1676

  // f1678
  logic [0:0] f1678_wen;
  logic [31:0] f1678_wdata;
  logic [0:0] f1678_clk;
  logic [0:0] f1678_rst;
  logic [31:0] f1678_rdata;
  sr_buffer_32_1 f1678(.wen(f1678_wen), .wdata(f1678_wdata), .clk(f1678_clk), .rst(f1678_rst), .rdata(f1678_rdata));
  assign f1678_clk = clk;
  assign f1678_rst = rst;
  // Bindings to f1678

  // f1680
  logic [0:0] f1680_wen;
  logic [31:0] f1680_wdata;
  logic [0:0] f1680_clk;
  logic [0:0] f1680_rst;
  logic [31:0] f1680_rdata;
  sr_buffer_32_1 f1680(.wen(f1680_wen), .wdata(f1680_wdata), .clk(f1680_clk), .rst(f1680_rst), .rdata(f1680_rdata));
  assign f1680_clk = clk;
  assign f1680_rst = rst;
  // Bindings to f1680

  // f1682
  logic [0:0] f1682_wen;
  logic [31:0] f1682_wdata;
  logic [0:0] f1682_clk;
  logic [0:0] f1682_rst;
  logic [31:0] f1682_rdata;
  sr_buffer_32_1 f1682(.wen(f1682_wen), .wdata(f1682_wdata), .clk(f1682_clk), .rst(f1682_rst), .rdata(f1682_rdata));
  assign f1682_clk = clk;
  assign f1682_rst = rst;
  // Bindings to f1682

  // f1684
  logic [0:0] f1684_wen;
  logic [31:0] f1684_wdata;
  logic [0:0] f1684_clk;
  logic [0:0] f1684_rst;
  logic [31:0] f1684_rdata;
  sr_buffer_32_1 f1684(.wen(f1684_wen), .wdata(f1684_wdata), .clk(f1684_clk), .rst(f1684_rst), .rdata(f1684_rdata));
  assign f1684_clk = clk;
  assign f1684_rst = rst;
  // Bindings to f1684

  // f1686
  logic [0:0] f1686_wen;
  logic [31:0] f1686_wdata;
  logic [0:0] f1686_clk;
  logic [0:0] f1686_rst;
  logic [31:0] f1686_rdata;
  sr_buffer_32_1 f1686(.wen(f1686_wen), .wdata(f1686_wdata), .clk(f1686_clk), .rst(f1686_rst), .rdata(f1686_rdata));
  assign f1686_clk = clk;
  assign f1686_rst = rst;
  // Bindings to f1686

  // f1688
  logic [0:0] f1688_wen;
  logic [31:0] f1688_wdata;
  logic [0:0] f1688_clk;
  logic [0:0] f1688_rst;
  logic [31:0] f1688_rdata;
  sr_buffer_32_1 f1688(.wen(f1688_wen), .wdata(f1688_wdata), .clk(f1688_clk), .rst(f1688_rst), .rdata(f1688_rdata));
  assign f1688_clk = clk;
  assign f1688_rst = rst;
  // Bindings to f1688

  // f1690
  logic [0:0] f1690_wen;
  logic [31:0] f1690_wdata;
  logic [0:0] f1690_clk;
  logic [0:0] f1690_rst;
  logic [31:0] f1690_rdata;
  sr_buffer_32_1 f1690(.wen(f1690_wen), .wdata(f1690_wdata), .clk(f1690_clk), .rst(f1690_rst), .rdata(f1690_rdata));
  assign f1690_clk = clk;
  assign f1690_rst = rst;
  // Bindings to f1690

  // f1692
  logic [0:0] f1692_wen;
  logic [31:0] f1692_wdata;
  logic [0:0] f1692_clk;
  logic [0:0] f1692_rst;
  logic [31:0] f1692_rdata;
  sr_buffer_32_1 f1692(.wen(f1692_wen), .wdata(f1692_wdata), .clk(f1692_clk), .rst(f1692_rst), .rdata(f1692_rdata));
  assign f1692_clk = clk;
  assign f1692_rst = rst;
  // Bindings to f1692

  // f1694
  logic [0:0] f1694_wen;
  logic [31:0] f1694_wdata;
  logic [0:0] f1694_clk;
  logic [0:0] f1694_rst;
  logic [31:0] f1694_rdata;
  sr_buffer_32_1 f1694(.wen(f1694_wen), .wdata(f1694_wdata), .clk(f1694_clk), .rst(f1694_rst), .rdata(f1694_rdata));
  assign f1694_clk = clk;
  assign f1694_rst = rst;
  // Bindings to f1694

  // f1696
  logic [0:0] f1696_wen;
  logic [31:0] f1696_wdata;
  logic [0:0] f1696_clk;
  logic [0:0] f1696_rst;
  logic [31:0] f1696_rdata;
  sr_buffer_32_1 f1696(.wen(f1696_wen), .wdata(f1696_wdata), .clk(f1696_clk), .rst(f1696_rst), .rdata(f1696_rdata));
  assign f1696_clk = clk;
  assign f1696_rst = rst;
  // Bindings to f1696

  // f1698
  logic [0:0] f1698_wen;
  logic [31:0] f1698_wdata;
  logic [0:0] f1698_clk;
  logic [0:0] f1698_rst;
  logic [31:0] f1698_rdata;
  sr_buffer_32_1 f1698(.wen(f1698_wen), .wdata(f1698_wdata), .clk(f1698_clk), .rst(f1698_rst), .rdata(f1698_rdata));
  assign f1698_clk = clk;
  assign f1698_rst = rst;
  // Bindings to f1698

  // f1700
  logic [0:0] f1700_wen;
  logic [31:0] f1700_wdata;
  logic [0:0] f1700_clk;
  logic [0:0] f1700_rst;
  logic [31:0] f1700_rdata;
  sr_buffer_32_1 f1700(.wen(f1700_wen), .wdata(f1700_wdata), .clk(f1700_clk), .rst(f1700_rst), .rdata(f1700_rdata));
  assign f1700_clk = clk;
  assign f1700_rst = rst;
  // Bindings to f1700

  // f1702
  logic [0:0] f1702_wen;
  logic [31:0] f1702_wdata;
  logic [0:0] f1702_clk;
  logic [0:0] f1702_rst;
  logic [31:0] f1702_rdata;
  sr_buffer_32_1 f1702(.wen(f1702_wen), .wdata(f1702_wdata), .clk(f1702_clk), .rst(f1702_rst), .rdata(f1702_rdata));
  assign f1702_clk = clk;
  assign f1702_rst = rst;
  // Bindings to f1702

  // f1704
  logic [0:0] f1704_wen;
  logic [31:0] f1704_wdata;
  logic [0:0] f1704_clk;
  logic [0:0] f1704_rst;
  logic [31:0] f1704_rdata;
  sr_buffer_32_1 f1704(.wen(f1704_wen), .wdata(f1704_wdata), .clk(f1704_clk), .rst(f1704_rst), .rdata(f1704_rdata));
  assign f1704_clk = clk;
  assign f1704_rst = rst;
  // Bindings to f1704

  // f1706
  logic [0:0] f1706_wen;
  logic [31:0] f1706_wdata;
  logic [0:0] f1706_clk;
  logic [0:0] f1706_rst;
  logic [31:0] f1706_rdata;
  sr_buffer_32_1 f1706(.wen(f1706_wen), .wdata(f1706_wdata), .clk(f1706_clk), .rst(f1706_rst), .rdata(f1706_rdata));
  assign f1706_clk = clk;
  assign f1706_rst = rst;
  // Bindings to f1706

  // f1708
  logic [0:0] f1708_wen;
  logic [31:0] f1708_wdata;
  logic [0:0] f1708_clk;
  logic [0:0] f1708_rst;
  logic [31:0] f1708_rdata;
  sr_buffer_32_1 f1708(.wen(f1708_wen), .wdata(f1708_wdata), .clk(f1708_clk), .rst(f1708_rst), .rdata(f1708_rdata));
  assign f1708_clk = clk;
  assign f1708_rst = rst;
  // Bindings to f1708

  // f1710
  logic [0:0] f1710_wen;
  logic [31:0] f1710_wdata;
  logic [0:0] f1710_clk;
  logic [0:0] f1710_rst;
  logic [31:0] f1710_rdata;
  sr_buffer_32_1 f1710(.wen(f1710_wen), .wdata(f1710_wdata), .clk(f1710_clk), .rst(f1710_rst), .rdata(f1710_rdata));
  assign f1710_clk = clk;
  assign f1710_rst = rst;
  // Bindings to f1710

  // f1712
  logic [0:0] f1712_wen;
  logic [31:0] f1712_wdata;
  logic [0:0] f1712_clk;
  logic [0:0] f1712_rst;
  logic [31:0] f1712_rdata;
  sr_buffer_32_1 f1712(.wen(f1712_wen), .wdata(f1712_wdata), .clk(f1712_clk), .rst(f1712_rst), .rdata(f1712_rdata));
  assign f1712_clk = clk;
  assign f1712_rst = rst;
  // Bindings to f1712

  // f1714
  logic [0:0] f1714_wen;
  logic [31:0] f1714_wdata;
  logic [0:0] f1714_clk;
  logic [0:0] f1714_rst;
  logic [31:0] f1714_rdata;
  sr_buffer_32_1 f1714(.wen(f1714_wen), .wdata(f1714_wdata), .clk(f1714_clk), .rst(f1714_rst), .rdata(f1714_rdata));
  assign f1714_clk = clk;
  assign f1714_rst = rst;
  // Bindings to f1714

  // f1716
  logic [0:0] f1716_wen;
  logic [31:0] f1716_wdata;
  logic [0:0] f1716_clk;
  logic [0:0] f1716_rst;
  logic [31:0] f1716_rdata;
  sr_buffer_32_1 f1716(.wen(f1716_wen), .wdata(f1716_wdata), .clk(f1716_clk), .rst(f1716_rst), .rdata(f1716_rdata));
  assign f1716_clk = clk;
  assign f1716_rst = rst;
  // Bindings to f1716

  // f1718
  logic [0:0] f1718_wen;
  logic [31:0] f1718_wdata;
  logic [0:0] f1718_clk;
  logic [0:0] f1718_rst;
  logic [31:0] f1718_rdata;
  sr_buffer_32_1 f1718(.wen(f1718_wen), .wdata(f1718_wdata), .clk(f1718_clk), .rst(f1718_rst), .rdata(f1718_rdata));
  assign f1718_clk = clk;
  assign f1718_rst = rst;
  // Bindings to f1718

  // f1720
  logic [0:0] f1720_wen;
  logic [31:0] f1720_wdata;
  logic [0:0] f1720_clk;
  logic [0:0] f1720_rst;
  logic [31:0] f1720_rdata;
  sr_buffer_32_1 f1720(.wen(f1720_wen), .wdata(f1720_wdata), .clk(f1720_clk), .rst(f1720_rst), .rdata(f1720_rdata));
  assign f1720_clk = clk;
  assign f1720_rst = rst;
  // Bindings to f1720

  // f1722
  logic [0:0] f1722_wen;
  logic [31:0] f1722_wdata;
  logic [0:0] f1722_clk;
  logic [0:0] f1722_rst;
  logic [31:0] f1722_rdata;
  sr_buffer_32_1 f1722(.wen(f1722_wen), .wdata(f1722_wdata), .clk(f1722_clk), .rst(f1722_rst), .rdata(f1722_rdata));
  assign f1722_clk = clk;
  assign f1722_rst = rst;
  // Bindings to f1722

  // f1724
  logic [0:0] f1724_wen;
  logic [31:0] f1724_wdata;
  logic [0:0] f1724_clk;
  logic [0:0] f1724_rst;
  logic [31:0] f1724_rdata;
  sr_buffer_32_1 f1724(.wen(f1724_wen), .wdata(f1724_wdata), .clk(f1724_clk), .rst(f1724_rst), .rdata(f1724_rdata));
  assign f1724_clk = clk;
  assign f1724_rst = rst;
  // Bindings to f1724

  // f1726
  logic [0:0] f1726_wen;
  logic [31:0] f1726_wdata;
  logic [0:0] f1726_clk;
  logic [0:0] f1726_rst;
  logic [31:0] f1726_rdata;
  sr_buffer_32_1 f1726(.wen(f1726_wen), .wdata(f1726_wdata), .clk(f1726_clk), .rst(f1726_rst), .rdata(f1726_rdata));
  assign f1726_clk = clk;
  assign f1726_rst = rst;
  // Bindings to f1726

  // f1728
  logic [0:0] f1728_wen;
  logic [31:0] f1728_wdata;
  logic [0:0] f1728_clk;
  logic [0:0] f1728_rst;
  logic [31:0] f1728_rdata;
  sr_buffer_32_1 f1728(.wen(f1728_wen), .wdata(f1728_wdata), .clk(f1728_clk), .rst(f1728_rst), .rdata(f1728_rdata));
  assign f1728_clk = clk;
  assign f1728_rst = rst;
  // Bindings to f1728

  // f1730
  logic [0:0] f1730_wen;
  logic [31:0] f1730_wdata;
  logic [0:0] f1730_clk;
  logic [0:0] f1730_rst;
  logic [31:0] f1730_rdata;
  sr_buffer_32_1 f1730(.wen(f1730_wen), .wdata(f1730_wdata), .clk(f1730_clk), .rst(f1730_rst), .rdata(f1730_rdata));
  assign f1730_clk = clk;
  assign f1730_rst = rst;
  // Bindings to f1730

  // f1732
  logic [0:0] f1732_wen;
  logic [31:0] f1732_wdata;
  logic [0:0] f1732_clk;
  logic [0:0] f1732_rst;
  logic [31:0] f1732_rdata;
  sr_buffer_32_1 f1732(.wen(f1732_wen), .wdata(f1732_wdata), .clk(f1732_clk), .rst(f1732_rst), .rdata(f1732_rdata));
  assign f1732_clk = clk;
  assign f1732_rst = rst;
  // Bindings to f1732

  // f1734
  logic [0:0] f1734_wen;
  logic [31:0] f1734_wdata;
  logic [0:0] f1734_clk;
  logic [0:0] f1734_rst;
  logic [31:0] f1734_rdata;
  sr_buffer_32_1 f1734(.wen(f1734_wen), .wdata(f1734_wdata), .clk(f1734_clk), .rst(f1734_rst), .rdata(f1734_rdata));
  assign f1734_clk = clk;
  assign f1734_rst = rst;
  // Bindings to f1734

  // f1736
  logic [0:0] f1736_wen;
  logic [31:0] f1736_wdata;
  logic [0:0] f1736_clk;
  logic [0:0] f1736_rst;
  logic [31:0] f1736_rdata;
  sr_buffer_32_1 f1736(.wen(f1736_wen), .wdata(f1736_wdata), .clk(f1736_clk), .rst(f1736_rst), .rdata(f1736_rdata));
  assign f1736_clk = clk;
  assign f1736_rst = rst;
  // Bindings to f1736

  // f1738
  logic [0:0] f1738_wen;
  logic [31:0] f1738_wdata;
  logic [0:0] f1738_clk;
  logic [0:0] f1738_rst;
  logic [31:0] f1738_rdata;
  sr_buffer_32_1 f1738(.wen(f1738_wen), .wdata(f1738_wdata), .clk(f1738_clk), .rst(f1738_rst), .rdata(f1738_rdata));
  assign f1738_clk = clk;
  assign f1738_rst = rst;
  // Bindings to f1738

  // f1740
  logic [0:0] f1740_wen;
  logic [31:0] f1740_wdata;
  logic [0:0] f1740_clk;
  logic [0:0] f1740_rst;
  logic [31:0] f1740_rdata;
  sr_buffer_32_1 f1740(.wen(f1740_wen), .wdata(f1740_wdata), .clk(f1740_clk), .rst(f1740_rst), .rdata(f1740_rdata));
  assign f1740_clk = clk;
  assign f1740_rst = rst;
  // Bindings to f1740

  // f1742
  logic [0:0] f1742_wen;
  logic [31:0] f1742_wdata;
  logic [0:0] f1742_clk;
  logic [0:0] f1742_rst;
  logic [31:0] f1742_rdata;
  sr_buffer_32_1 f1742(.wen(f1742_wen), .wdata(f1742_wdata), .clk(f1742_clk), .rst(f1742_rst), .rdata(f1742_rdata));
  assign f1742_clk = clk;
  assign f1742_rst = rst;
  // Bindings to f1742

  // f1744
  logic [0:0] f1744_wen;
  logic [31:0] f1744_wdata;
  logic [0:0] f1744_clk;
  logic [0:0] f1744_rst;
  logic [31:0] f1744_rdata;
  sr_buffer_32_1 f1744(.wen(f1744_wen), .wdata(f1744_wdata), .clk(f1744_clk), .rst(f1744_rst), .rdata(f1744_rdata));
  assign f1744_clk = clk;
  assign f1744_rst = rst;
  // Bindings to f1744

  // f1746
  logic [0:0] f1746_wen;
  logic [31:0] f1746_wdata;
  logic [0:0] f1746_clk;
  logic [0:0] f1746_rst;
  logic [31:0] f1746_rdata;
  sr_buffer_32_1 f1746(.wen(f1746_wen), .wdata(f1746_wdata), .clk(f1746_clk), .rst(f1746_rst), .rdata(f1746_rdata));
  assign f1746_clk = clk;
  assign f1746_rst = rst;
  // Bindings to f1746

  // f1748
  logic [0:0] f1748_wen;
  logic [31:0] f1748_wdata;
  logic [0:0] f1748_clk;
  logic [0:0] f1748_rst;
  logic [31:0] f1748_rdata;
  sr_buffer_32_1 f1748(.wen(f1748_wen), .wdata(f1748_wdata), .clk(f1748_clk), .rst(f1748_rst), .rdata(f1748_rdata));
  assign f1748_clk = clk;
  assign f1748_rst = rst;
  // Bindings to f1748

  // f1750
  logic [0:0] f1750_wen;
  logic [31:0] f1750_wdata;
  logic [0:0] f1750_clk;
  logic [0:0] f1750_rst;
  logic [31:0] f1750_rdata;
  sr_buffer_32_1 f1750(.wen(f1750_wen), .wdata(f1750_wdata), .clk(f1750_clk), .rst(f1750_rst), .rdata(f1750_rdata));
  assign f1750_clk = clk;
  assign f1750_rst = rst;
  // Bindings to f1750

  // f1752
  logic [0:0] f1752_wen;
  logic [31:0] f1752_wdata;
  logic [0:0] f1752_clk;
  logic [0:0] f1752_rst;
  logic [31:0] f1752_rdata;
  sr_buffer_32_1 f1752(.wen(f1752_wen), .wdata(f1752_wdata), .clk(f1752_clk), .rst(f1752_rst), .rdata(f1752_rdata));
  assign f1752_clk = clk;
  assign f1752_rst = rst;
  // Bindings to f1752

  // f1754
  logic [0:0] f1754_wen;
  logic [31:0] f1754_wdata;
  logic [0:0] f1754_clk;
  logic [0:0] f1754_rst;
  logic [31:0] f1754_rdata;
  sr_buffer_32_1 f1754(.wen(f1754_wen), .wdata(f1754_wdata), .clk(f1754_clk), .rst(f1754_rst), .rdata(f1754_rdata));
  assign f1754_clk = clk;
  assign f1754_rst = rst;
  // Bindings to f1754

  // f1756
  logic [0:0] f1756_wen;
  logic [31:0] f1756_wdata;
  logic [0:0] f1756_clk;
  logic [0:0] f1756_rst;
  logic [31:0] f1756_rdata;
  sr_buffer_32_1 f1756(.wen(f1756_wen), .wdata(f1756_wdata), .clk(f1756_clk), .rst(f1756_rst), .rdata(f1756_rdata));
  assign f1756_clk = clk;
  assign f1756_rst = rst;
  // Bindings to f1756

  // f1758
  logic [0:0] f1758_wen;
  logic [31:0] f1758_wdata;
  logic [0:0] f1758_clk;
  logic [0:0] f1758_rst;
  logic [31:0] f1758_rdata;
  sr_buffer_32_1 f1758(.wen(f1758_wen), .wdata(f1758_wdata), .clk(f1758_clk), .rst(f1758_rst), .rdata(f1758_rdata));
  assign f1758_clk = clk;
  assign f1758_rst = rst;
  // Bindings to f1758

  // f1760
  logic [0:0] f1760_wen;
  logic [31:0] f1760_wdata;
  logic [0:0] f1760_clk;
  logic [0:0] f1760_rst;
  logic [31:0] f1760_rdata;
  sr_buffer_32_1 f1760(.wen(f1760_wen), .wdata(f1760_wdata), .clk(f1760_clk), .rst(f1760_rst), .rdata(f1760_rdata));
  assign f1760_clk = clk;
  assign f1760_rst = rst;
  // Bindings to f1760

  // f1762
  logic [0:0] f1762_wen;
  logic [31:0] f1762_wdata;
  logic [0:0] f1762_clk;
  logic [0:0] f1762_rst;
  logic [31:0] f1762_rdata;
  sr_buffer_32_1 f1762(.wen(f1762_wen), .wdata(f1762_wdata), .clk(f1762_clk), .rst(f1762_rst), .rdata(f1762_rdata));
  assign f1762_clk = clk;
  assign f1762_rst = rst;
  // Bindings to f1762

  // f1764
  logic [0:0] f1764_wen;
  logic [31:0] f1764_wdata;
  logic [0:0] f1764_clk;
  logic [0:0] f1764_rst;
  logic [31:0] f1764_rdata;
  sr_buffer_32_1 f1764(.wen(f1764_wen), .wdata(f1764_wdata), .clk(f1764_clk), .rst(f1764_rst), .rdata(f1764_rdata));
  assign f1764_clk = clk;
  assign f1764_rst = rst;
  // Bindings to f1764

  // f1766
  logic [0:0] f1766_wen;
  logic [31:0] f1766_wdata;
  logic [0:0] f1766_clk;
  logic [0:0] f1766_rst;
  logic [31:0] f1766_rdata;
  sr_buffer_32_1 f1766(.wen(f1766_wen), .wdata(f1766_wdata), .clk(f1766_clk), .rst(f1766_rst), .rdata(f1766_rdata));
  assign f1766_clk = clk;
  assign f1766_rst = rst;
  // Bindings to f1766

  // f1768
  logic [0:0] f1768_wen;
  logic [31:0] f1768_wdata;
  logic [0:0] f1768_clk;
  logic [0:0] f1768_rst;
  logic [31:0] f1768_rdata;
  sr_buffer_32_1 f1768(.wen(f1768_wen), .wdata(f1768_wdata), .clk(f1768_clk), .rst(f1768_rst), .rdata(f1768_rdata));
  assign f1768_clk = clk;
  assign f1768_rst = rst;
  // Bindings to f1768

  // f1770
  logic [0:0] f1770_wen;
  logic [31:0] f1770_wdata;
  logic [0:0] f1770_clk;
  logic [0:0] f1770_rst;
  logic [31:0] f1770_rdata;
  sr_buffer_32_1 f1770(.wen(f1770_wen), .wdata(f1770_wdata), .clk(f1770_clk), .rst(f1770_rst), .rdata(f1770_rdata));
  assign f1770_clk = clk;
  assign f1770_rst = rst;
  // Bindings to f1770

  // f1772
  logic [0:0] f1772_wen;
  logic [31:0] f1772_wdata;
  logic [0:0] f1772_clk;
  logic [0:0] f1772_rst;
  logic [31:0] f1772_rdata;
  sr_buffer_32_1 f1772(.wen(f1772_wen), .wdata(f1772_wdata), .clk(f1772_clk), .rst(f1772_rst), .rdata(f1772_rdata));
  assign f1772_clk = clk;
  assign f1772_rst = rst;
  // Bindings to f1772

  // f1774
  logic [0:0] f1774_wen;
  logic [31:0] f1774_wdata;
  logic [0:0] f1774_clk;
  logic [0:0] f1774_rst;
  logic [31:0] f1774_rdata;
  sr_buffer_32_1 f1774(.wen(f1774_wen), .wdata(f1774_wdata), .clk(f1774_clk), .rst(f1774_rst), .rdata(f1774_rdata));
  assign f1774_clk = clk;
  assign f1774_rst = rst;
  // Bindings to f1774

  // f1776
  logic [0:0] f1776_wen;
  logic [31:0] f1776_wdata;
  logic [0:0] f1776_clk;
  logic [0:0] f1776_rst;
  logic [31:0] f1776_rdata;
  sr_buffer_32_1 f1776(.wen(f1776_wen), .wdata(f1776_wdata), .clk(f1776_clk), .rst(f1776_rst), .rdata(f1776_rdata));
  assign f1776_clk = clk;
  assign f1776_rst = rst;
  // Bindings to f1776

  // f1778
  logic [0:0] f1778_wen;
  logic [31:0] f1778_wdata;
  logic [0:0] f1778_clk;
  logic [0:0] f1778_rst;
  logic [31:0] f1778_rdata;
  sr_buffer_32_1 f1778(.wen(f1778_wen), .wdata(f1778_wdata), .clk(f1778_clk), .rst(f1778_rst), .rdata(f1778_rdata));
  assign f1778_clk = clk;
  assign f1778_rst = rst;
  // Bindings to f1778

  // f1780
  logic [0:0] f1780_wen;
  logic [31:0] f1780_wdata;
  logic [0:0] f1780_clk;
  logic [0:0] f1780_rst;
  logic [31:0] f1780_rdata;
  sr_buffer_32_1 f1780(.wen(f1780_wen), .wdata(f1780_wdata), .clk(f1780_clk), .rst(f1780_rst), .rdata(f1780_rdata));
  assign f1780_clk = clk;
  assign f1780_rst = rst;
  // Bindings to f1780

  // f1782
  logic [0:0] f1782_wen;
  logic [31:0] f1782_wdata;
  logic [0:0] f1782_clk;
  logic [0:0] f1782_rst;
  logic [31:0] f1782_rdata;
  sr_buffer_32_1 f1782(.wen(f1782_wen), .wdata(f1782_wdata), .clk(f1782_clk), .rst(f1782_rst), .rdata(f1782_rdata));
  assign f1782_clk = clk;
  assign f1782_rst = rst;
  // Bindings to f1782

  // f1784
  logic [0:0] f1784_wen;
  logic [31:0] f1784_wdata;
  logic [0:0] f1784_clk;
  logic [0:0] f1784_rst;
  logic [31:0] f1784_rdata;
  sr_buffer_32_1 f1784(.wen(f1784_wen), .wdata(f1784_wdata), .clk(f1784_clk), .rst(f1784_rst), .rdata(f1784_rdata));
  assign f1784_clk = clk;
  assign f1784_rst = rst;
  // Bindings to f1784

  // f1786
  logic [0:0] f1786_wen;
  logic [31:0] f1786_wdata;
  logic [0:0] f1786_clk;
  logic [0:0] f1786_rst;
  logic [31:0] f1786_rdata;
  sr_buffer_32_1 f1786(.wen(f1786_wen), .wdata(f1786_wdata), .clk(f1786_clk), .rst(f1786_rst), .rdata(f1786_rdata));
  assign f1786_clk = clk;
  assign f1786_rst = rst;
  // Bindings to f1786

  // f1788
  logic [0:0] f1788_wen;
  logic [31:0] f1788_wdata;
  logic [0:0] f1788_clk;
  logic [0:0] f1788_rst;
  logic [31:0] f1788_rdata;
  sr_buffer_32_1 f1788(.wen(f1788_wen), .wdata(f1788_wdata), .clk(f1788_clk), .rst(f1788_rst), .rdata(f1788_rdata));
  assign f1788_clk = clk;
  assign f1788_rst = rst;
  // Bindings to f1788

  // f1790
  logic [0:0] f1790_wen;
  logic [31:0] f1790_wdata;
  logic [0:0] f1790_clk;
  logic [0:0] f1790_rst;
  logic [31:0] f1790_rdata;
  sr_buffer_32_1 f1790(.wen(f1790_wen), .wdata(f1790_wdata), .clk(f1790_clk), .rst(f1790_rst), .rdata(f1790_rdata));
  assign f1790_clk = clk;
  assign f1790_rst = rst;
  // Bindings to f1790

  // f1792
  logic [0:0] f1792_wen;
  logic [31:0] f1792_wdata;
  logic [0:0] f1792_clk;
  logic [0:0] f1792_rst;
  logic [31:0] f1792_rdata;
  sr_buffer_32_1 f1792(.wen(f1792_wen), .wdata(f1792_wdata), .clk(f1792_clk), .rst(f1792_rst), .rdata(f1792_rdata));
  assign f1792_clk = clk;
  assign f1792_rst = rst;
  // Bindings to f1792

  // f1794
  logic [0:0] f1794_wen;
  logic [31:0] f1794_wdata;
  logic [0:0] f1794_clk;
  logic [0:0] f1794_rst;
  logic [31:0] f1794_rdata;
  sr_buffer_32_1 f1794(.wen(f1794_wen), .wdata(f1794_wdata), .clk(f1794_clk), .rst(f1794_rst), .rdata(f1794_rdata));
  assign f1794_clk = clk;
  assign f1794_rst = rst;
  // Bindings to f1794

  // f1796
  logic [0:0] f1796_wen;
  logic [31:0] f1796_wdata;
  logic [0:0] f1796_clk;
  logic [0:0] f1796_rst;
  logic [31:0] f1796_rdata;
  sr_buffer_32_1 f1796(.wen(f1796_wen), .wdata(f1796_wdata), .clk(f1796_clk), .rst(f1796_rst), .rdata(f1796_rdata));
  assign f1796_clk = clk;
  assign f1796_rst = rst;
  // Bindings to f1796

  // f1798
  logic [0:0] f1798_wen;
  logic [31:0] f1798_wdata;
  logic [0:0] f1798_clk;
  logic [0:0] f1798_rst;
  logic [31:0] f1798_rdata;
  sr_buffer_32_1 f1798(.wen(f1798_wen), .wdata(f1798_wdata), .clk(f1798_clk), .rst(f1798_rst), .rdata(f1798_rdata));
  assign f1798_clk = clk;
  assign f1798_rst = rst;
  // Bindings to f1798

  // f1800
  logic [0:0] f1800_wen;
  logic [31:0] f1800_wdata;
  logic [0:0] f1800_clk;
  logic [0:0] f1800_rst;
  logic [31:0] f1800_rdata;
  sr_buffer_32_1 f1800(.wen(f1800_wen), .wdata(f1800_wdata), .clk(f1800_clk), .rst(f1800_rst), .rdata(f1800_rdata));
  assign f1800_clk = clk;
  assign f1800_rst = rst;
  // Bindings to f1800

  // f1802
  logic [0:0] f1802_wen;
  logic [31:0] f1802_wdata;
  logic [0:0] f1802_clk;
  logic [0:0] f1802_rst;
  logic [31:0] f1802_rdata;
  sr_buffer_32_1 f1802(.wen(f1802_wen), .wdata(f1802_wdata), .clk(f1802_clk), .rst(f1802_rst), .rdata(f1802_rdata));
  assign f1802_clk = clk;
  assign f1802_rst = rst;
  // Bindings to f1802

  // f1804
  logic [0:0] f1804_wen;
  logic [31:0] f1804_wdata;
  logic [0:0] f1804_clk;
  logic [0:0] f1804_rst;
  logic [31:0] f1804_rdata;
  sr_buffer_32_1 f1804(.wen(f1804_wen), .wdata(f1804_wdata), .clk(f1804_clk), .rst(f1804_rst), .rdata(f1804_rdata));
  assign f1804_clk = clk;
  assign f1804_rst = rst;
  // Bindings to f1804

  // f1806
  logic [0:0] f1806_wen;
  logic [31:0] f1806_wdata;
  logic [0:0] f1806_clk;
  logic [0:0] f1806_rst;
  logic [31:0] f1806_rdata;
  sr_buffer_32_1 f1806(.wen(f1806_wen), .wdata(f1806_wdata), .clk(f1806_clk), .rst(f1806_rst), .rdata(f1806_rdata));
  assign f1806_clk = clk;
  assign f1806_rst = rst;
  // Bindings to f1806

  // f1808
  logic [0:0] f1808_wen;
  logic [31:0] f1808_wdata;
  logic [0:0] f1808_clk;
  logic [0:0] f1808_rst;
  logic [31:0] f1808_rdata;
  sr_buffer_32_1 f1808(.wen(f1808_wen), .wdata(f1808_wdata), .clk(f1808_clk), .rst(f1808_rst), .rdata(f1808_rdata));
  assign f1808_clk = clk;
  assign f1808_rst = rst;
  // Bindings to f1808

  // f1810
  logic [0:0] f1810_wen;
  logic [31:0] f1810_wdata;
  logic [0:0] f1810_clk;
  logic [0:0] f1810_rst;
  logic [31:0] f1810_rdata;
  sr_buffer_32_1 f1810(.wen(f1810_wen), .wdata(f1810_wdata), .clk(f1810_clk), .rst(f1810_rst), .rdata(f1810_rdata));
  assign f1810_clk = clk;
  assign f1810_rst = rst;
  // Bindings to f1810

  // f1812
  logic [0:0] f1812_wen;
  logic [31:0] f1812_wdata;
  logic [0:0] f1812_clk;
  logic [0:0] f1812_rst;
  logic [31:0] f1812_rdata;
  sr_buffer_32_1 f1812(.wen(f1812_wen), .wdata(f1812_wdata), .clk(f1812_clk), .rst(f1812_rst), .rdata(f1812_rdata));
  assign f1812_clk = clk;
  assign f1812_rst = rst;
  // Bindings to f1812

  // f1814
  logic [0:0] f1814_wen;
  logic [31:0] f1814_wdata;
  logic [0:0] f1814_clk;
  logic [0:0] f1814_rst;
  logic [31:0] f1814_rdata;
  sr_buffer_32_1 f1814(.wen(f1814_wen), .wdata(f1814_wdata), .clk(f1814_clk), .rst(f1814_rst), .rdata(f1814_rdata));
  assign f1814_clk = clk;
  assign f1814_rst = rst;
  // Bindings to f1814

  // f1816
  logic [0:0] f1816_wen;
  logic [31:0] f1816_wdata;
  logic [0:0] f1816_clk;
  logic [0:0] f1816_rst;
  logic [31:0] f1816_rdata;
  sr_buffer_32_1 f1816(.wen(f1816_wen), .wdata(f1816_wdata), .clk(f1816_clk), .rst(f1816_rst), .rdata(f1816_rdata));
  assign f1816_clk = clk;
  assign f1816_rst = rst;
  // Bindings to f1816

  // f1818
  logic [0:0] f1818_wen;
  logic [31:0] f1818_wdata;
  logic [0:0] f1818_clk;
  logic [0:0] f1818_rst;
  logic [31:0] f1818_rdata;
  sr_buffer_32_1 f1818(.wen(f1818_wen), .wdata(f1818_wdata), .clk(f1818_clk), .rst(f1818_rst), .rdata(f1818_rdata));
  assign f1818_clk = clk;
  assign f1818_rst = rst;
  // Bindings to f1818

  // f1820
  logic [0:0] f1820_wen;
  logic [31:0] f1820_wdata;
  logic [0:0] f1820_clk;
  logic [0:0] f1820_rst;
  logic [31:0] f1820_rdata;
  sr_buffer_32_1 f1820(.wen(f1820_wen), .wdata(f1820_wdata), .clk(f1820_clk), .rst(f1820_rst), .rdata(f1820_rdata));
  assign f1820_clk = clk;
  assign f1820_rst = rst;
  // Bindings to f1820

  // f1822
  logic [0:0] f1822_wen;
  logic [31:0] f1822_wdata;
  logic [0:0] f1822_clk;
  logic [0:0] f1822_rst;
  logic [31:0] f1822_rdata;
  sr_buffer_32_1 f1822(.wen(f1822_wen), .wdata(f1822_wdata), .clk(f1822_clk), .rst(f1822_rst), .rdata(f1822_rdata));
  assign f1822_clk = clk;
  assign f1822_rst = rst;
  // Bindings to f1822

  // f1824
  logic [0:0] f1824_wen;
  logic [31:0] f1824_wdata;
  logic [0:0] f1824_clk;
  logic [0:0] f1824_rst;
  logic [31:0] f1824_rdata;
  sr_buffer_32_1 f1824(.wen(f1824_wen), .wdata(f1824_wdata), .clk(f1824_clk), .rst(f1824_rst), .rdata(f1824_rdata));
  assign f1824_clk = clk;
  assign f1824_rst = rst;
  // Bindings to f1824

  // f1826
  logic [0:0] f1826_wen;
  logic [31:0] f1826_wdata;
  logic [0:0] f1826_clk;
  logic [0:0] f1826_rst;
  logic [31:0] f1826_rdata;
  sr_buffer_32_1 f1826(.wen(f1826_wen), .wdata(f1826_wdata), .clk(f1826_clk), .rst(f1826_rst), .rdata(f1826_rdata));
  assign f1826_clk = clk;
  assign f1826_rst = rst;
  // Bindings to f1826

  // f1828
  logic [0:0] f1828_wen;
  logic [31:0] f1828_wdata;
  logic [0:0] f1828_clk;
  logic [0:0] f1828_rst;
  logic [31:0] f1828_rdata;
  sr_buffer_32_1 f1828(.wen(f1828_wen), .wdata(f1828_wdata), .clk(f1828_clk), .rst(f1828_rst), .rdata(f1828_rdata));
  assign f1828_clk = clk;
  assign f1828_rst = rst;
  // Bindings to f1828

  // f1830
  logic [0:0] f1830_wen;
  logic [31:0] f1830_wdata;
  logic [0:0] f1830_clk;
  logic [0:0] f1830_rst;
  logic [31:0] f1830_rdata;
  sr_buffer_32_1 f1830(.wen(f1830_wen), .wdata(f1830_wdata), .clk(f1830_clk), .rst(f1830_rst), .rdata(f1830_rdata));
  assign f1830_clk = clk;
  assign f1830_rst = rst;
  // Bindings to f1830

  // f1832
  logic [0:0] f1832_wen;
  logic [31:0] f1832_wdata;
  logic [0:0] f1832_clk;
  logic [0:0] f1832_rst;
  logic [31:0] f1832_rdata;
  sr_buffer_32_1 f1832(.wen(f1832_wen), .wdata(f1832_wdata), .clk(f1832_clk), .rst(f1832_rst), .rdata(f1832_rdata));
  assign f1832_clk = clk;
  assign f1832_rst = rst;
  // Bindings to f1832

  // f1834
  logic [0:0] f1834_wen;
  logic [31:0] f1834_wdata;
  logic [0:0] f1834_clk;
  logic [0:0] f1834_rst;
  logic [31:0] f1834_rdata;
  sr_buffer_32_1 f1834(.wen(f1834_wen), .wdata(f1834_wdata), .clk(f1834_clk), .rst(f1834_rst), .rdata(f1834_rdata));
  assign f1834_clk = clk;
  assign f1834_rst = rst;
  // Bindings to f1834

  // f1836
  logic [0:0] f1836_wen;
  logic [31:0] f1836_wdata;
  logic [0:0] f1836_clk;
  logic [0:0] f1836_rst;
  logic [31:0] f1836_rdata;
  sr_buffer_32_1 f1836(.wen(f1836_wen), .wdata(f1836_wdata), .clk(f1836_clk), .rst(f1836_rst), .rdata(f1836_rdata));
  assign f1836_clk = clk;
  assign f1836_rst = rst;
  // Bindings to f1836

  // f1838
  logic [0:0] f1838_wen;
  logic [31:0] f1838_wdata;
  logic [0:0] f1838_clk;
  logic [0:0] f1838_rst;
  logic [31:0] f1838_rdata;
  sr_buffer_32_1 f1838(.wen(f1838_wen), .wdata(f1838_wdata), .clk(f1838_clk), .rst(f1838_rst), .rdata(f1838_rdata));
  assign f1838_clk = clk;
  assign f1838_rst = rst;
  // Bindings to f1838

  // f1840
  logic [0:0] f1840_wen;
  logic [31:0] f1840_wdata;
  logic [0:0] f1840_clk;
  logic [0:0] f1840_rst;
  logic [31:0] f1840_rdata;
  sr_buffer_32_1 f1840(.wen(f1840_wen), .wdata(f1840_wdata), .clk(f1840_clk), .rst(f1840_rst), .rdata(f1840_rdata));
  assign f1840_clk = clk;
  assign f1840_rst = rst;
  // Bindings to f1840

  // f1842
  logic [0:0] f1842_wen;
  logic [31:0] f1842_wdata;
  logic [0:0] f1842_clk;
  logic [0:0] f1842_rst;
  logic [31:0] f1842_rdata;
  sr_buffer_32_1 f1842(.wen(f1842_wen), .wdata(f1842_wdata), .clk(f1842_clk), .rst(f1842_rst), .rdata(f1842_rdata));
  assign f1842_clk = clk;
  assign f1842_rst = rst;
  // Bindings to f1842

  // f1844
  logic [0:0] f1844_wen;
  logic [31:0] f1844_wdata;
  logic [0:0] f1844_clk;
  logic [0:0] f1844_rst;
  logic [31:0] f1844_rdata;
  sr_buffer_32_1 f1844(.wen(f1844_wen), .wdata(f1844_wdata), .clk(f1844_clk), .rst(f1844_rst), .rdata(f1844_rdata));
  assign f1844_clk = clk;
  assign f1844_rst = rst;
  // Bindings to f1844

  // f1846
  logic [0:0] f1846_wen;
  logic [31:0] f1846_wdata;
  logic [0:0] f1846_clk;
  logic [0:0] f1846_rst;
  logic [31:0] f1846_rdata;
  sr_buffer_32_1 f1846(.wen(f1846_wen), .wdata(f1846_wdata), .clk(f1846_clk), .rst(f1846_rst), .rdata(f1846_rdata));
  assign f1846_clk = clk;
  assign f1846_rst = rst;
  // Bindings to f1846

  // f1848
  logic [0:0] f1848_wen;
  logic [31:0] f1848_wdata;
  logic [0:0] f1848_clk;
  logic [0:0] f1848_rst;
  logic [31:0] f1848_rdata;
  sr_buffer_32_1 f1848(.wen(f1848_wen), .wdata(f1848_wdata), .clk(f1848_clk), .rst(f1848_rst), .rdata(f1848_rdata));
  assign f1848_clk = clk;
  assign f1848_rst = rst;
  // Bindings to f1848

  // f1850
  logic [0:0] f1850_wen;
  logic [31:0] f1850_wdata;
  logic [0:0] f1850_clk;
  logic [0:0] f1850_rst;
  logic [31:0] f1850_rdata;
  sr_buffer_32_1 f1850(.wen(f1850_wen), .wdata(f1850_wdata), .clk(f1850_clk), .rst(f1850_rst), .rdata(f1850_rdata));
  assign f1850_clk = clk;
  assign f1850_rst = rst;
  // Bindings to f1850

  // f1852
  logic [0:0] f1852_wen;
  logic [31:0] f1852_wdata;
  logic [0:0] f1852_clk;
  logic [0:0] f1852_rst;
  logic [31:0] f1852_rdata;
  sr_buffer_32_1 f1852(.wen(f1852_wen), .wdata(f1852_wdata), .clk(f1852_clk), .rst(f1852_rst), .rdata(f1852_rdata));
  assign f1852_clk = clk;
  assign f1852_rst = rst;
  // Bindings to f1852

  // f1854
  logic [0:0] f1854_wen;
  logic [31:0] f1854_wdata;
  logic [0:0] f1854_clk;
  logic [0:0] f1854_rst;
  logic [31:0] f1854_rdata;
  sr_buffer_32_1 f1854(.wen(f1854_wen), .wdata(f1854_wdata), .clk(f1854_clk), .rst(f1854_rst), .rdata(f1854_rdata));
  assign f1854_clk = clk;
  assign f1854_rst = rst;
  // Bindings to f1854

  // f1856
  logic [0:0] f1856_wen;
  logic [31:0] f1856_wdata;
  logic [0:0] f1856_clk;
  logic [0:0] f1856_rst;
  logic [31:0] f1856_rdata;
  sr_buffer_32_1 f1856(.wen(f1856_wen), .wdata(f1856_wdata), .clk(f1856_clk), .rst(f1856_rst), .rdata(f1856_rdata));
  assign f1856_clk = clk;
  assign f1856_rst = rst;
  // Bindings to f1856

  // f1858
  logic [0:0] f1858_wen;
  logic [31:0] f1858_wdata;
  logic [0:0] f1858_clk;
  logic [0:0] f1858_rst;
  logic [31:0] f1858_rdata;
  sr_buffer_32_1 f1858(.wen(f1858_wen), .wdata(f1858_wdata), .clk(f1858_clk), .rst(f1858_rst), .rdata(f1858_rdata));
  assign f1858_clk = clk;
  assign f1858_rst = rst;
  // Bindings to f1858

  // f1860
  logic [0:0] f1860_wen;
  logic [31:0] f1860_wdata;
  logic [0:0] f1860_clk;
  logic [0:0] f1860_rst;
  logic [31:0] f1860_rdata;
  sr_buffer_32_1 f1860(.wen(f1860_wen), .wdata(f1860_wdata), .clk(f1860_clk), .rst(f1860_rst), .rdata(f1860_rdata));
  assign f1860_clk = clk;
  assign f1860_rst = rst;
  // Bindings to f1860

  // f1862
  logic [0:0] f1862_wen;
  logic [31:0] f1862_wdata;
  logic [0:0] f1862_clk;
  logic [0:0] f1862_rst;
  logic [31:0] f1862_rdata;
  sr_buffer_32_1 f1862(.wen(f1862_wen), .wdata(f1862_wdata), .clk(f1862_clk), .rst(f1862_rst), .rdata(f1862_rdata));
  assign f1862_clk = clk;
  assign f1862_rst = rst;
  // Bindings to f1862

  // f1864
  logic [0:0] f1864_wen;
  logic [31:0] f1864_wdata;
  logic [0:0] f1864_clk;
  logic [0:0] f1864_rst;
  logic [31:0] f1864_rdata;
  sr_buffer_32_1 f1864(.wen(f1864_wen), .wdata(f1864_wdata), .clk(f1864_clk), .rst(f1864_rst), .rdata(f1864_rdata));
  assign f1864_clk = clk;
  assign f1864_rst = rst;
  // Bindings to f1864

  // f1866
  logic [0:0] f1866_wen;
  logic [31:0] f1866_wdata;
  logic [0:0] f1866_clk;
  logic [0:0] f1866_rst;
  logic [31:0] f1866_rdata;
  sr_buffer_32_1 f1866(.wen(f1866_wen), .wdata(f1866_wdata), .clk(f1866_clk), .rst(f1866_rst), .rdata(f1866_rdata));
  assign f1866_clk = clk;
  assign f1866_rst = rst;
  // Bindings to f1866

  // f1868
  logic [0:0] f1868_wen;
  logic [31:0] f1868_wdata;
  logic [0:0] f1868_clk;
  logic [0:0] f1868_rst;
  logic [31:0] f1868_rdata;
  sr_buffer_32_1 f1868(.wen(f1868_wen), .wdata(f1868_wdata), .clk(f1868_clk), .rst(f1868_rst), .rdata(f1868_rdata));
  assign f1868_clk = clk;
  assign f1868_rst = rst;
  // Bindings to f1868

  // f1870
  logic [0:0] f1870_wen;
  logic [31:0] f1870_wdata;
  logic [0:0] f1870_clk;
  logic [0:0] f1870_rst;
  logic [31:0] f1870_rdata;
  sr_buffer_32_1 f1870(.wen(f1870_wen), .wdata(f1870_wdata), .clk(f1870_clk), .rst(f1870_rst), .rdata(f1870_rdata));
  assign f1870_clk = clk;
  assign f1870_rst = rst;
  // Bindings to f1870

  // f1872
  logic [0:0] f1872_wen;
  logic [31:0] f1872_wdata;
  logic [0:0] f1872_clk;
  logic [0:0] f1872_rst;
  logic [31:0] f1872_rdata;
  sr_buffer_32_1 f1872(.wen(f1872_wen), .wdata(f1872_wdata), .clk(f1872_clk), .rst(f1872_rst), .rdata(f1872_rdata));
  assign f1872_clk = clk;
  assign f1872_rst = rst;
  // Bindings to f1872

  // f1874
  logic [0:0] f1874_wen;
  logic [31:0] f1874_wdata;
  logic [0:0] f1874_clk;
  logic [0:0] f1874_rst;
  logic [31:0] f1874_rdata;
  sr_buffer_32_1 f1874(.wen(f1874_wen), .wdata(f1874_wdata), .clk(f1874_clk), .rst(f1874_rst), .rdata(f1874_rdata));
  assign f1874_clk = clk;
  assign f1874_rst = rst;
  // Bindings to f1874

  // f1876
  logic [0:0] f1876_wen;
  logic [31:0] f1876_wdata;
  logic [0:0] f1876_clk;
  logic [0:0] f1876_rst;
  logic [31:0] f1876_rdata;
  sr_buffer_32_1 f1876(.wen(f1876_wen), .wdata(f1876_wdata), .clk(f1876_clk), .rst(f1876_rst), .rdata(f1876_rdata));
  assign f1876_clk = clk;
  assign f1876_rst = rst;
  // Bindings to f1876

  // f1878
  logic [0:0] f1878_wen;
  logic [31:0] f1878_wdata;
  logic [0:0] f1878_clk;
  logic [0:0] f1878_rst;
  logic [31:0] f1878_rdata;
  sr_buffer_32_1 f1878(.wen(f1878_wen), .wdata(f1878_wdata), .clk(f1878_clk), .rst(f1878_rst), .rdata(f1878_rdata));
  assign f1878_clk = clk;
  assign f1878_rst = rst;
  // Bindings to f1878

  // f1880
  logic [0:0] f1880_wen;
  logic [31:0] f1880_wdata;
  logic [0:0] f1880_clk;
  logic [0:0] f1880_rst;
  logic [31:0] f1880_rdata;
  sr_buffer_32_1 f1880(.wen(f1880_wen), .wdata(f1880_wdata), .clk(f1880_clk), .rst(f1880_rst), .rdata(f1880_rdata));
  assign f1880_clk = clk;
  assign f1880_rst = rst;
  // Bindings to f1880

  // f1882
  logic [0:0] f1882_wen;
  logic [31:0] f1882_wdata;
  logic [0:0] f1882_clk;
  logic [0:0] f1882_rst;
  logic [31:0] f1882_rdata;
  sr_buffer_32_1 f1882(.wen(f1882_wen), .wdata(f1882_wdata), .clk(f1882_clk), .rst(f1882_rst), .rdata(f1882_rdata));
  assign f1882_clk = clk;
  assign f1882_rst = rst;
  // Bindings to f1882

  // f1884
  logic [0:0] f1884_wen;
  logic [31:0] f1884_wdata;
  logic [0:0] f1884_clk;
  logic [0:0] f1884_rst;
  logic [31:0] f1884_rdata;
  sr_buffer_32_1 f1884(.wen(f1884_wen), .wdata(f1884_wdata), .clk(f1884_clk), .rst(f1884_rst), .rdata(f1884_rdata));
  assign f1884_clk = clk;
  assign f1884_rst = rst;
  // Bindings to f1884

  // f1886
  logic [0:0] f1886_wen;
  logic [31:0] f1886_wdata;
  logic [0:0] f1886_clk;
  logic [0:0] f1886_rst;
  logic [31:0] f1886_rdata;
  sr_buffer_32_1 f1886(.wen(f1886_wen), .wdata(f1886_wdata), .clk(f1886_clk), .rst(f1886_rst), .rdata(f1886_rdata));
  assign f1886_clk = clk;
  assign f1886_rst = rst;
  // Bindings to f1886

  // f1888
  logic [0:0] f1888_wen;
  logic [31:0] f1888_wdata;
  logic [0:0] f1888_clk;
  logic [0:0] f1888_rst;
  logic [31:0] f1888_rdata;
  sr_buffer_32_1 f1888(.wen(f1888_wen), .wdata(f1888_wdata), .clk(f1888_clk), .rst(f1888_rst), .rdata(f1888_rdata));
  assign f1888_clk = clk;
  assign f1888_rst = rst;
  // Bindings to f1888

  // f1890
  logic [0:0] f1890_wen;
  logic [31:0] f1890_wdata;
  logic [0:0] f1890_clk;
  logic [0:0] f1890_rst;
  logic [31:0] f1890_rdata;
  sr_buffer_32_1 f1890(.wen(f1890_wen), .wdata(f1890_wdata), .clk(f1890_clk), .rst(f1890_rst), .rdata(f1890_rdata));
  assign f1890_clk = clk;
  assign f1890_rst = rst;
  // Bindings to f1890

  // f1892
  logic [0:0] f1892_wen;
  logic [31:0] f1892_wdata;
  logic [0:0] f1892_clk;
  logic [0:0] f1892_rst;
  logic [31:0] f1892_rdata;
  sr_buffer_32_1 f1892(.wen(f1892_wen), .wdata(f1892_wdata), .clk(f1892_clk), .rst(f1892_rst), .rdata(f1892_rdata));
  assign f1892_clk = clk;
  assign f1892_rst = rst;
  // Bindings to f1892

  // f1894
  logic [0:0] f1894_wen;
  logic [31:0] f1894_wdata;
  logic [0:0] f1894_clk;
  logic [0:0] f1894_rst;
  logic [31:0] f1894_rdata;
  sr_buffer_32_1 f1894(.wen(f1894_wen), .wdata(f1894_wdata), .clk(f1894_clk), .rst(f1894_rst), .rdata(f1894_rdata));
  assign f1894_clk = clk;
  assign f1894_rst = rst;
  // Bindings to f1894

  // f1896
  logic [0:0] f1896_wen;
  logic [31:0] f1896_wdata;
  logic [0:0] f1896_clk;
  logic [0:0] f1896_rst;
  logic [31:0] f1896_rdata;
  sr_buffer_32_1 f1896(.wen(f1896_wen), .wdata(f1896_wdata), .clk(f1896_clk), .rst(f1896_rst), .rdata(f1896_rdata));
  assign f1896_clk = clk;
  assign f1896_rst = rst;
  // Bindings to f1896

  // f1898
  logic [0:0] f1898_wen;
  logic [31:0] f1898_wdata;
  logic [0:0] f1898_clk;
  logic [0:0] f1898_rst;
  logic [31:0] f1898_rdata;
  sr_buffer_32_1 f1898(.wen(f1898_wen), .wdata(f1898_wdata), .clk(f1898_clk), .rst(f1898_rst), .rdata(f1898_rdata));
  assign f1898_clk = clk;
  assign f1898_rst = rst;
  // Bindings to f1898

  // f1900
  logic [0:0] f1900_wen;
  logic [31:0] f1900_wdata;
  logic [0:0] f1900_clk;
  logic [0:0] f1900_rst;
  logic [31:0] f1900_rdata;
  sr_buffer_32_1 f1900(.wen(f1900_wen), .wdata(f1900_wdata), .clk(f1900_clk), .rst(f1900_rst), .rdata(f1900_rdata));
  assign f1900_clk = clk;
  assign f1900_rst = rst;
  // Bindings to f1900

  // f1902
  logic [0:0] f1902_wen;
  logic [31:0] f1902_wdata;
  logic [0:0] f1902_clk;
  logic [0:0] f1902_rst;
  logic [31:0] f1902_rdata;
  sr_buffer_32_1 f1902(.wen(f1902_wen), .wdata(f1902_wdata), .clk(f1902_clk), .rst(f1902_rst), .rdata(f1902_rdata));
  assign f1902_clk = clk;
  assign f1902_rst = rst;
  // Bindings to f1902

  // f1904
  logic [0:0] f1904_wen;
  logic [31:0] f1904_wdata;
  logic [0:0] f1904_clk;
  logic [0:0] f1904_rst;
  logic [31:0] f1904_rdata;
  sr_buffer_32_1 f1904(.wen(f1904_wen), .wdata(f1904_wdata), .clk(f1904_clk), .rst(f1904_rst), .rdata(f1904_rdata));
  assign f1904_clk = clk;
  assign f1904_rst = rst;
  // Bindings to f1904

  // f1906
  logic [0:0] f1906_wen;
  logic [31:0] f1906_wdata;
  logic [0:0] f1906_clk;
  logic [0:0] f1906_rst;
  logic [31:0] f1906_rdata;
  sr_buffer_32_1 f1906(.wen(f1906_wen), .wdata(f1906_wdata), .clk(f1906_clk), .rst(f1906_rst), .rdata(f1906_rdata));
  assign f1906_clk = clk;
  assign f1906_rst = rst;
  // Bindings to f1906

  // f1908
  logic [0:0] f1908_wen;
  logic [31:0] f1908_wdata;
  logic [0:0] f1908_clk;
  logic [0:0] f1908_rst;
  logic [31:0] f1908_rdata;
  sr_buffer_32_1 f1908(.wen(f1908_wen), .wdata(f1908_wdata), .clk(f1908_clk), .rst(f1908_rst), .rdata(f1908_rdata));
  assign f1908_clk = clk;
  assign f1908_rst = rst;
  // Bindings to f1908

  // f1910
  logic [0:0] f1910_wen;
  logic [31:0] f1910_wdata;
  logic [0:0] f1910_clk;
  logic [0:0] f1910_rst;
  logic [31:0] f1910_rdata;
  sr_buffer_32_1 f1910(.wen(f1910_wen), .wdata(f1910_wdata), .clk(f1910_clk), .rst(f1910_rst), .rdata(f1910_rdata));
  assign f1910_clk = clk;
  assign f1910_rst = rst;
  // Bindings to f1910

  // f1912
  logic [0:0] f1912_wen;
  logic [31:0] f1912_wdata;
  logic [0:0] f1912_clk;
  logic [0:0] f1912_rst;
  logic [31:0] f1912_rdata;
  sr_buffer_32_1 f1912(.wen(f1912_wen), .wdata(f1912_wdata), .clk(f1912_clk), .rst(f1912_rst), .rdata(f1912_rdata));
  assign f1912_clk = clk;
  assign f1912_rst = rst;
  // Bindings to f1912

  // f1914
  logic [0:0] f1914_wen;
  logic [31:0] f1914_wdata;
  logic [0:0] f1914_clk;
  logic [0:0] f1914_rst;
  logic [31:0] f1914_rdata;
  sr_buffer_32_1 f1914(.wen(f1914_wen), .wdata(f1914_wdata), .clk(f1914_clk), .rst(f1914_rst), .rdata(f1914_rdata));
  assign f1914_clk = clk;
  assign f1914_rst = rst;
  // Bindings to f1914

  // f1916
  logic [0:0] f1916_wen;
  logic [31:0] f1916_wdata;
  logic [0:0] f1916_clk;
  logic [0:0] f1916_rst;
  logic [31:0] f1916_rdata;
  sr_buffer_32_1 f1916(.wen(f1916_wen), .wdata(f1916_wdata), .clk(f1916_clk), .rst(f1916_rst), .rdata(f1916_rdata));
  assign f1916_clk = clk;
  assign f1916_rst = rst;
  // Bindings to f1916

  // f1918
  logic [0:0] f1918_wen;
  logic [31:0] f1918_wdata;
  logic [0:0] f1918_clk;
  logic [0:0] f1918_rst;
  logic [31:0] f1918_rdata;
  sr_buffer_32_1 f1918(.wen(f1918_wen), .wdata(f1918_wdata), .clk(f1918_clk), .rst(f1918_rst), .rdata(f1918_rdata));
  assign f1918_clk = clk;
  assign f1918_rst = rst;
  // Bindings to f1918

  // f1920
  logic [0:0] f1920_wen;
  logic [31:0] f1920_wdata;
  logic [0:0] f1920_clk;
  logic [0:0] f1920_rst;
  logic [31:0] f1920_rdata;
  sr_buffer_32_1 f1920(.wen(f1920_wen), .wdata(f1920_wdata), .clk(f1920_clk), .rst(f1920_rst), .rdata(f1920_rdata));
  assign f1920_clk = clk;
  assign f1920_rst = rst;
  // Bindings to f1920

  // f1922
  logic [0:0] f1922_wen;
  logic [31:0] f1922_wdata;
  logic [0:0] f1922_clk;
  logic [0:0] f1922_rst;
  logic [31:0] f1922_rdata;
  sr_buffer_32_1 f1922(.wen(f1922_wen), .wdata(f1922_wdata), .clk(f1922_clk), .rst(f1922_rst), .rdata(f1922_rdata));
  assign f1922_clk = clk;
  assign f1922_rst = rst;
  // Bindings to f1922

  // f1924
  logic [0:0] f1924_wen;
  logic [31:0] f1924_wdata;
  logic [0:0] f1924_clk;
  logic [0:0] f1924_rst;
  logic [31:0] f1924_rdata;
  sr_buffer_32_1 f1924(.wen(f1924_wen), .wdata(f1924_wdata), .clk(f1924_clk), .rst(f1924_rst), .rdata(f1924_rdata));
  assign f1924_clk = clk;
  assign f1924_rst = rst;
  // Bindings to f1924

  // f1926
  logic [0:0] f1926_wen;
  logic [31:0] f1926_wdata;
  logic [0:0] f1926_clk;
  logic [0:0] f1926_rst;
  logic [31:0] f1926_rdata;
  sr_buffer_32_1 f1926(.wen(f1926_wen), .wdata(f1926_wdata), .clk(f1926_clk), .rst(f1926_rst), .rdata(f1926_rdata));
  assign f1926_clk = clk;
  assign f1926_rst = rst;
  // Bindings to f1926

  // f1928
  logic [0:0] f1928_wen;
  logic [31:0] f1928_wdata;
  logic [0:0] f1928_clk;
  logic [0:0] f1928_rst;
  logic [31:0] f1928_rdata;
  sr_buffer_32_1 f1928(.wen(f1928_wen), .wdata(f1928_wdata), .clk(f1928_clk), .rst(f1928_rst), .rdata(f1928_rdata));
  assign f1928_clk = clk;
  assign f1928_rst = rst;
  // Bindings to f1928

  // f1930
  logic [0:0] f1930_wen;
  logic [31:0] f1930_wdata;
  logic [0:0] f1930_clk;
  logic [0:0] f1930_rst;
  logic [31:0] f1930_rdata;
  sr_buffer_32_1 f1930(.wen(f1930_wen), .wdata(f1930_wdata), .clk(f1930_clk), .rst(f1930_rst), .rdata(f1930_rdata));
  assign f1930_clk = clk;
  assign f1930_rst = rst;
  // Bindings to f1930

  // f1932
  logic [0:0] f1932_wen;
  logic [31:0] f1932_wdata;
  logic [0:0] f1932_clk;
  logic [0:0] f1932_rst;
  logic [31:0] f1932_rdata;
  sr_buffer_32_1 f1932(.wen(f1932_wen), .wdata(f1932_wdata), .clk(f1932_clk), .rst(f1932_rst), .rdata(f1932_rdata));
  assign f1932_clk = clk;
  assign f1932_rst = rst;
  // Bindings to f1932

  // f1934
  logic [0:0] f1934_wen;
  logic [31:0] f1934_wdata;
  logic [0:0] f1934_clk;
  logic [0:0] f1934_rst;
  logic [31:0] f1934_rdata;
  sr_buffer_32_1 f1934(.wen(f1934_wen), .wdata(f1934_wdata), .clk(f1934_clk), .rst(f1934_rst), .rdata(f1934_rdata));
  assign f1934_clk = clk;
  assign f1934_rst = rst;
  // Bindings to f1934

  // f1936
  logic [0:0] f1936_wen;
  logic [31:0] f1936_wdata;
  logic [0:0] f1936_clk;
  logic [0:0] f1936_rst;
  logic [31:0] f1936_rdata;
  sr_buffer_32_1 f1936(.wen(f1936_wen), .wdata(f1936_wdata), .clk(f1936_clk), .rst(f1936_rst), .rdata(f1936_rdata));
  assign f1936_clk = clk;
  assign f1936_rst = rst;
  // Bindings to f1936

  // f1938
  logic [0:0] f1938_wen;
  logic [31:0] f1938_wdata;
  logic [0:0] f1938_clk;
  logic [0:0] f1938_rst;
  logic [31:0] f1938_rdata;
  sr_buffer_32_1 f1938(.wen(f1938_wen), .wdata(f1938_wdata), .clk(f1938_clk), .rst(f1938_rst), .rdata(f1938_rdata));
  assign f1938_clk = clk;
  assign f1938_rst = rst;
  // Bindings to f1938

  // f1940
  logic [0:0] f1940_wen;
  logic [31:0] f1940_wdata;
  logic [0:0] f1940_clk;
  logic [0:0] f1940_rst;
  logic [31:0] f1940_rdata;
  sr_buffer_32_1 f1940(.wen(f1940_wen), .wdata(f1940_wdata), .clk(f1940_clk), .rst(f1940_rst), .rdata(f1940_rdata));
  assign f1940_clk = clk;
  assign f1940_rst = rst;
  // Bindings to f1940

  // f1942
  logic [0:0] f1942_wen;
  logic [31:0] f1942_wdata;
  logic [0:0] f1942_clk;
  logic [0:0] f1942_rst;
  logic [31:0] f1942_rdata;
  sr_buffer_32_1 f1942(.wen(f1942_wen), .wdata(f1942_wdata), .clk(f1942_clk), .rst(f1942_rst), .rdata(f1942_rdata));
  assign f1942_clk = clk;
  assign f1942_rst = rst;
  // Bindings to f1942

  // f1944
  logic [0:0] f1944_wen;
  logic [31:0] f1944_wdata;
  logic [0:0] f1944_clk;
  logic [0:0] f1944_rst;
  logic [31:0] f1944_rdata;
  sr_buffer_32_1 f1944(.wen(f1944_wen), .wdata(f1944_wdata), .clk(f1944_clk), .rst(f1944_rst), .rdata(f1944_rdata));
  assign f1944_clk = clk;
  assign f1944_rst = rst;
  // Bindings to f1944

  // f1946
  logic [0:0] f1946_wen;
  logic [31:0] f1946_wdata;
  logic [0:0] f1946_clk;
  logic [0:0] f1946_rst;
  logic [31:0] f1946_rdata;
  sr_buffer_32_1 f1946(.wen(f1946_wen), .wdata(f1946_wdata), .clk(f1946_clk), .rst(f1946_rst), .rdata(f1946_rdata));
  assign f1946_clk = clk;
  assign f1946_rst = rst;
  // Bindings to f1946

  // f1948
  logic [0:0] f1948_wen;
  logic [31:0] f1948_wdata;
  logic [0:0] f1948_clk;
  logic [0:0] f1948_rst;
  logic [31:0] f1948_rdata;
  sr_buffer_32_1 f1948(.wen(f1948_wen), .wdata(f1948_wdata), .clk(f1948_clk), .rst(f1948_rst), .rdata(f1948_rdata));
  assign f1948_clk = clk;
  assign f1948_rst = rst;
  // Bindings to f1948

  // f1950
  logic [0:0] f1950_wen;
  logic [31:0] f1950_wdata;
  logic [0:0] f1950_clk;
  logic [0:0] f1950_rst;
  logic [31:0] f1950_rdata;
  sr_buffer_32_1 f1950(.wen(f1950_wen), .wdata(f1950_wdata), .clk(f1950_clk), .rst(f1950_rst), .rdata(f1950_rdata));
  assign f1950_clk = clk;
  assign f1950_rst = rst;
  // Bindings to f1950

  // f1952
  logic [0:0] f1952_wen;
  logic [31:0] f1952_wdata;
  logic [0:0] f1952_clk;
  logic [0:0] f1952_rst;
  logic [31:0] f1952_rdata;
  sr_buffer_32_1 f1952(.wen(f1952_wen), .wdata(f1952_wdata), .clk(f1952_clk), .rst(f1952_rst), .rdata(f1952_rdata));
  assign f1952_clk = clk;
  assign f1952_rst = rst;
  // Bindings to f1952

  // f1954
  logic [0:0] f1954_wen;
  logic [31:0] f1954_wdata;
  logic [0:0] f1954_clk;
  logic [0:0] f1954_rst;
  logic [31:0] f1954_rdata;
  sr_buffer_32_1 f1954(.wen(f1954_wen), .wdata(f1954_wdata), .clk(f1954_clk), .rst(f1954_rst), .rdata(f1954_rdata));
  assign f1954_clk = clk;
  assign f1954_rst = rst;
  // Bindings to f1954

  // f1956
  logic [0:0] f1956_wen;
  logic [31:0] f1956_wdata;
  logic [0:0] f1956_clk;
  logic [0:0] f1956_rst;
  logic [31:0] f1956_rdata;
  sr_buffer_32_1 f1956(.wen(f1956_wen), .wdata(f1956_wdata), .clk(f1956_clk), .rst(f1956_rst), .rdata(f1956_rdata));
  assign f1956_clk = clk;
  assign f1956_rst = rst;
  // Bindings to f1956

  // f1958
  logic [0:0] f1958_wen;
  logic [31:0] f1958_wdata;
  logic [0:0] f1958_clk;
  logic [0:0] f1958_rst;
  logic [31:0] f1958_rdata;
  sr_buffer_32_1 f1958(.wen(f1958_wen), .wdata(f1958_wdata), .clk(f1958_clk), .rst(f1958_rst), .rdata(f1958_rdata));
  assign f1958_clk = clk;
  assign f1958_rst = rst;
  // Bindings to f1958

  // f1960
  logic [0:0] f1960_wen;
  logic [31:0] f1960_wdata;
  logic [0:0] f1960_clk;
  logic [0:0] f1960_rst;
  logic [31:0] f1960_rdata;
  sr_buffer_32_1 f1960(.wen(f1960_wen), .wdata(f1960_wdata), .clk(f1960_clk), .rst(f1960_rst), .rdata(f1960_rdata));
  assign f1960_clk = clk;
  assign f1960_rst = rst;
  // Bindings to f1960

  // f1962
  logic [0:0] f1962_wen;
  logic [31:0] f1962_wdata;
  logic [0:0] f1962_clk;
  logic [0:0] f1962_rst;
  logic [31:0] f1962_rdata;
  sr_buffer_32_1 f1962(.wen(f1962_wen), .wdata(f1962_wdata), .clk(f1962_clk), .rst(f1962_rst), .rdata(f1962_rdata));
  assign f1962_clk = clk;
  assign f1962_rst = rst;
  // Bindings to f1962

  // f1964
  logic [0:0] f1964_wen;
  logic [31:0] f1964_wdata;
  logic [0:0] f1964_clk;
  logic [0:0] f1964_rst;
  logic [31:0] f1964_rdata;
  sr_buffer_32_1 f1964(.wen(f1964_wen), .wdata(f1964_wdata), .clk(f1964_clk), .rst(f1964_rst), .rdata(f1964_rdata));
  assign f1964_clk = clk;
  assign f1964_rst = rst;
  // Bindings to f1964

  // f1966
  logic [0:0] f1966_wen;
  logic [31:0] f1966_wdata;
  logic [0:0] f1966_clk;
  logic [0:0] f1966_rst;
  logic [31:0] f1966_rdata;
  sr_buffer_32_1 f1966(.wen(f1966_wen), .wdata(f1966_wdata), .clk(f1966_clk), .rst(f1966_rst), .rdata(f1966_rdata));
  assign f1966_clk = clk;
  assign f1966_rst = rst;
  // Bindings to f1966

  // f1968
  logic [0:0] f1968_wen;
  logic [31:0] f1968_wdata;
  logic [0:0] f1968_clk;
  logic [0:0] f1968_rst;
  logic [31:0] f1968_rdata;
  sr_buffer_32_1 f1968(.wen(f1968_wen), .wdata(f1968_wdata), .clk(f1968_clk), .rst(f1968_rst), .rdata(f1968_rdata));
  assign f1968_clk = clk;
  assign f1968_rst = rst;
  // Bindings to f1968

  // f1970
  logic [0:0] f1970_wen;
  logic [31:0] f1970_wdata;
  logic [0:0] f1970_clk;
  logic [0:0] f1970_rst;
  logic [31:0] f1970_rdata;
  sr_buffer_32_1 f1970(.wen(f1970_wen), .wdata(f1970_wdata), .clk(f1970_clk), .rst(f1970_rst), .rdata(f1970_rdata));
  assign f1970_clk = clk;
  assign f1970_rst = rst;
  // Bindings to f1970

  // f1972
  logic [0:0] f1972_wen;
  logic [31:0] f1972_wdata;
  logic [0:0] f1972_clk;
  logic [0:0] f1972_rst;
  logic [31:0] f1972_rdata;
  sr_buffer_32_1 f1972(.wen(f1972_wen), .wdata(f1972_wdata), .clk(f1972_clk), .rst(f1972_rst), .rdata(f1972_rdata));
  assign f1972_clk = clk;
  assign f1972_rst = rst;
  // Bindings to f1972

  // f1974
  logic [0:0] f1974_wen;
  logic [31:0] f1974_wdata;
  logic [0:0] f1974_clk;
  logic [0:0] f1974_rst;
  logic [31:0] f1974_rdata;
  sr_buffer_32_1 f1974(.wen(f1974_wen), .wdata(f1974_wdata), .clk(f1974_clk), .rst(f1974_rst), .rdata(f1974_rdata));
  assign f1974_clk = clk;
  assign f1974_rst = rst;
  // Bindings to f1974

  // f1976
  logic [0:0] f1976_wen;
  logic [31:0] f1976_wdata;
  logic [0:0] f1976_clk;
  logic [0:0] f1976_rst;
  logic [31:0] f1976_rdata;
  sr_buffer_32_1 f1976(.wen(f1976_wen), .wdata(f1976_wdata), .clk(f1976_clk), .rst(f1976_rst), .rdata(f1976_rdata));
  assign f1976_clk = clk;
  assign f1976_rst = rst;
  // Bindings to f1976

  // f1978
  logic [0:0] f1978_wen;
  logic [31:0] f1978_wdata;
  logic [0:0] f1978_clk;
  logic [0:0] f1978_rst;
  logic [31:0] f1978_rdata;
  sr_buffer_32_1 f1978(.wen(f1978_wen), .wdata(f1978_wdata), .clk(f1978_clk), .rst(f1978_rst), .rdata(f1978_rdata));
  assign f1978_clk = clk;
  assign f1978_rst = rst;
  // Bindings to f1978

  // f1980
  logic [0:0] f1980_wen;
  logic [31:0] f1980_wdata;
  logic [0:0] f1980_clk;
  logic [0:0] f1980_rst;
  logic [31:0] f1980_rdata;
  sr_buffer_32_1 f1980(.wen(f1980_wen), .wdata(f1980_wdata), .clk(f1980_clk), .rst(f1980_rst), .rdata(f1980_rdata));
  assign f1980_clk = clk;
  assign f1980_rst = rst;
  // Bindings to f1980

  // f1982
  logic [0:0] f1982_wen;
  logic [31:0] f1982_wdata;
  logic [0:0] f1982_clk;
  logic [0:0] f1982_rst;
  logic [31:0] f1982_rdata;
  sr_buffer_32_1 f1982(.wen(f1982_wen), .wdata(f1982_wdata), .clk(f1982_clk), .rst(f1982_rst), .rdata(f1982_rdata));
  assign f1982_clk = clk;
  assign f1982_rst = rst;
  // Bindings to f1982

  // f1984
  logic [0:0] f1984_wen;
  logic [31:0] f1984_wdata;
  logic [0:0] f1984_clk;
  logic [0:0] f1984_rst;
  logic [31:0] f1984_rdata;
  sr_buffer_32_1 f1984(.wen(f1984_wen), .wdata(f1984_wdata), .clk(f1984_clk), .rst(f1984_rst), .rdata(f1984_rdata));
  assign f1984_clk = clk;
  assign f1984_rst = rst;
  // Bindings to f1984

  // f1986
  logic [0:0] f1986_wen;
  logic [31:0] f1986_wdata;
  logic [0:0] f1986_clk;
  logic [0:0] f1986_rst;
  logic [31:0] f1986_rdata;
  sr_buffer_32_1 f1986(.wen(f1986_wen), .wdata(f1986_wdata), .clk(f1986_clk), .rst(f1986_rst), .rdata(f1986_rdata));
  assign f1986_clk = clk;
  assign f1986_rst = rst;
  // Bindings to f1986

  // f1988
  logic [0:0] f1988_wen;
  logic [31:0] f1988_wdata;
  logic [0:0] f1988_clk;
  logic [0:0] f1988_rst;
  logic [31:0] f1988_rdata;
  sr_buffer_32_1 f1988(.wen(f1988_wen), .wdata(f1988_wdata), .clk(f1988_clk), .rst(f1988_rst), .rdata(f1988_rdata));
  assign f1988_clk = clk;
  assign f1988_rst = rst;
  // Bindings to f1988

  // f1990
  logic [0:0] f1990_wen;
  logic [31:0] f1990_wdata;
  logic [0:0] f1990_clk;
  logic [0:0] f1990_rst;
  logic [31:0] f1990_rdata;
  sr_buffer_32_1 f1990(.wen(f1990_wen), .wdata(f1990_wdata), .clk(f1990_clk), .rst(f1990_rst), .rdata(f1990_rdata));
  assign f1990_clk = clk;
  assign f1990_rst = rst;
  // Bindings to f1990

  // f1992
  logic [0:0] f1992_wen;
  logic [31:0] f1992_wdata;
  logic [0:0] f1992_clk;
  logic [0:0] f1992_rst;
  logic [31:0] f1992_rdata;
  sr_buffer_32_1 f1992(.wen(f1992_wen), .wdata(f1992_wdata), .clk(f1992_clk), .rst(f1992_rst), .rdata(f1992_rdata));
  assign f1992_clk = clk;
  assign f1992_rst = rst;
  // Bindings to f1992

  // f1994
  logic [0:0] f1994_wen;
  logic [31:0] f1994_wdata;
  logic [0:0] f1994_clk;
  logic [0:0] f1994_rst;
  logic [31:0] f1994_rdata;
  sr_buffer_32_1 f1994(.wen(f1994_wen), .wdata(f1994_wdata), .clk(f1994_clk), .rst(f1994_rst), .rdata(f1994_rdata));
  assign f1994_clk = clk;
  assign f1994_rst = rst;
  // Bindings to f1994

  // f1996
  logic [0:0] f1996_wen;
  logic [31:0] f1996_wdata;
  logic [0:0] f1996_clk;
  logic [0:0] f1996_rst;
  logic [31:0] f1996_rdata;
  sr_buffer_32_1 f1996(.wen(f1996_wen), .wdata(f1996_wdata), .clk(f1996_clk), .rst(f1996_rst), .rdata(f1996_rdata));
  assign f1996_clk = clk;
  assign f1996_rst = rst;
  // Bindings to f1996

  // f1998
  logic [0:0] f1998_wen;
  logic [31:0] f1998_wdata;
  logic [0:0] f1998_clk;
  logic [0:0] f1998_rst;
  logic [31:0] f1998_rdata;
  sr_buffer_32_1 f1998(.wen(f1998_wen), .wdata(f1998_wdata), .clk(f1998_clk), .rst(f1998_rst), .rdata(f1998_rdata));
  assign f1998_clk = clk;
  assign f1998_rst = rst;
  // Bindings to f1998

  // f2000
  logic [0:0] f2000_wen;
  logic [31:0] f2000_wdata;
  logic [0:0] f2000_clk;
  logic [0:0] f2000_rst;
  logic [31:0] f2000_rdata;
  sr_buffer_32_1 f2000(.wen(f2000_wen), .wdata(f2000_wdata), .clk(f2000_clk), .rst(f2000_rst), .rdata(f2000_rdata));
  assign f2000_clk = clk;
  assign f2000_rst = rst;
  // Bindings to f2000

  // f2002
  logic [0:0] f2002_wen;
  logic [31:0] f2002_wdata;
  logic [0:0] f2002_clk;
  logic [0:0] f2002_rst;
  logic [31:0] f2002_rdata;
  sr_buffer_32_1 f2002(.wen(f2002_wen), .wdata(f2002_wdata), .clk(f2002_clk), .rst(f2002_rst), .rdata(f2002_rdata));
  assign f2002_clk = clk;
  assign f2002_rst = rst;
  // Bindings to f2002

  // f2004
  logic [0:0] f2004_wen;
  logic [31:0] f2004_wdata;
  logic [0:0] f2004_clk;
  logic [0:0] f2004_rst;
  logic [31:0] f2004_rdata;
  sr_buffer_32_1 f2004(.wen(f2004_wen), .wdata(f2004_wdata), .clk(f2004_clk), .rst(f2004_rst), .rdata(f2004_rdata));
  assign f2004_clk = clk;
  assign f2004_rst = rst;
  // Bindings to f2004

  // f2006
  logic [0:0] f2006_wen;
  logic [31:0] f2006_wdata;
  logic [0:0] f2006_clk;
  logic [0:0] f2006_rst;
  logic [31:0] f2006_rdata;
  sr_buffer_32_1 f2006(.wen(f2006_wen), .wdata(f2006_wdata), .clk(f2006_clk), .rst(f2006_rst), .rdata(f2006_rdata));
  assign f2006_clk = clk;
  assign f2006_rst = rst;
  // Bindings to f2006

  // f2008
  logic [0:0] f2008_wen;
  logic [31:0] f2008_wdata;
  logic [0:0] f2008_clk;
  logic [0:0] f2008_rst;
  logic [31:0] f2008_rdata;
  sr_buffer_32_1 f2008(.wen(f2008_wen), .wdata(f2008_wdata), .clk(f2008_clk), .rst(f2008_rst), .rdata(f2008_rdata));
  assign f2008_clk = clk;
  assign f2008_rst = rst;
  // Bindings to f2008

  // f2010
  logic [0:0] f2010_wen;
  logic [31:0] f2010_wdata;
  logic [0:0] f2010_clk;
  logic [0:0] f2010_rst;
  logic [31:0] f2010_rdata;
  sr_buffer_32_1 f2010(.wen(f2010_wen), .wdata(f2010_wdata), .clk(f2010_clk), .rst(f2010_rst), .rdata(f2010_rdata));
  assign f2010_clk = clk;
  assign f2010_rst = rst;
  // Bindings to f2010

  // f2012
  logic [0:0] f2012_wen;
  logic [31:0] f2012_wdata;
  logic [0:0] f2012_clk;
  logic [0:0] f2012_rst;
  logic [31:0] f2012_rdata;
  sr_buffer_32_1 f2012(.wen(f2012_wen), .wdata(f2012_wdata), .clk(f2012_clk), .rst(f2012_rst), .rdata(f2012_rdata));
  assign f2012_clk = clk;
  assign f2012_rst = rst;
  // Bindings to f2012

  // f2014
  logic [0:0] f2014_wen;
  logic [31:0] f2014_wdata;
  logic [0:0] f2014_clk;
  logic [0:0] f2014_rst;
  logic [31:0] f2014_rdata;
  sr_buffer_32_1 f2014(.wen(f2014_wen), .wdata(f2014_wdata), .clk(f2014_clk), .rst(f2014_rst), .rdata(f2014_rdata));
  assign f2014_clk = clk;
  assign f2014_rst = rst;
  // Bindings to f2014

  // f2016
  logic [0:0] f2016_wen;
  logic [31:0] f2016_wdata;
  logic [0:0] f2016_clk;
  logic [0:0] f2016_rst;
  logic [31:0] f2016_rdata;
  sr_buffer_32_1 f2016(.wen(f2016_wen), .wdata(f2016_wdata), .clk(f2016_clk), .rst(f2016_rst), .rdata(f2016_rdata));
  assign f2016_clk = clk;
  assign f2016_rst = rst;
  // Bindings to f2016

  // f2018
  logic [0:0] f2018_wen;
  logic [31:0] f2018_wdata;
  logic [0:0] f2018_clk;
  logic [0:0] f2018_rst;
  logic [31:0] f2018_rdata;
  sr_buffer_32_1 f2018(.wen(f2018_wen), .wdata(f2018_wdata), .clk(f2018_clk), .rst(f2018_rst), .rdata(f2018_rdata));
  assign f2018_clk = clk;
  assign f2018_rst = rst;
  // Bindings to f2018

  // f2020
  logic [0:0] f2020_wen;
  logic [31:0] f2020_wdata;
  logic [0:0] f2020_clk;
  logic [0:0] f2020_rst;
  logic [31:0] f2020_rdata;
  sr_buffer_32_1 f2020(.wen(f2020_wen), .wdata(f2020_wdata), .clk(f2020_clk), .rst(f2020_rst), .rdata(f2020_rdata));
  assign f2020_clk = clk;
  assign f2020_rst = rst;
  // Bindings to f2020

  // f2022
  logic [0:0] f2022_wen;
  logic [31:0] f2022_wdata;
  logic [0:0] f2022_clk;
  logic [0:0] f2022_rst;
  logic [31:0] f2022_rdata;
  sr_buffer_32_1 f2022(.wen(f2022_wen), .wdata(f2022_wdata), .clk(f2022_clk), .rst(f2022_rst), .rdata(f2022_rdata));
  assign f2022_clk = clk;
  assign f2022_rst = rst;
  // Bindings to f2022

  // f2024
  logic [0:0] f2024_wen;
  logic [31:0] f2024_wdata;
  logic [0:0] f2024_clk;
  logic [0:0] f2024_rst;
  logic [31:0] f2024_rdata;
  sr_buffer_32_1 f2024(.wen(f2024_wen), .wdata(f2024_wdata), .clk(f2024_clk), .rst(f2024_rst), .rdata(f2024_rdata));
  assign f2024_clk = clk;
  assign f2024_rst = rst;
  // Bindings to f2024

  // f2026
  logic [0:0] f2026_wen;
  logic [31:0] f2026_wdata;
  logic [0:0] f2026_clk;
  logic [0:0] f2026_rst;
  logic [31:0] f2026_rdata;
  sr_buffer_32_1 f2026(.wen(f2026_wen), .wdata(f2026_wdata), .clk(f2026_clk), .rst(f2026_rst), .rdata(f2026_rdata));
  assign f2026_clk = clk;
  assign f2026_rst = rst;
  // Bindings to f2026

  // f2028
  logic [0:0] f2028_wen;
  logic [31:0] f2028_wdata;
  logic [0:0] f2028_clk;
  logic [0:0] f2028_rst;
  logic [31:0] f2028_rdata;
  sr_buffer_32_1 f2028(.wen(f2028_wen), .wdata(f2028_wdata), .clk(f2028_clk), .rst(f2028_rst), .rdata(f2028_rdata));
  assign f2028_clk = clk;
  assign f2028_rst = rst;
  // Bindings to f2028

  // f2030
  logic [0:0] f2030_wen;
  logic [31:0] f2030_wdata;
  logic [0:0] f2030_clk;
  logic [0:0] f2030_rst;
  logic [31:0] f2030_rdata;
  sr_buffer_32_1 f2030(.wen(f2030_wen), .wdata(f2030_wdata), .clk(f2030_clk), .rst(f2030_rst), .rdata(f2030_rdata));
  assign f2030_clk = clk;
  assign f2030_rst = rst;
  // Bindings to f2030

  // f2032
  logic [0:0] f2032_wen;
  logic [31:0] f2032_wdata;
  logic [0:0] f2032_clk;
  logic [0:0] f2032_rst;
  logic [31:0] f2032_rdata;
  sr_buffer_32_1 f2032(.wen(f2032_wen), .wdata(f2032_wdata), .clk(f2032_clk), .rst(f2032_rst), .rdata(f2032_rdata));
  assign f2032_clk = clk;
  assign f2032_rst = rst;
  // Bindings to f2032

  // f2034
  logic [0:0] f2034_wen;
  logic [31:0] f2034_wdata;
  logic [0:0] f2034_clk;
  logic [0:0] f2034_rst;
  logic [31:0] f2034_rdata;
  sr_buffer_32_1 f2034(.wen(f2034_wen), .wdata(f2034_wdata), .clk(f2034_clk), .rst(f2034_rst), .rdata(f2034_rdata));
  assign f2034_clk = clk;
  assign f2034_rst = rst;
  // Bindings to f2034

  // f2036
  logic [0:0] f2036_wen;
  logic [31:0] f2036_wdata;
  logic [0:0] f2036_clk;
  logic [0:0] f2036_rst;
  logic [31:0] f2036_rdata;
  sr_buffer_32_1 f2036(.wen(f2036_wen), .wdata(f2036_wdata), .clk(f2036_clk), .rst(f2036_rst), .rdata(f2036_rdata));
  assign f2036_clk = clk;
  assign f2036_rst = rst;
  // Bindings to f2036

  // f2038
  logic [0:0] f2038_wen;
  logic [31:0] f2038_wdata;
  logic [0:0] f2038_clk;
  logic [0:0] f2038_rst;
  logic [31:0] f2038_rdata;
  sr_buffer_32_1 f2038(.wen(f2038_wen), .wdata(f2038_wdata), .clk(f2038_clk), .rst(f2038_rst), .rdata(f2038_rdata));
  assign f2038_clk = clk;
  assign f2038_rst = rst;
  // Bindings to f2038

  // f2040
  logic [0:0] f2040_wen;
  logic [31:0] f2040_wdata;
  logic [0:0] f2040_clk;
  logic [0:0] f2040_rst;
  logic [31:0] f2040_rdata;
  sr_buffer_32_1 f2040(.wen(f2040_wen), .wdata(f2040_wdata), .clk(f2040_clk), .rst(f2040_rst), .rdata(f2040_rdata));
  assign f2040_clk = clk;
  assign f2040_rst = rst;
  // Bindings to f2040

  // f2042
  logic [0:0] f2042_wen;
  logic [31:0] f2042_wdata;
  logic [0:0] f2042_clk;
  logic [0:0] f2042_rst;
  logic [31:0] f2042_rdata;
  sr_buffer_32_1 f2042(.wen(f2042_wen), .wdata(f2042_wdata), .clk(f2042_clk), .rst(f2042_rst), .rdata(f2042_rdata));
  assign f2042_clk = clk;
  assign f2042_rst = rst;
  // Bindings to f2042

  // f2044
  logic [0:0] f2044_wen;
  logic [31:0] f2044_wdata;
  logic [0:0] f2044_clk;
  logic [0:0] f2044_rst;
  logic [31:0] f2044_rdata;
  sr_buffer_32_1 f2044(.wen(f2044_wen), .wdata(f2044_wdata), .clk(f2044_clk), .rst(f2044_rst), .rdata(f2044_rdata));
  assign f2044_clk = clk;
  assign f2044_rst = rst;
  // Bindings to f2044

  // f2046
  logic [0:0] f2046_wen;
  logic [31:0] f2046_wdata;
  logic [0:0] f2046_clk;
  logic [0:0] f2046_rst;
  logic [31:0] f2046_rdata;
  sr_buffer_32_1 f2046(.wen(f2046_wen), .wdata(f2046_wdata), .clk(f2046_clk), .rst(f2046_rst), .rdata(f2046_rdata));
  assign f2046_clk = clk;
  assign f2046_rst = rst;
  // Bindings to f2046

  // f2048
  logic [0:0] f2048_wen;
  logic [31:0] f2048_wdata;
  logic [0:0] f2048_clk;
  logic [0:0] f2048_rst;
  logic [31:0] f2048_rdata;
  sr_buffer_32_1 f2048(.wen(f2048_wen), .wdata(f2048_wdata), .clk(f2048_clk), .rst(f2048_rst), .rdata(f2048_rdata));
  assign f2048_clk = clk;
  assign f2048_rst = rst;
  // Bindings to f2048

  // f2050
  logic [0:0] f2050_wen;
  logic [31:0] f2050_wdata;
  logic [0:0] f2050_clk;
  logic [0:0] f2050_rst;
  logic [31:0] f2050_rdata;
  sr_buffer_32_1 f2050(.wen(f2050_wen), .wdata(f2050_wdata), .clk(f2050_clk), .rst(f2050_rst), .rdata(f2050_rdata));
  assign f2050_clk = clk;
  assign f2050_rst = rst;
  // Bindings to f2050

  // f2052
  logic [0:0] f2052_wen;
  logic [31:0] f2052_wdata;
  logic [0:0] f2052_clk;
  logic [0:0] f2052_rst;
  logic [31:0] f2052_rdata;
  sr_buffer_32_1 f2052(.wen(f2052_wen), .wdata(f2052_wdata), .clk(f2052_clk), .rst(f2052_rst), .rdata(f2052_rdata));
  assign f2052_clk = clk;
  assign f2052_rst = rst;
  // Bindings to f2052

  // f2054
  logic [0:0] f2054_wen;
  logic [31:0] f2054_wdata;
  logic [0:0] f2054_clk;
  logic [0:0] f2054_rst;
  logic [31:0] f2054_rdata;
  sr_buffer_32_1 f2054(.wen(f2054_wen), .wdata(f2054_wdata), .clk(f2054_clk), .rst(f2054_rst), .rdata(f2054_rdata));
  assign f2054_clk = clk;
  assign f2054_rst = rst;
  // Bindings to f2054

  // f2056
  logic [0:0] f2056_wen;
  logic [31:0] f2056_wdata;
  logic [0:0] f2056_clk;
  logic [0:0] f2056_rst;
  logic [31:0] f2056_rdata;
  sr_buffer_32_1 f2056(.wen(f2056_wen), .wdata(f2056_wdata), .clk(f2056_clk), .rst(f2056_rst), .rdata(f2056_rdata));
  assign f2056_clk = clk;
  assign f2056_rst = rst;
  // Bindings to f2056

  // f2058
  logic [0:0] f2058_wen;
  logic [31:0] f2058_wdata;
  logic [0:0] f2058_clk;
  logic [0:0] f2058_rst;
  logic [31:0] f2058_rdata;
  sr_buffer_32_1 f2058(.wen(f2058_wen), .wdata(f2058_wdata), .clk(f2058_clk), .rst(f2058_rst), .rdata(f2058_rdata));
  assign f2058_clk = clk;
  assign f2058_rst = rst;
  // Bindings to f2058

  // f2060
  logic [0:0] f2060_wen;
  logic [31:0] f2060_wdata;
  logic [0:0] f2060_clk;
  logic [0:0] f2060_rst;
  logic [31:0] f2060_rdata;
  sr_buffer_32_1 f2060(.wen(f2060_wen), .wdata(f2060_wdata), .clk(f2060_clk), .rst(f2060_rst), .rdata(f2060_rdata));
  assign f2060_clk = clk;
  assign f2060_rst = rst;
  // Bindings to f2060

  // f2062
  logic [0:0] f2062_wen;
  logic [31:0] f2062_wdata;
  logic [0:0] f2062_clk;
  logic [0:0] f2062_rst;
  logic [31:0] f2062_rdata;
  sr_buffer_32_1 f2062(.wen(f2062_wen), .wdata(f2062_wdata), .clk(f2062_clk), .rst(f2062_rst), .rdata(f2062_rdata));
  assign f2062_clk = clk;
  assign f2062_rst = rst;
  // Bindings to f2062

  // f2064
  logic [0:0] f2064_wen;
  logic [31:0] f2064_wdata;
  logic [0:0] f2064_clk;
  logic [0:0] f2064_rst;
  logic [31:0] f2064_rdata;
  sr_buffer_32_1 f2064(.wen(f2064_wen), .wdata(f2064_wdata), .clk(f2064_clk), .rst(f2064_rst), .rdata(f2064_rdata));
  assign f2064_clk = clk;
  assign f2064_rst = rst;
  // Bindings to f2064

  // f2066
  logic [0:0] f2066_wen;
  logic [31:0] f2066_wdata;
  logic [0:0] f2066_clk;
  logic [0:0] f2066_rst;
  logic [31:0] f2066_rdata;
  sr_buffer_32_1 f2066(.wen(f2066_wen), .wdata(f2066_wdata), .clk(f2066_clk), .rst(f2066_rst), .rdata(f2066_rdata));
  assign f2066_clk = clk;
  assign f2066_rst = rst;
  // Bindings to f2066

  // f2068
  logic [0:0] f2068_wen;
  logic [31:0] f2068_wdata;
  logic [0:0] f2068_clk;
  logic [0:0] f2068_rst;
  logic [31:0] f2068_rdata;
  sr_buffer_32_1 f2068(.wen(f2068_wen), .wdata(f2068_wdata), .clk(f2068_clk), .rst(f2068_rst), .rdata(f2068_rdata));
  assign f2068_clk = clk;
  assign f2068_rst = rst;
  // Bindings to f2068

  // f2070
  logic [0:0] f2070_wen;
  logic [31:0] f2070_wdata;
  logic [0:0] f2070_clk;
  logic [0:0] f2070_rst;
  logic [31:0] f2070_rdata;
  sr_buffer_32_1 f2070(.wen(f2070_wen), .wdata(f2070_wdata), .clk(f2070_clk), .rst(f2070_rst), .rdata(f2070_rdata));
  assign f2070_clk = clk;
  assign f2070_rst = rst;
  // Bindings to f2070

  // f2072
  logic [0:0] f2072_wen;
  logic [31:0] f2072_wdata;
  logic [0:0] f2072_clk;
  logic [0:0] f2072_rst;
  logic [31:0] f2072_rdata;
  sr_buffer_32_1 f2072(.wen(f2072_wen), .wdata(f2072_wdata), .clk(f2072_clk), .rst(f2072_rst), .rdata(f2072_rdata));
  assign f2072_clk = clk;
  assign f2072_rst = rst;
  // Bindings to f2072

  // f2074
  logic [0:0] f2074_wen;
  logic [31:0] f2074_wdata;
  logic [0:0] f2074_clk;
  logic [0:0] f2074_rst;
  logic [31:0] f2074_rdata;
  sr_buffer_32_1 f2074(.wen(f2074_wen), .wdata(f2074_wdata), .clk(f2074_clk), .rst(f2074_rst), .rdata(f2074_rdata));
  assign f2074_clk = clk;
  assign f2074_rst = rst;
  // Bindings to f2074

  // f2076
  logic [0:0] f2076_wen;
  logic [31:0] f2076_wdata;
  logic [0:0] f2076_clk;
  logic [0:0] f2076_rst;
  logic [31:0] f2076_rdata;
  sr_buffer_32_1 f2076(.wen(f2076_wen), .wdata(f2076_wdata), .clk(f2076_clk), .rst(f2076_rst), .rdata(f2076_rdata));
  assign f2076_clk = clk;
  assign f2076_rst = rst;
  // Bindings to f2076

  // f2078
  logic [0:0] f2078_wen;
  logic [31:0] f2078_wdata;
  logic [0:0] f2078_clk;
  logic [0:0] f2078_rst;
  logic [31:0] f2078_rdata;
  sr_buffer_32_1 f2078(.wen(f2078_wen), .wdata(f2078_wdata), .clk(f2078_clk), .rst(f2078_rst), .rdata(f2078_rdata));
  assign f2078_clk = clk;
  assign f2078_rst = rst;
  // Bindings to f2078

  // f2080
  logic [0:0] f2080_wen;
  logic [31:0] f2080_wdata;
  logic [0:0] f2080_clk;
  logic [0:0] f2080_rst;
  logic [31:0] f2080_rdata;
  sr_buffer_32_1 f2080(.wen(f2080_wen), .wdata(f2080_wdata), .clk(f2080_clk), .rst(f2080_rst), .rdata(f2080_rdata));
  assign f2080_clk = clk;
  assign f2080_rst = rst;
  // Bindings to f2080

  // f2082
  logic [0:0] f2082_wen;
  logic [31:0] f2082_wdata;
  logic [0:0] f2082_clk;
  logic [0:0] f2082_rst;
  logic [31:0] f2082_rdata;
  sr_buffer_32_1 f2082(.wen(f2082_wen), .wdata(f2082_wdata), .clk(f2082_clk), .rst(f2082_rst), .rdata(f2082_rdata));
  assign f2082_clk = clk;
  assign f2082_rst = rst;
  // Bindings to f2082

  // f2084
  logic [0:0] f2084_wen;
  logic [31:0] f2084_wdata;
  logic [0:0] f2084_clk;
  logic [0:0] f2084_rst;
  logic [31:0] f2084_rdata;
  sr_buffer_32_1 f2084(.wen(f2084_wen), .wdata(f2084_wdata), .clk(f2084_clk), .rst(f2084_rst), .rdata(f2084_rdata));
  assign f2084_clk = clk;
  assign f2084_rst = rst;
  // Bindings to f2084

  // f2086
  logic [0:0] f2086_wen;
  logic [31:0] f2086_wdata;
  logic [0:0] f2086_clk;
  logic [0:0] f2086_rst;
  logic [31:0] f2086_rdata;
  sr_buffer_32_1 f2086(.wen(f2086_wen), .wdata(f2086_wdata), .clk(f2086_clk), .rst(f2086_rst), .rdata(f2086_rdata));
  assign f2086_clk = clk;
  assign f2086_rst = rst;
  // Bindings to f2086

  // f2088
  logic [0:0] f2088_wen;
  logic [31:0] f2088_wdata;
  logic [0:0] f2088_clk;
  logic [0:0] f2088_rst;
  logic [31:0] f2088_rdata;
  sr_buffer_32_1 f2088(.wen(f2088_wen), .wdata(f2088_wdata), .clk(f2088_clk), .rst(f2088_rst), .rdata(f2088_rdata));
  assign f2088_clk = clk;
  assign f2088_rst = rst;
  // Bindings to f2088

  // f2090
  logic [0:0] f2090_wen;
  logic [31:0] f2090_wdata;
  logic [0:0] f2090_clk;
  logic [0:0] f2090_rst;
  logic [31:0] f2090_rdata;
  sr_buffer_32_1 f2090(.wen(f2090_wen), .wdata(f2090_wdata), .clk(f2090_clk), .rst(f2090_rst), .rdata(f2090_rdata));
  assign f2090_clk = clk;
  assign f2090_rst = rst;
  // Bindings to f2090

  // f2092
  logic [0:0] f2092_wen;
  logic [31:0] f2092_wdata;
  logic [0:0] f2092_clk;
  logic [0:0] f2092_rst;
  logic [31:0] f2092_rdata;
  sr_buffer_32_1 f2092(.wen(f2092_wen), .wdata(f2092_wdata), .clk(f2092_clk), .rst(f2092_rst), .rdata(f2092_rdata));
  assign f2092_clk = clk;
  assign f2092_rst = rst;
  // Bindings to f2092

  // f2094
  logic [0:0] f2094_wen;
  logic [31:0] f2094_wdata;
  logic [0:0] f2094_clk;
  logic [0:0] f2094_rst;
  logic [31:0] f2094_rdata;
  sr_buffer_32_1 f2094(.wen(f2094_wen), .wdata(f2094_wdata), .clk(f2094_clk), .rst(f2094_rst), .rdata(f2094_rdata));
  assign f2094_clk = clk;
  assign f2094_rst = rst;
  // Bindings to f2094

  // f2096
  logic [0:0] f2096_wen;
  logic [31:0] f2096_wdata;
  logic [0:0] f2096_clk;
  logic [0:0] f2096_rst;
  logic [31:0] f2096_rdata;
  sr_buffer_32_1 f2096(.wen(f2096_wen), .wdata(f2096_wdata), .clk(f2096_clk), .rst(f2096_rst), .rdata(f2096_rdata));
  assign f2096_clk = clk;
  assign f2096_rst = rst;
  // Bindings to f2096

  // f2098
  logic [0:0] f2098_wen;
  logic [31:0] f2098_wdata;
  logic [0:0] f2098_clk;
  logic [0:0] f2098_rst;
  logic [31:0] f2098_rdata;
  sr_buffer_32_1 f2098(.wen(f2098_wen), .wdata(f2098_wdata), .clk(f2098_clk), .rst(f2098_rst), .rdata(f2098_rdata));
  assign f2098_clk = clk;
  assign f2098_rst = rst;
  // Bindings to f2098

  // f2100
  logic [0:0] f2100_wen;
  logic [31:0] f2100_wdata;
  logic [0:0] f2100_clk;
  logic [0:0] f2100_rst;
  logic [31:0] f2100_rdata;
  sr_buffer_32_1 f2100(.wen(f2100_wen), .wdata(f2100_wdata), .clk(f2100_clk), .rst(f2100_rst), .rdata(f2100_rdata));
  assign f2100_clk = clk;
  assign f2100_rst = rst;
  // Bindings to f2100

  // f2102
  logic [0:0] f2102_wen;
  logic [31:0] f2102_wdata;
  logic [0:0] f2102_clk;
  logic [0:0] f2102_rst;
  logic [31:0] f2102_rdata;
  sr_buffer_32_1 f2102(.wen(f2102_wen), .wdata(f2102_wdata), .clk(f2102_clk), .rst(f2102_rst), .rdata(f2102_rdata));
  assign f2102_clk = clk;
  assign f2102_rst = rst;
  // Bindings to f2102

  // f2104
  logic [0:0] f2104_wen;
  logic [31:0] f2104_wdata;
  logic [0:0] f2104_clk;
  logic [0:0] f2104_rst;
  logic [31:0] f2104_rdata;
  sr_buffer_32_1 f2104(.wen(f2104_wen), .wdata(f2104_wdata), .clk(f2104_clk), .rst(f2104_rst), .rdata(f2104_rdata));
  assign f2104_clk = clk;
  assign f2104_rst = rst;
  // Bindings to f2104

  // f2106
  logic [0:0] f2106_wen;
  logic [31:0] f2106_wdata;
  logic [0:0] f2106_clk;
  logic [0:0] f2106_rst;
  logic [31:0] f2106_rdata;
  sr_buffer_32_1 f2106(.wen(f2106_wen), .wdata(f2106_wdata), .clk(f2106_clk), .rst(f2106_rst), .rdata(f2106_rdata));
  assign f2106_clk = clk;
  assign f2106_rst = rst;
  // Bindings to f2106

  // f2108
  logic [0:0] f2108_wen;
  logic [31:0] f2108_wdata;
  logic [0:0] f2108_clk;
  logic [0:0] f2108_rst;
  logic [31:0] f2108_rdata;
  sr_buffer_32_1 f2108(.wen(f2108_wen), .wdata(f2108_wdata), .clk(f2108_clk), .rst(f2108_rst), .rdata(f2108_rdata));
  assign f2108_clk = clk;
  assign f2108_rst = rst;
  // Bindings to f2108

  // f2110
  logic [0:0] f2110_wen;
  logic [31:0] f2110_wdata;
  logic [0:0] f2110_clk;
  logic [0:0] f2110_rst;
  logic [31:0] f2110_rdata;
  sr_buffer_32_1 f2110(.wen(f2110_wen), .wdata(f2110_wdata), .clk(f2110_clk), .rst(f2110_rst), .rdata(f2110_rdata));
  assign f2110_clk = clk;
  assign f2110_rst = rst;
  // Bindings to f2110

  // f2112
  logic [0:0] f2112_wen;
  logic [31:0] f2112_wdata;
  logic [0:0] f2112_clk;
  logic [0:0] f2112_rst;
  logic [31:0] f2112_rdata;
  sr_buffer_32_1 f2112(.wen(f2112_wen), .wdata(f2112_wdata), .clk(f2112_clk), .rst(f2112_rst), .rdata(f2112_rdata));
  assign f2112_clk = clk;
  assign f2112_rst = rst;
  // Bindings to f2112

  // f2114
  logic [0:0] f2114_wen;
  logic [31:0] f2114_wdata;
  logic [0:0] f2114_clk;
  logic [0:0] f2114_rst;
  logic [31:0] f2114_rdata;
  sr_buffer_32_1 f2114(.wen(f2114_wen), .wdata(f2114_wdata), .clk(f2114_clk), .rst(f2114_rst), .rdata(f2114_rdata));
  assign f2114_clk = clk;
  assign f2114_rst = rst;
  // Bindings to f2114

  // f2116
  logic [0:0] f2116_wen;
  logic [31:0] f2116_wdata;
  logic [0:0] f2116_clk;
  logic [0:0] f2116_rst;
  logic [31:0] f2116_rdata;
  sr_buffer_32_1 f2116(.wen(f2116_wen), .wdata(f2116_wdata), .clk(f2116_clk), .rst(f2116_rst), .rdata(f2116_rdata));
  assign f2116_clk = clk;
  assign f2116_rst = rst;
  // Bindings to f2116

  // f2118
  logic [0:0] f2118_wen;
  logic [31:0] f2118_wdata;
  logic [0:0] f2118_clk;
  logic [0:0] f2118_rst;
  logic [31:0] f2118_rdata;
  sr_buffer_32_1 f2118(.wen(f2118_wen), .wdata(f2118_wdata), .clk(f2118_clk), .rst(f2118_rst), .rdata(f2118_rdata));
  assign f2118_clk = clk;
  assign f2118_rst = rst;
  // Bindings to f2118

  // f2120
  logic [0:0] f2120_wen;
  logic [31:0] f2120_wdata;
  logic [0:0] f2120_clk;
  logic [0:0] f2120_rst;
  logic [31:0] f2120_rdata;
  sr_buffer_32_1 f2120(.wen(f2120_wen), .wdata(f2120_wdata), .clk(f2120_clk), .rst(f2120_rst), .rdata(f2120_rdata));
  assign f2120_clk = clk;
  assign f2120_rst = rst;
  // Bindings to f2120

  // f2122
  logic [0:0] f2122_wen;
  logic [31:0] f2122_wdata;
  logic [0:0] f2122_clk;
  logic [0:0] f2122_rst;
  logic [31:0] f2122_rdata;
  sr_buffer_32_1 f2122(.wen(f2122_wen), .wdata(f2122_wdata), .clk(f2122_clk), .rst(f2122_rst), .rdata(f2122_rdata));
  assign f2122_clk = clk;
  assign f2122_rst = rst;
  // Bindings to f2122

  // f2124
  logic [0:0] f2124_wen;
  logic [31:0] f2124_wdata;
  logic [0:0] f2124_clk;
  logic [0:0] f2124_rst;
  logic [31:0] f2124_rdata;
  sr_buffer_32_1 f2124(.wen(f2124_wen), .wdata(f2124_wdata), .clk(f2124_clk), .rst(f2124_rst), .rdata(f2124_rdata));
  assign f2124_clk = clk;
  assign f2124_rst = rst;
  // Bindings to f2124

  // f2126
  logic [0:0] f2126_wen;
  logic [31:0] f2126_wdata;
  logic [0:0] f2126_clk;
  logic [0:0] f2126_rst;
  logic [31:0] f2126_rdata;
  sr_buffer_32_1 f2126(.wen(f2126_wen), .wdata(f2126_wdata), .clk(f2126_clk), .rst(f2126_rst), .rdata(f2126_rdata));
  assign f2126_clk = clk;
  assign f2126_rst = rst;
  // Bindings to f2126

  // f2128
  logic [0:0] f2128_wen;
  logic [31:0] f2128_wdata;
  logic [0:0] f2128_clk;
  logic [0:0] f2128_rst;
  logic [31:0] f2128_rdata;
  sr_buffer_32_1 f2128(.wen(f2128_wen), .wdata(f2128_wdata), .clk(f2128_clk), .rst(f2128_rst), .rdata(f2128_rdata));
  assign f2128_clk = clk;
  assign f2128_rst = rst;
  // Bindings to f2128

  // f2130
  logic [0:0] f2130_wen;
  logic [31:0] f2130_wdata;
  logic [0:0] f2130_clk;
  logic [0:0] f2130_rst;
  logic [31:0] f2130_rdata;
  sr_buffer_32_1 f2130(.wen(f2130_wen), .wdata(f2130_wdata), .clk(f2130_clk), .rst(f2130_rst), .rdata(f2130_rdata));
  assign f2130_clk = clk;
  assign f2130_rst = rst;
  // Bindings to f2130

  // f2132
  logic [0:0] f2132_wen;
  logic [31:0] f2132_wdata;
  logic [0:0] f2132_clk;
  logic [0:0] f2132_rst;
  logic [31:0] f2132_rdata;
  sr_buffer_32_1 f2132(.wen(f2132_wen), .wdata(f2132_wdata), .clk(f2132_clk), .rst(f2132_rst), .rdata(f2132_rdata));
  assign f2132_clk = clk;
  assign f2132_rst = rst;
  // Bindings to f2132

  // f2134
  logic [0:0] f2134_wen;
  logic [31:0] f2134_wdata;
  logic [0:0] f2134_clk;
  logic [0:0] f2134_rst;
  logic [31:0] f2134_rdata;
  sr_buffer_32_1 f2134(.wen(f2134_wen), .wdata(f2134_wdata), .clk(f2134_clk), .rst(f2134_rst), .rdata(f2134_rdata));
  assign f2134_clk = clk;
  assign f2134_rst = rst;
  // Bindings to f2134

  // f2136
  logic [0:0] f2136_wen;
  logic [31:0] f2136_wdata;
  logic [0:0] f2136_clk;
  logic [0:0] f2136_rst;
  logic [31:0] f2136_rdata;
  sr_buffer_32_1 f2136(.wen(f2136_wen), .wdata(f2136_wdata), .clk(f2136_clk), .rst(f2136_rst), .rdata(f2136_rdata));
  assign f2136_clk = clk;
  assign f2136_rst = rst;
  // Bindings to f2136

  // f2138
  logic [0:0] f2138_wen;
  logic [31:0] f2138_wdata;
  logic [0:0] f2138_clk;
  logic [0:0] f2138_rst;
  logic [31:0] f2138_rdata;
  sr_buffer_32_1 f2138(.wen(f2138_wen), .wdata(f2138_wdata), .clk(f2138_clk), .rst(f2138_rst), .rdata(f2138_rdata));
  assign f2138_clk = clk;
  assign f2138_rst = rst;
  // Bindings to f2138

  // f2140
  logic [0:0] f2140_wen;
  logic [31:0] f2140_wdata;
  logic [0:0] f2140_clk;
  logic [0:0] f2140_rst;
  logic [31:0] f2140_rdata;
  sr_buffer_32_1 f2140(.wen(f2140_wen), .wdata(f2140_wdata), .clk(f2140_clk), .rst(f2140_rst), .rdata(f2140_rdata));
  assign f2140_clk = clk;
  assign f2140_rst = rst;
  // Bindings to f2140

  // f2142
  logic [0:0] f2142_wen;
  logic [31:0] f2142_wdata;
  logic [0:0] f2142_clk;
  logic [0:0] f2142_rst;
  logic [31:0] f2142_rdata;
  sr_buffer_32_1 f2142(.wen(f2142_wen), .wdata(f2142_wdata), .clk(f2142_clk), .rst(f2142_rst), .rdata(f2142_rdata));
  assign f2142_clk = clk;
  assign f2142_rst = rst;
  // Bindings to f2142

  // f2144
  logic [0:0] f2144_wen;
  logic [31:0] f2144_wdata;
  logic [0:0] f2144_clk;
  logic [0:0] f2144_rst;
  logic [31:0] f2144_rdata;
  sr_buffer_32_1 f2144(.wen(f2144_wen), .wdata(f2144_wdata), .clk(f2144_clk), .rst(f2144_rst), .rdata(f2144_rdata));
  assign f2144_clk = clk;
  assign f2144_rst = rst;
  // Bindings to f2144

  // f2146
  logic [0:0] f2146_wen;
  logic [31:0] f2146_wdata;
  logic [0:0] f2146_clk;
  logic [0:0] f2146_rst;
  logic [31:0] f2146_rdata;
  sr_buffer_32_1 f2146(.wen(f2146_wen), .wdata(f2146_wdata), .clk(f2146_clk), .rst(f2146_rst), .rdata(f2146_rdata));
  assign f2146_clk = clk;
  assign f2146_rst = rst;
  // Bindings to f2146

  // f2148
  logic [0:0] f2148_wen;
  logic [31:0] f2148_wdata;
  logic [0:0] f2148_clk;
  logic [0:0] f2148_rst;
  logic [31:0] f2148_rdata;
  sr_buffer_32_1 f2148(.wen(f2148_wen), .wdata(f2148_wdata), .clk(f2148_clk), .rst(f2148_rst), .rdata(f2148_rdata));
  assign f2148_clk = clk;
  assign f2148_rst = rst;
  // Bindings to f2148

  // f2150
  logic [0:0] f2150_wen;
  logic [31:0] f2150_wdata;
  logic [0:0] f2150_clk;
  logic [0:0] f2150_rst;
  logic [31:0] f2150_rdata;
  sr_buffer_32_1 f2150(.wen(f2150_wen), .wdata(f2150_wdata), .clk(f2150_clk), .rst(f2150_rst), .rdata(f2150_rdata));
  assign f2150_clk = clk;
  assign f2150_rst = rst;
  // Bindings to f2150

  // f2152
  logic [0:0] f2152_wen;
  logic [31:0] f2152_wdata;
  logic [0:0] f2152_clk;
  logic [0:0] f2152_rst;
  logic [31:0] f2152_rdata;
  sr_buffer_32_1 f2152(.wen(f2152_wen), .wdata(f2152_wdata), .clk(f2152_clk), .rst(f2152_rst), .rdata(f2152_rdata));
  assign f2152_clk = clk;
  assign f2152_rst = rst;
  // Bindings to f2152

  // f2154
  logic [0:0] f2154_wen;
  logic [31:0] f2154_wdata;
  logic [0:0] f2154_clk;
  logic [0:0] f2154_rst;
  logic [31:0] f2154_rdata;
  sr_buffer_32_1 f2154(.wen(f2154_wen), .wdata(f2154_wdata), .clk(f2154_clk), .rst(f2154_rst), .rdata(f2154_rdata));
  assign f2154_clk = clk;
  assign f2154_rst = rst;
  // Bindings to f2154

  // f2156
  logic [0:0] f2156_wen;
  logic [31:0] f2156_wdata;
  logic [0:0] f2156_clk;
  logic [0:0] f2156_rst;
  logic [31:0] f2156_rdata;
  sr_buffer_32_1 f2156(.wen(f2156_wen), .wdata(f2156_wdata), .clk(f2156_clk), .rst(f2156_rst), .rdata(f2156_rdata));
  assign f2156_clk = clk;
  assign f2156_rst = rst;
  // Bindings to f2156

  // f2158
  logic [0:0] f2158_wen;
  logic [31:0] f2158_wdata;
  logic [0:0] f2158_clk;
  logic [0:0] f2158_rst;
  logic [31:0] f2158_rdata;
  sr_buffer_32_1 f2158(.wen(f2158_wen), .wdata(f2158_wdata), .clk(f2158_clk), .rst(f2158_rst), .rdata(f2158_rdata));
  assign f2158_clk = clk;
  assign f2158_rst = rst;
  // Bindings to f2158

  // f2160
  logic [0:0] f2160_wen;
  logic [31:0] f2160_wdata;
  logic [0:0] f2160_clk;
  logic [0:0] f2160_rst;
  logic [31:0] f2160_rdata;
  sr_buffer_32_1 f2160(.wen(f2160_wen), .wdata(f2160_wdata), .clk(f2160_clk), .rst(f2160_rst), .rdata(f2160_rdata));
  assign f2160_clk = clk;
  assign f2160_rst = rst;
  // Bindings to f2160

  // f2162
  logic [0:0] f2162_wen;
  logic [31:0] f2162_wdata;
  logic [0:0] f2162_clk;
  logic [0:0] f2162_rst;
  logic [31:0] f2162_rdata;
  sr_buffer_32_1 f2162(.wen(f2162_wen), .wdata(f2162_wdata), .clk(f2162_clk), .rst(f2162_rst), .rdata(f2162_rdata));
  assign f2162_clk = clk;
  assign f2162_rst = rst;
  // Bindings to f2162

  // f2164
  logic [0:0] f2164_wen;
  logic [31:0] f2164_wdata;
  logic [0:0] f2164_clk;
  logic [0:0] f2164_rst;
  logic [31:0] f2164_rdata;
  sr_buffer_32_1 f2164(.wen(f2164_wen), .wdata(f2164_wdata), .clk(f2164_clk), .rst(f2164_rst), .rdata(f2164_rdata));
  assign f2164_clk = clk;
  assign f2164_rst = rst;
  // Bindings to f2164

  // f2166
  logic [0:0] f2166_wen;
  logic [31:0] f2166_wdata;
  logic [0:0] f2166_clk;
  logic [0:0] f2166_rst;
  logic [31:0] f2166_rdata;
  sr_buffer_32_1 f2166(.wen(f2166_wen), .wdata(f2166_wdata), .clk(f2166_clk), .rst(f2166_rst), .rdata(f2166_rdata));
  assign f2166_clk = clk;
  assign f2166_rst = rst;
  // Bindings to f2166

  // f2168
  logic [0:0] f2168_wen;
  logic [31:0] f2168_wdata;
  logic [0:0] f2168_clk;
  logic [0:0] f2168_rst;
  logic [31:0] f2168_rdata;
  sr_buffer_32_1 f2168(.wen(f2168_wen), .wdata(f2168_wdata), .clk(f2168_clk), .rst(f2168_rst), .rdata(f2168_rdata));
  assign f2168_clk = clk;
  assign f2168_rst = rst;
  // Bindings to f2168

  // f2170
  logic [0:0] f2170_wen;
  logic [31:0] f2170_wdata;
  logic [0:0] f2170_clk;
  logic [0:0] f2170_rst;
  logic [31:0] f2170_rdata;
  sr_buffer_32_1 f2170(.wen(f2170_wen), .wdata(f2170_wdata), .clk(f2170_clk), .rst(f2170_rst), .rdata(f2170_rdata));
  assign f2170_clk = clk;
  assign f2170_rst = rst;
  // Bindings to f2170

  // f2172
  logic [0:0] f2172_wen;
  logic [31:0] f2172_wdata;
  logic [0:0] f2172_clk;
  logic [0:0] f2172_rst;
  logic [31:0] f2172_rdata;
  sr_buffer_32_1 f2172(.wen(f2172_wen), .wdata(f2172_wdata), .clk(f2172_clk), .rst(f2172_rst), .rdata(f2172_rdata));
  assign f2172_clk = clk;
  assign f2172_rst = rst;
  // Bindings to f2172

  // f2174
  logic [0:0] f2174_wen;
  logic [31:0] f2174_wdata;
  logic [0:0] f2174_clk;
  logic [0:0] f2174_rst;
  logic [31:0] f2174_rdata;
  sr_buffer_32_1 f2174(.wen(f2174_wen), .wdata(f2174_wdata), .clk(f2174_clk), .rst(f2174_rst), .rdata(f2174_rdata));
  assign f2174_clk = clk;
  assign f2174_rst = rst;
  // Bindings to f2174

  // f2176
  logic [0:0] f2176_wen;
  logic [31:0] f2176_wdata;
  logic [0:0] f2176_clk;
  logic [0:0] f2176_rst;
  logic [31:0] f2176_rdata;
  sr_buffer_32_1 f2176(.wen(f2176_wen), .wdata(f2176_wdata), .clk(f2176_clk), .rst(f2176_rst), .rdata(f2176_rdata));
  assign f2176_clk = clk;
  assign f2176_rst = rst;
  // Bindings to f2176

  // f2178
  logic [0:0] f2178_wen;
  logic [31:0] f2178_wdata;
  logic [0:0] f2178_clk;
  logic [0:0] f2178_rst;
  logic [31:0] f2178_rdata;
  sr_buffer_32_1 f2178(.wen(f2178_wen), .wdata(f2178_wdata), .clk(f2178_clk), .rst(f2178_rst), .rdata(f2178_rdata));
  assign f2178_clk = clk;
  assign f2178_rst = rst;
  // Bindings to f2178

  // f2180
  logic [0:0] f2180_wen;
  logic [31:0] f2180_wdata;
  logic [0:0] f2180_clk;
  logic [0:0] f2180_rst;
  logic [31:0] f2180_rdata;
  sr_buffer_32_1 f2180(.wen(f2180_wen), .wdata(f2180_wdata), .clk(f2180_clk), .rst(f2180_rst), .rdata(f2180_rdata));
  assign f2180_clk = clk;
  assign f2180_rst = rst;
  // Bindings to f2180

  // f2182
  logic [0:0] f2182_wen;
  logic [31:0] f2182_wdata;
  logic [0:0] f2182_clk;
  logic [0:0] f2182_rst;
  logic [31:0] f2182_rdata;
  sr_buffer_32_1 f2182(.wen(f2182_wen), .wdata(f2182_wdata), .clk(f2182_clk), .rst(f2182_rst), .rdata(f2182_rdata));
  assign f2182_clk = clk;
  assign f2182_rst = rst;
  // Bindings to f2182

  // f2184
  logic [0:0] f2184_wen;
  logic [31:0] f2184_wdata;
  logic [0:0] f2184_clk;
  logic [0:0] f2184_rst;
  logic [31:0] f2184_rdata;
  sr_buffer_32_1 f2184(.wen(f2184_wen), .wdata(f2184_wdata), .clk(f2184_clk), .rst(f2184_rst), .rdata(f2184_rdata));
  assign f2184_clk = clk;
  assign f2184_rst = rst;
  // Bindings to f2184

  // f2186
  logic [0:0] f2186_wen;
  logic [31:0] f2186_wdata;
  logic [0:0] f2186_clk;
  logic [0:0] f2186_rst;
  logic [31:0] f2186_rdata;
  sr_buffer_32_1 f2186(.wen(f2186_wen), .wdata(f2186_wdata), .clk(f2186_clk), .rst(f2186_rst), .rdata(f2186_rdata));
  assign f2186_clk = clk;
  assign f2186_rst = rst;
  // Bindings to f2186

  // f2188
  logic [0:0] f2188_wen;
  logic [31:0] f2188_wdata;
  logic [0:0] f2188_clk;
  logic [0:0] f2188_rst;
  logic [31:0] f2188_rdata;
  sr_buffer_32_1 f2188(.wen(f2188_wen), .wdata(f2188_wdata), .clk(f2188_clk), .rst(f2188_rst), .rdata(f2188_rdata));
  assign f2188_clk = clk;
  assign f2188_rst = rst;
  // Bindings to f2188

  // f2190
  logic [0:0] f2190_wen;
  logic [31:0] f2190_wdata;
  logic [0:0] f2190_clk;
  logic [0:0] f2190_rst;
  logic [31:0] f2190_rdata;
  sr_buffer_32_1 f2190(.wen(f2190_wen), .wdata(f2190_wdata), .clk(f2190_clk), .rst(f2190_rst), .rdata(f2190_rdata));
  assign f2190_clk = clk;
  assign f2190_rst = rst;
  // Bindings to f2190

  // f2192
  logic [0:0] f2192_wen;
  logic [31:0] f2192_wdata;
  logic [0:0] f2192_clk;
  logic [0:0] f2192_rst;
  logic [31:0] f2192_rdata;
  sr_buffer_32_1 f2192(.wen(f2192_wen), .wdata(f2192_wdata), .clk(f2192_clk), .rst(f2192_rst), .rdata(f2192_rdata));
  assign f2192_clk = clk;
  assign f2192_rst = rst;
  // Bindings to f2192

  // f2194
  logic [0:0] f2194_wen;
  logic [31:0] f2194_wdata;
  logic [0:0] f2194_clk;
  logic [0:0] f2194_rst;
  logic [31:0] f2194_rdata;
  sr_buffer_32_1 f2194(.wen(f2194_wen), .wdata(f2194_wdata), .clk(f2194_clk), .rst(f2194_rst), .rdata(f2194_rdata));
  assign f2194_clk = clk;
  assign f2194_rst = rst;
  // Bindings to f2194

  // f2196
  logic [0:0] f2196_wen;
  logic [31:0] f2196_wdata;
  logic [0:0] f2196_clk;
  logic [0:0] f2196_rst;
  logic [31:0] f2196_rdata;
  sr_buffer_32_1 f2196(.wen(f2196_wen), .wdata(f2196_wdata), .clk(f2196_clk), .rst(f2196_rst), .rdata(f2196_rdata));
  assign f2196_clk = clk;
  assign f2196_rst = rst;
  // Bindings to f2196

  // f2198
  logic [0:0] f2198_wen;
  logic [31:0] f2198_wdata;
  logic [0:0] f2198_clk;
  logic [0:0] f2198_rst;
  logic [31:0] f2198_rdata;
  sr_buffer_32_1 f2198(.wen(f2198_wen), .wdata(f2198_wdata), .clk(f2198_clk), .rst(f2198_rst), .rdata(f2198_rdata));
  assign f2198_clk = clk;
  assign f2198_rst = rst;
  // Bindings to f2198

  // f2200
  logic [0:0] f2200_wen;
  logic [31:0] f2200_wdata;
  logic [0:0] f2200_clk;
  logic [0:0] f2200_rst;
  logic [31:0] f2200_rdata;
  sr_buffer_32_1 f2200(.wen(f2200_wen), .wdata(f2200_wdata), .clk(f2200_clk), .rst(f2200_rst), .rdata(f2200_rdata));
  assign f2200_clk = clk;
  assign f2200_rst = rst;
  // Bindings to f2200

  // f2202
  logic [0:0] f2202_wen;
  logic [31:0] f2202_wdata;
  logic [0:0] f2202_clk;
  logic [0:0] f2202_rst;
  logic [31:0] f2202_rdata;
  sr_buffer_32_1 f2202(.wen(f2202_wen), .wdata(f2202_wdata), .clk(f2202_clk), .rst(f2202_rst), .rdata(f2202_rdata));
  assign f2202_clk = clk;
  assign f2202_rst = rst;
  // Bindings to f2202

  // f2204
  logic [0:0] f2204_wen;
  logic [31:0] f2204_wdata;
  logic [0:0] f2204_clk;
  logic [0:0] f2204_rst;
  logic [31:0] f2204_rdata;
  sr_buffer_32_1 f2204(.wen(f2204_wen), .wdata(f2204_wdata), .clk(f2204_clk), .rst(f2204_rst), .rdata(f2204_rdata));
  assign f2204_clk = clk;
  assign f2204_rst = rst;
  // Bindings to f2204

  // f2206
  logic [0:0] f2206_wen;
  logic [31:0] f2206_wdata;
  logic [0:0] f2206_clk;
  logic [0:0] f2206_rst;
  logic [31:0] f2206_rdata;
  sr_buffer_32_1 f2206(.wen(f2206_wen), .wdata(f2206_wdata), .clk(f2206_clk), .rst(f2206_rst), .rdata(f2206_rdata));
  assign f2206_clk = clk;
  assign f2206_rst = rst;
  // Bindings to f2206

  // f2208
  logic [0:0] f2208_wen;
  logic [31:0] f2208_wdata;
  logic [0:0] f2208_clk;
  logic [0:0] f2208_rst;
  logic [31:0] f2208_rdata;
  sr_buffer_32_1 f2208(.wen(f2208_wen), .wdata(f2208_wdata), .clk(f2208_clk), .rst(f2208_rst), .rdata(f2208_rdata));
  assign f2208_clk = clk;
  assign f2208_rst = rst;
  // Bindings to f2208

  // f2210
  logic [0:0] f2210_wen;
  logic [31:0] f2210_wdata;
  logic [0:0] f2210_clk;
  logic [0:0] f2210_rst;
  logic [31:0] f2210_rdata;
  sr_buffer_32_1 f2210(.wen(f2210_wen), .wdata(f2210_wdata), .clk(f2210_clk), .rst(f2210_rst), .rdata(f2210_rdata));
  assign f2210_clk = clk;
  assign f2210_rst = rst;
  // Bindings to f2210

  // f2212
  logic [0:0] f2212_wen;
  logic [31:0] f2212_wdata;
  logic [0:0] f2212_clk;
  logic [0:0] f2212_rst;
  logic [31:0] f2212_rdata;
  sr_buffer_32_1 f2212(.wen(f2212_wen), .wdata(f2212_wdata), .clk(f2212_clk), .rst(f2212_rst), .rdata(f2212_rdata));
  assign f2212_clk = clk;
  assign f2212_rst = rst;
  // Bindings to f2212

  // f2214
  logic [0:0] f2214_wen;
  logic [31:0] f2214_wdata;
  logic [0:0] f2214_clk;
  logic [0:0] f2214_rst;
  logic [31:0] f2214_rdata;
  sr_buffer_32_1 f2214(.wen(f2214_wen), .wdata(f2214_wdata), .clk(f2214_clk), .rst(f2214_rst), .rdata(f2214_rdata));
  assign f2214_clk = clk;
  assign f2214_rst = rst;
  // Bindings to f2214

  // f2216
  logic [0:0] f2216_wen;
  logic [31:0] f2216_wdata;
  logic [0:0] f2216_clk;
  logic [0:0] f2216_rst;
  logic [31:0] f2216_rdata;
  sr_buffer_32_1 f2216(.wen(f2216_wen), .wdata(f2216_wdata), .clk(f2216_clk), .rst(f2216_rst), .rdata(f2216_rdata));
  assign f2216_clk = clk;
  assign f2216_rst = rst;
  // Bindings to f2216

  // f2218
  logic [0:0] f2218_wen;
  logic [31:0] f2218_wdata;
  logic [0:0] f2218_clk;
  logic [0:0] f2218_rst;
  logic [31:0] f2218_rdata;
  sr_buffer_32_1 f2218(.wen(f2218_wen), .wdata(f2218_wdata), .clk(f2218_clk), .rst(f2218_rst), .rdata(f2218_rdata));
  assign f2218_clk = clk;
  assign f2218_rst = rst;
  // Bindings to f2218

  // f2220
  logic [0:0] f2220_wen;
  logic [31:0] f2220_wdata;
  logic [0:0] f2220_clk;
  logic [0:0] f2220_rst;
  logic [31:0] f2220_rdata;
  sr_buffer_32_1 f2220(.wen(f2220_wen), .wdata(f2220_wdata), .clk(f2220_clk), .rst(f2220_rst), .rdata(f2220_rdata));
  assign f2220_clk = clk;
  assign f2220_rst = rst;
  // Bindings to f2220

  // f2222
  logic [0:0] f2222_wen;
  logic [31:0] f2222_wdata;
  logic [0:0] f2222_clk;
  logic [0:0] f2222_rst;
  logic [31:0] f2222_rdata;
  sr_buffer_32_1 f2222(.wen(f2222_wen), .wdata(f2222_wdata), .clk(f2222_clk), .rst(f2222_rst), .rdata(f2222_rdata));
  assign f2222_clk = clk;
  assign f2222_rst = rst;
  // Bindings to f2222

  // f2224
  logic [0:0] f2224_wen;
  logic [31:0] f2224_wdata;
  logic [0:0] f2224_clk;
  logic [0:0] f2224_rst;
  logic [31:0] f2224_rdata;
  sr_buffer_32_1 f2224(.wen(f2224_wen), .wdata(f2224_wdata), .clk(f2224_clk), .rst(f2224_rst), .rdata(f2224_rdata));
  assign f2224_clk = clk;
  assign f2224_rst = rst;
  // Bindings to f2224

  // f2226
  logic [0:0] f2226_wen;
  logic [31:0] f2226_wdata;
  logic [0:0] f2226_clk;
  logic [0:0] f2226_rst;
  logic [31:0] f2226_rdata;
  sr_buffer_32_1 f2226(.wen(f2226_wen), .wdata(f2226_wdata), .clk(f2226_clk), .rst(f2226_rst), .rdata(f2226_rdata));
  assign f2226_clk = clk;
  assign f2226_rst = rst;
  // Bindings to f2226

  // f2228
  logic [0:0] f2228_wen;
  logic [31:0] f2228_wdata;
  logic [0:0] f2228_clk;
  logic [0:0] f2228_rst;
  logic [31:0] f2228_rdata;
  sr_buffer_32_1 f2228(.wen(f2228_wen), .wdata(f2228_wdata), .clk(f2228_clk), .rst(f2228_rst), .rdata(f2228_rdata));
  assign f2228_clk = clk;
  assign f2228_rst = rst;
  // Bindings to f2228

  // f2230
  logic [0:0] f2230_wen;
  logic [31:0] f2230_wdata;
  logic [0:0] f2230_clk;
  logic [0:0] f2230_rst;
  logic [31:0] f2230_rdata;
  sr_buffer_32_1 f2230(.wen(f2230_wen), .wdata(f2230_wdata), .clk(f2230_clk), .rst(f2230_rst), .rdata(f2230_rdata));
  assign f2230_clk = clk;
  assign f2230_rst = rst;
  // Bindings to f2230

  // f2232
  logic [0:0] f2232_wen;
  logic [31:0] f2232_wdata;
  logic [0:0] f2232_clk;
  logic [0:0] f2232_rst;
  logic [31:0] f2232_rdata;
  sr_buffer_32_1 f2232(.wen(f2232_wen), .wdata(f2232_wdata), .clk(f2232_clk), .rst(f2232_rst), .rdata(f2232_rdata));
  assign f2232_clk = clk;
  assign f2232_rst = rst;
  // Bindings to f2232

  // f2234
  logic [0:0] f2234_wen;
  logic [31:0] f2234_wdata;
  logic [0:0] f2234_clk;
  logic [0:0] f2234_rst;
  logic [31:0] f2234_rdata;
  sr_buffer_32_1 f2234(.wen(f2234_wen), .wdata(f2234_wdata), .clk(f2234_clk), .rst(f2234_rst), .rdata(f2234_rdata));
  assign f2234_clk = clk;
  assign f2234_rst = rst;
  // Bindings to f2234

  // f2236
  logic [0:0] f2236_wen;
  logic [31:0] f2236_wdata;
  logic [0:0] f2236_clk;
  logic [0:0] f2236_rst;
  logic [31:0] f2236_rdata;
  sr_buffer_32_1 f2236(.wen(f2236_wen), .wdata(f2236_wdata), .clk(f2236_clk), .rst(f2236_rst), .rdata(f2236_rdata));
  assign f2236_clk = clk;
  assign f2236_rst = rst;
  // Bindings to f2236

  // f2238
  logic [0:0] f2238_wen;
  logic [31:0] f2238_wdata;
  logic [0:0] f2238_clk;
  logic [0:0] f2238_rst;
  logic [31:0] f2238_rdata;
  sr_buffer_32_1 f2238(.wen(f2238_wen), .wdata(f2238_wdata), .clk(f2238_clk), .rst(f2238_rst), .rdata(f2238_rdata));
  assign f2238_clk = clk;
  assign f2238_rst = rst;
  // Bindings to f2238

  // f2240
  logic [0:0] f2240_wen;
  logic [31:0] f2240_wdata;
  logic [0:0] f2240_clk;
  logic [0:0] f2240_rst;
  logic [31:0] f2240_rdata;
  sr_buffer_32_1 f2240(.wen(f2240_wen), .wdata(f2240_wdata), .clk(f2240_clk), .rst(f2240_rst), .rdata(f2240_rdata));
  assign f2240_clk = clk;
  assign f2240_rst = rst;
  // Bindings to f2240

  // f2242
  logic [0:0] f2242_wen;
  logic [31:0] f2242_wdata;
  logic [0:0] f2242_clk;
  logic [0:0] f2242_rst;
  logic [31:0] f2242_rdata;
  sr_buffer_32_1 f2242(.wen(f2242_wen), .wdata(f2242_wdata), .clk(f2242_clk), .rst(f2242_rst), .rdata(f2242_rdata));
  assign f2242_clk = clk;
  assign f2242_rst = rst;
  // Bindings to f2242

  // f2244
  logic [0:0] f2244_wen;
  logic [31:0] f2244_wdata;
  logic [0:0] f2244_clk;
  logic [0:0] f2244_rst;
  logic [31:0] f2244_rdata;
  sr_buffer_32_1 f2244(.wen(f2244_wen), .wdata(f2244_wdata), .clk(f2244_clk), .rst(f2244_rst), .rdata(f2244_rdata));
  assign f2244_clk = clk;
  assign f2244_rst = rst;
  // Bindings to f2244

  // f2246
  logic [0:0] f2246_wen;
  logic [31:0] f2246_wdata;
  logic [0:0] f2246_clk;
  logic [0:0] f2246_rst;
  logic [31:0] f2246_rdata;
  sr_buffer_32_1 f2246(.wen(f2246_wen), .wdata(f2246_wdata), .clk(f2246_clk), .rst(f2246_rst), .rdata(f2246_rdata));
  assign f2246_clk = clk;
  assign f2246_rst = rst;
  // Bindings to f2246

  // f2248
  logic [0:0] f2248_wen;
  logic [31:0] f2248_wdata;
  logic [0:0] f2248_clk;
  logic [0:0] f2248_rst;
  logic [31:0] f2248_rdata;
  sr_buffer_32_1 f2248(.wen(f2248_wen), .wdata(f2248_wdata), .clk(f2248_clk), .rst(f2248_rst), .rdata(f2248_rdata));
  assign f2248_clk = clk;
  assign f2248_rst = rst;
  // Bindings to f2248

  // f2250
  logic [0:0] f2250_wen;
  logic [31:0] f2250_wdata;
  logic [0:0] f2250_clk;
  logic [0:0] f2250_rst;
  logic [31:0] f2250_rdata;
  sr_buffer_32_1 f2250(.wen(f2250_wen), .wdata(f2250_wdata), .clk(f2250_clk), .rst(f2250_rst), .rdata(f2250_rdata));
  assign f2250_clk = clk;
  assign f2250_rst = rst;
  // Bindings to f2250

  // f2252
  logic [0:0] f2252_wen;
  logic [31:0] f2252_wdata;
  logic [0:0] f2252_clk;
  logic [0:0] f2252_rst;
  logic [31:0] f2252_rdata;
  sr_buffer_32_1 f2252(.wen(f2252_wen), .wdata(f2252_wdata), .clk(f2252_clk), .rst(f2252_rst), .rdata(f2252_rdata));
  assign f2252_clk = clk;
  assign f2252_rst = rst;
  // Bindings to f2252

  // f2254
  logic [0:0] f2254_wen;
  logic [31:0] f2254_wdata;
  logic [0:0] f2254_clk;
  logic [0:0] f2254_rst;
  logic [31:0] f2254_rdata;
  sr_buffer_32_1 f2254(.wen(f2254_wen), .wdata(f2254_wdata), .clk(f2254_clk), .rst(f2254_rst), .rdata(f2254_rdata));
  assign f2254_clk = clk;
  assign f2254_rst = rst;
  // Bindings to f2254

  // f2256
  logic [0:0] f2256_wen;
  logic [31:0] f2256_wdata;
  logic [0:0] f2256_clk;
  logic [0:0] f2256_rst;
  logic [31:0] f2256_rdata;
  sr_buffer_32_1 f2256(.wen(f2256_wen), .wdata(f2256_wdata), .clk(f2256_clk), .rst(f2256_rst), .rdata(f2256_rdata));
  assign f2256_clk = clk;
  assign f2256_rst = rst;
  // Bindings to f2256

  // f2258
  logic [0:0] f2258_wen;
  logic [31:0] f2258_wdata;
  logic [0:0] f2258_clk;
  logic [0:0] f2258_rst;
  logic [31:0] f2258_rdata;
  sr_buffer_32_1 f2258(.wen(f2258_wen), .wdata(f2258_wdata), .clk(f2258_clk), .rst(f2258_rst), .rdata(f2258_rdata));
  assign f2258_clk = clk;
  assign f2258_rst = rst;
  // Bindings to f2258

  // f2260
  logic [0:0] f2260_wen;
  logic [31:0] f2260_wdata;
  logic [0:0] f2260_clk;
  logic [0:0] f2260_rst;
  logic [31:0] f2260_rdata;
  sr_buffer_32_1 f2260(.wen(f2260_wen), .wdata(f2260_wdata), .clk(f2260_clk), .rst(f2260_rst), .rdata(f2260_rdata));
  assign f2260_clk = clk;
  assign f2260_rst = rst;
  // Bindings to f2260

  // f2262
  logic [0:0] f2262_wen;
  logic [31:0] f2262_wdata;
  logic [0:0] f2262_clk;
  logic [0:0] f2262_rst;
  logic [31:0] f2262_rdata;
  sr_buffer_32_1 f2262(.wen(f2262_wen), .wdata(f2262_wdata), .clk(f2262_clk), .rst(f2262_rst), .rdata(f2262_rdata));
  assign f2262_clk = clk;
  assign f2262_rst = rst;
  // Bindings to f2262

  // f2264
  logic [0:0] f2264_wen;
  logic [31:0] f2264_wdata;
  logic [0:0] f2264_clk;
  logic [0:0] f2264_rst;
  logic [31:0] f2264_rdata;
  sr_buffer_32_1 f2264(.wen(f2264_wen), .wdata(f2264_wdata), .clk(f2264_clk), .rst(f2264_rst), .rdata(f2264_rdata));
  assign f2264_clk = clk;
  assign f2264_rst = rst;
  // Bindings to f2264

  // f2266
  logic [0:0] f2266_wen;
  logic [31:0] f2266_wdata;
  logic [0:0] f2266_clk;
  logic [0:0] f2266_rst;
  logic [31:0] f2266_rdata;
  sr_buffer_32_1 f2266(.wen(f2266_wen), .wdata(f2266_wdata), .clk(f2266_clk), .rst(f2266_rst), .rdata(f2266_rdata));
  assign f2266_clk = clk;
  assign f2266_rst = rst;
  // Bindings to f2266

  // f2268
  logic [0:0] f2268_wen;
  logic [31:0] f2268_wdata;
  logic [0:0] f2268_clk;
  logic [0:0] f2268_rst;
  logic [31:0] f2268_rdata;
  sr_buffer_32_1 f2268(.wen(f2268_wen), .wdata(f2268_wdata), .clk(f2268_clk), .rst(f2268_rst), .rdata(f2268_rdata));
  assign f2268_clk = clk;
  assign f2268_rst = rst;
  // Bindings to f2268

  // f2270
  logic [0:0] f2270_wen;
  logic [31:0] f2270_wdata;
  logic [0:0] f2270_clk;
  logic [0:0] f2270_rst;
  logic [31:0] f2270_rdata;
  sr_buffer_32_1 f2270(.wen(f2270_wen), .wdata(f2270_wdata), .clk(f2270_clk), .rst(f2270_rst), .rdata(f2270_rdata));
  assign f2270_clk = clk;
  assign f2270_rst = rst;
  // Bindings to f2270

  // f2272
  logic [0:0] f2272_wen;
  logic [31:0] f2272_wdata;
  logic [0:0] f2272_clk;
  logic [0:0] f2272_rst;
  logic [31:0] f2272_rdata;
  sr_buffer_32_1 f2272(.wen(f2272_wen), .wdata(f2272_wdata), .clk(f2272_clk), .rst(f2272_rst), .rdata(f2272_rdata));
  assign f2272_clk = clk;
  assign f2272_rst = rst;
  // Bindings to f2272

  // f2274
  logic [0:0] f2274_wen;
  logic [31:0] f2274_wdata;
  logic [0:0] f2274_clk;
  logic [0:0] f2274_rst;
  logic [31:0] f2274_rdata;
  sr_buffer_32_1 f2274(.wen(f2274_wen), .wdata(f2274_wdata), .clk(f2274_clk), .rst(f2274_rst), .rdata(f2274_rdata));
  assign f2274_clk = clk;
  assign f2274_rst = rst;
  // Bindings to f2274

  // f2276
  logic [0:0] f2276_wen;
  logic [31:0] f2276_wdata;
  logic [0:0] f2276_clk;
  logic [0:0] f2276_rst;
  logic [31:0] f2276_rdata;
  sr_buffer_32_1 f2276(.wen(f2276_wen), .wdata(f2276_wdata), .clk(f2276_clk), .rst(f2276_rst), .rdata(f2276_rdata));
  assign f2276_clk = clk;
  assign f2276_rst = rst;
  // Bindings to f2276

  // f2278
  logic [0:0] f2278_wen;
  logic [31:0] f2278_wdata;
  logic [0:0] f2278_clk;
  logic [0:0] f2278_rst;
  logic [31:0] f2278_rdata;
  sr_buffer_32_1 f2278(.wen(f2278_wen), .wdata(f2278_wdata), .clk(f2278_clk), .rst(f2278_rst), .rdata(f2278_rdata));
  assign f2278_clk = clk;
  assign f2278_rst = rst;
  // Bindings to f2278

  // f2280
  logic [0:0] f2280_wen;
  logic [31:0] f2280_wdata;
  logic [0:0] f2280_clk;
  logic [0:0] f2280_rst;
  logic [31:0] f2280_rdata;
  sr_buffer_32_1 f2280(.wen(f2280_wen), .wdata(f2280_wdata), .clk(f2280_clk), .rst(f2280_rst), .rdata(f2280_rdata));
  assign f2280_clk = clk;
  assign f2280_rst = rst;
  // Bindings to f2280

  // f2282
  logic [0:0] f2282_wen;
  logic [31:0] f2282_wdata;
  logic [0:0] f2282_clk;
  logic [0:0] f2282_rst;
  logic [31:0] f2282_rdata;
  sr_buffer_32_1 f2282(.wen(f2282_wen), .wdata(f2282_wdata), .clk(f2282_clk), .rst(f2282_rst), .rdata(f2282_rdata));
  assign f2282_clk = clk;
  assign f2282_rst = rst;
  // Bindings to f2282

  // f2284
  logic [0:0] f2284_wen;
  logic [31:0] f2284_wdata;
  logic [0:0] f2284_clk;
  logic [0:0] f2284_rst;
  logic [31:0] f2284_rdata;
  sr_buffer_32_1 f2284(.wen(f2284_wen), .wdata(f2284_wdata), .clk(f2284_clk), .rst(f2284_rst), .rdata(f2284_rdata));
  assign f2284_clk = clk;
  assign f2284_rst = rst;
  // Bindings to f2284

  // f2286
  logic [0:0] f2286_wen;
  logic [31:0] f2286_wdata;
  logic [0:0] f2286_clk;
  logic [0:0] f2286_rst;
  logic [31:0] f2286_rdata;
  sr_buffer_32_1 f2286(.wen(f2286_wen), .wdata(f2286_wdata), .clk(f2286_clk), .rst(f2286_rst), .rdata(f2286_rdata));
  assign f2286_clk = clk;
  assign f2286_rst = rst;
  // Bindings to f2286

  // f2288
  logic [0:0] f2288_wen;
  logic [31:0] f2288_wdata;
  logic [0:0] f2288_clk;
  logic [0:0] f2288_rst;
  logic [31:0] f2288_rdata;
  sr_buffer_32_1 f2288(.wen(f2288_wen), .wdata(f2288_wdata), .clk(f2288_clk), .rst(f2288_rst), .rdata(f2288_rdata));
  assign f2288_clk = clk;
  assign f2288_rst = rst;
  // Bindings to f2288

  // f2290
  logic [0:0] f2290_wen;
  logic [31:0] f2290_wdata;
  logic [0:0] f2290_clk;
  logic [0:0] f2290_rst;
  logic [31:0] f2290_rdata;
  sr_buffer_32_1 f2290(.wen(f2290_wen), .wdata(f2290_wdata), .clk(f2290_clk), .rst(f2290_rst), .rdata(f2290_rdata));
  assign f2290_clk = clk;
  assign f2290_rst = rst;
  // Bindings to f2290

  // f2292
  logic [0:0] f2292_wen;
  logic [31:0] f2292_wdata;
  logic [0:0] f2292_clk;
  logic [0:0] f2292_rst;
  logic [31:0] f2292_rdata;
  sr_buffer_32_1 f2292(.wen(f2292_wen), .wdata(f2292_wdata), .clk(f2292_clk), .rst(f2292_rst), .rdata(f2292_rdata));
  assign f2292_clk = clk;
  assign f2292_rst = rst;
  // Bindings to f2292

  // f2294
  logic [0:0] f2294_wen;
  logic [31:0] f2294_wdata;
  logic [0:0] f2294_clk;
  logic [0:0] f2294_rst;
  logic [31:0] f2294_rdata;
  sr_buffer_32_1 f2294(.wen(f2294_wen), .wdata(f2294_wdata), .clk(f2294_clk), .rst(f2294_rst), .rdata(f2294_rdata));
  assign f2294_clk = clk;
  assign f2294_rst = rst;
  // Bindings to f2294

  // f2296
  logic [0:0] f2296_wen;
  logic [31:0] f2296_wdata;
  logic [0:0] f2296_clk;
  logic [0:0] f2296_rst;
  logic [31:0] f2296_rdata;
  sr_buffer_32_1 f2296(.wen(f2296_wen), .wdata(f2296_wdata), .clk(f2296_clk), .rst(f2296_rst), .rdata(f2296_rdata));
  assign f2296_clk = clk;
  assign f2296_rst = rst;
  // Bindings to f2296

  // f2298
  logic [0:0] f2298_wen;
  logic [31:0] f2298_wdata;
  logic [0:0] f2298_clk;
  logic [0:0] f2298_rst;
  logic [31:0] f2298_rdata;
  sr_buffer_32_1 f2298(.wen(f2298_wen), .wdata(f2298_wdata), .clk(f2298_clk), .rst(f2298_rst), .rdata(f2298_rdata));
  assign f2298_clk = clk;
  assign f2298_rst = rst;
  // Bindings to f2298

  // f2300
  logic [0:0] f2300_wen;
  logic [31:0] f2300_wdata;
  logic [0:0] f2300_clk;
  logic [0:0] f2300_rst;
  logic [31:0] f2300_rdata;
  sr_buffer_32_1 f2300(.wen(f2300_wen), .wdata(f2300_wdata), .clk(f2300_clk), .rst(f2300_rst), .rdata(f2300_rdata));
  assign f2300_clk = clk;
  assign f2300_rst = rst;
  // Bindings to f2300

  // f2302
  logic [0:0] f2302_wen;
  logic [31:0] f2302_wdata;
  logic [0:0] f2302_clk;
  logic [0:0] f2302_rst;
  logic [31:0] f2302_rdata;
  sr_buffer_32_1 f2302(.wen(f2302_wen), .wdata(f2302_wdata), .clk(f2302_clk), .rst(f2302_rst), .rdata(f2302_rdata));
  assign f2302_clk = clk;
  assign f2302_rst = rst;
  // Bindings to f2302

  // f2304
  logic [0:0] f2304_wen;
  logic [31:0] f2304_wdata;
  logic [0:0] f2304_clk;
  logic [0:0] f2304_rst;
  logic [31:0] f2304_rdata;
  sr_buffer_32_1 f2304(.wen(f2304_wen), .wdata(f2304_wdata), .clk(f2304_clk), .rst(f2304_rst), .rdata(f2304_rdata));
  assign f2304_clk = clk;
  assign f2304_rst = rst;
  // Bindings to f2304

  // f2306
  logic [0:0] f2306_wen;
  logic [31:0] f2306_wdata;
  logic [0:0] f2306_clk;
  logic [0:0] f2306_rst;
  logic [31:0] f2306_rdata;
  sr_buffer_32_1 f2306(.wen(f2306_wen), .wdata(f2306_wdata), .clk(f2306_clk), .rst(f2306_rst), .rdata(f2306_rdata));
  assign f2306_clk = clk;
  assign f2306_rst = rst;
  // Bindings to f2306

  // f2308
  logic [0:0] f2308_wen;
  logic [31:0] f2308_wdata;
  logic [0:0] f2308_clk;
  logic [0:0] f2308_rst;
  logic [31:0] f2308_rdata;
  sr_buffer_32_1 f2308(.wen(f2308_wen), .wdata(f2308_wdata), .clk(f2308_clk), .rst(f2308_rst), .rdata(f2308_rdata));
  assign f2308_clk = clk;
  assign f2308_rst = rst;
  // Bindings to f2308

  // f2310
  logic [0:0] f2310_wen;
  logic [31:0] f2310_wdata;
  logic [0:0] f2310_clk;
  logic [0:0] f2310_rst;
  logic [31:0] f2310_rdata;
  sr_buffer_32_1 f2310(.wen(f2310_wen), .wdata(f2310_wdata), .clk(f2310_clk), .rst(f2310_rst), .rdata(f2310_rdata));
  assign f2310_clk = clk;
  assign f2310_rst = rst;
  // Bindings to f2310

  // f2312
  logic [0:0] f2312_wen;
  logic [31:0] f2312_wdata;
  logic [0:0] f2312_clk;
  logic [0:0] f2312_rst;
  logic [31:0] f2312_rdata;
  sr_buffer_32_1 f2312(.wen(f2312_wen), .wdata(f2312_wdata), .clk(f2312_clk), .rst(f2312_rst), .rdata(f2312_rdata));
  assign f2312_clk = clk;
  assign f2312_rst = rst;
  // Bindings to f2312

  // f2314
  logic [0:0] f2314_wen;
  logic [31:0] f2314_wdata;
  logic [0:0] f2314_clk;
  logic [0:0] f2314_rst;
  logic [31:0] f2314_rdata;
  sr_buffer_32_1 f2314(.wen(f2314_wen), .wdata(f2314_wdata), .clk(f2314_clk), .rst(f2314_rst), .rdata(f2314_rdata));
  assign f2314_clk = clk;
  assign f2314_rst = rst;
  // Bindings to f2314

  // f2316
  logic [0:0] f2316_wen;
  logic [31:0] f2316_wdata;
  logic [0:0] f2316_clk;
  logic [0:0] f2316_rst;
  logic [31:0] f2316_rdata;
  sr_buffer_32_1 f2316(.wen(f2316_wen), .wdata(f2316_wdata), .clk(f2316_clk), .rst(f2316_rst), .rdata(f2316_rdata));
  assign f2316_clk = clk;
  assign f2316_rst = rst;
  // Bindings to f2316

  // f2318
  logic [0:0] f2318_wen;
  logic [31:0] f2318_wdata;
  logic [0:0] f2318_clk;
  logic [0:0] f2318_rst;
  logic [31:0] f2318_rdata;
  sr_buffer_32_1 f2318(.wen(f2318_wen), .wdata(f2318_wdata), .clk(f2318_clk), .rst(f2318_rst), .rdata(f2318_rdata));
  assign f2318_clk = clk;
  assign f2318_rst = rst;
  // Bindings to f2318

  // f2320
  logic [0:0] f2320_wen;
  logic [31:0] f2320_wdata;
  logic [0:0] f2320_clk;
  logic [0:0] f2320_rst;
  logic [31:0] f2320_rdata;
  sr_buffer_32_1 f2320(.wen(f2320_wen), .wdata(f2320_wdata), .clk(f2320_clk), .rst(f2320_rst), .rdata(f2320_rdata));
  assign f2320_clk = clk;
  assign f2320_rst = rst;
  // Bindings to f2320

  // f2322
  logic [0:0] f2322_wen;
  logic [31:0] f2322_wdata;
  logic [0:0] f2322_clk;
  logic [0:0] f2322_rst;
  logic [31:0] f2322_rdata;
  sr_buffer_32_1 f2322(.wen(f2322_wen), .wdata(f2322_wdata), .clk(f2322_clk), .rst(f2322_rst), .rdata(f2322_rdata));
  assign f2322_clk = clk;
  assign f2322_rst = rst;
  // Bindings to f2322

  // f2324
  logic [0:0] f2324_wen;
  logic [31:0] f2324_wdata;
  logic [0:0] f2324_clk;
  logic [0:0] f2324_rst;
  logic [31:0] f2324_rdata;
  sr_buffer_32_1 f2324(.wen(f2324_wen), .wdata(f2324_wdata), .clk(f2324_clk), .rst(f2324_rst), .rdata(f2324_rdata));
  assign f2324_clk = clk;
  assign f2324_rst = rst;
  // Bindings to f2324

  // f2326
  logic [0:0] f2326_wen;
  logic [31:0] f2326_wdata;
  logic [0:0] f2326_clk;
  logic [0:0] f2326_rst;
  logic [31:0] f2326_rdata;
  sr_buffer_32_1 f2326(.wen(f2326_wen), .wdata(f2326_wdata), .clk(f2326_clk), .rst(f2326_rst), .rdata(f2326_rdata));
  assign f2326_clk = clk;
  assign f2326_rst = rst;
  // Bindings to f2326

  // f2328
  logic [0:0] f2328_wen;
  logic [31:0] f2328_wdata;
  logic [0:0] f2328_clk;
  logic [0:0] f2328_rst;
  logic [31:0] f2328_rdata;
  sr_buffer_32_1 f2328(.wen(f2328_wen), .wdata(f2328_wdata), .clk(f2328_clk), .rst(f2328_rst), .rdata(f2328_rdata));
  assign f2328_clk = clk;
  assign f2328_rst = rst;
  // Bindings to f2328

  // f2330
  logic [0:0] f2330_wen;
  logic [31:0] f2330_wdata;
  logic [0:0] f2330_clk;
  logic [0:0] f2330_rst;
  logic [31:0] f2330_rdata;
  sr_buffer_32_1 f2330(.wen(f2330_wen), .wdata(f2330_wdata), .clk(f2330_clk), .rst(f2330_rst), .rdata(f2330_rdata));
  assign f2330_clk = clk;
  assign f2330_rst = rst;
  // Bindings to f2330

  // f2332
  logic [0:0] f2332_wen;
  logic [31:0] f2332_wdata;
  logic [0:0] f2332_clk;
  logic [0:0] f2332_rst;
  logic [31:0] f2332_rdata;
  sr_buffer_32_1 f2332(.wen(f2332_wen), .wdata(f2332_wdata), .clk(f2332_clk), .rst(f2332_rst), .rdata(f2332_rdata));
  assign f2332_clk = clk;
  assign f2332_rst = rst;
  // Bindings to f2332

  // f2334
  logic [0:0] f2334_wen;
  logic [31:0] f2334_wdata;
  logic [0:0] f2334_clk;
  logic [0:0] f2334_rst;
  logic [31:0] f2334_rdata;
  sr_buffer_32_1 f2334(.wen(f2334_wen), .wdata(f2334_wdata), .clk(f2334_clk), .rst(f2334_rst), .rdata(f2334_rdata));
  assign f2334_clk = clk;
  assign f2334_rst = rst;
  // Bindings to f2334

  // f2336
  logic [0:0] f2336_wen;
  logic [31:0] f2336_wdata;
  logic [0:0] f2336_clk;
  logic [0:0] f2336_rst;
  logic [31:0] f2336_rdata;
  sr_buffer_32_1 f2336(.wen(f2336_wen), .wdata(f2336_wdata), .clk(f2336_clk), .rst(f2336_rst), .rdata(f2336_rdata));
  assign f2336_clk = clk;
  assign f2336_rst = rst;
  // Bindings to f2336

  // f2338
  logic [0:0] f2338_wen;
  logic [31:0] f2338_wdata;
  logic [0:0] f2338_clk;
  logic [0:0] f2338_rst;
  logic [31:0] f2338_rdata;
  sr_buffer_32_1 f2338(.wen(f2338_wen), .wdata(f2338_wdata), .clk(f2338_clk), .rst(f2338_rst), .rdata(f2338_rdata));
  assign f2338_clk = clk;
  assign f2338_rst = rst;
  // Bindings to f2338

  // f2340
  logic [0:0] f2340_wen;
  logic [31:0] f2340_wdata;
  logic [0:0] f2340_clk;
  logic [0:0] f2340_rst;
  logic [31:0] f2340_rdata;
  sr_buffer_32_1 f2340(.wen(f2340_wen), .wdata(f2340_wdata), .clk(f2340_clk), .rst(f2340_rst), .rdata(f2340_rdata));
  assign f2340_clk = clk;
  assign f2340_rst = rst;
  // Bindings to f2340

  // f2342
  logic [0:0] f2342_wen;
  logic [31:0] f2342_wdata;
  logic [0:0] f2342_clk;
  logic [0:0] f2342_rst;
  logic [31:0] f2342_rdata;
  sr_buffer_32_1 f2342(.wen(f2342_wen), .wdata(f2342_wdata), .clk(f2342_clk), .rst(f2342_rst), .rdata(f2342_rdata));
  assign f2342_clk = clk;
  assign f2342_rst = rst;
  // Bindings to f2342

  // f2344
  logic [0:0] f2344_wen;
  logic [31:0] f2344_wdata;
  logic [0:0] f2344_clk;
  logic [0:0] f2344_rst;
  logic [31:0] f2344_rdata;
  sr_buffer_32_1 f2344(.wen(f2344_wen), .wdata(f2344_wdata), .clk(f2344_clk), .rst(f2344_rst), .rdata(f2344_rdata));
  assign f2344_clk = clk;
  assign f2344_rst = rst;
  // Bindings to f2344

  // f2346
  logic [0:0] f2346_wen;
  logic [31:0] f2346_wdata;
  logic [0:0] f2346_clk;
  logic [0:0] f2346_rst;
  logic [31:0] f2346_rdata;
  sr_buffer_32_1 f2346(.wen(f2346_wen), .wdata(f2346_wdata), .clk(f2346_clk), .rst(f2346_rst), .rdata(f2346_rdata));
  assign f2346_clk = clk;
  assign f2346_rst = rst;
  // Bindings to f2346

  // f2348
  logic [0:0] f2348_wen;
  logic [31:0] f2348_wdata;
  logic [0:0] f2348_clk;
  logic [0:0] f2348_rst;
  logic [31:0] f2348_rdata;
  sr_buffer_32_1 f2348(.wen(f2348_wen), .wdata(f2348_wdata), .clk(f2348_clk), .rst(f2348_rst), .rdata(f2348_rdata));
  assign f2348_clk = clk;
  assign f2348_rst = rst;
  // Bindings to f2348

  // f2350
  logic [0:0] f2350_wen;
  logic [31:0] f2350_wdata;
  logic [0:0] f2350_clk;
  logic [0:0] f2350_rst;
  logic [31:0] f2350_rdata;
  sr_buffer_32_1 f2350(.wen(f2350_wen), .wdata(f2350_wdata), .clk(f2350_clk), .rst(f2350_rst), .rdata(f2350_rdata));
  assign f2350_clk = clk;
  assign f2350_rst = rst;
  // Bindings to f2350

  // f2352
  logic [0:0] f2352_wen;
  logic [31:0] f2352_wdata;
  logic [0:0] f2352_clk;
  logic [0:0] f2352_rst;
  logic [31:0] f2352_rdata;
  sr_buffer_32_1 f2352(.wen(f2352_wen), .wdata(f2352_wdata), .clk(f2352_clk), .rst(f2352_rst), .rdata(f2352_rdata));
  assign f2352_clk = clk;
  assign f2352_rst = rst;
  // Bindings to f2352

  // f2354
  logic [0:0] f2354_wen;
  logic [31:0] f2354_wdata;
  logic [0:0] f2354_clk;
  logic [0:0] f2354_rst;
  logic [31:0] f2354_rdata;
  sr_buffer_32_1 f2354(.wen(f2354_wen), .wdata(f2354_wdata), .clk(f2354_clk), .rst(f2354_rst), .rdata(f2354_rdata));
  assign f2354_clk = clk;
  assign f2354_rst = rst;
  // Bindings to f2354

  // f2356
  logic [0:0] f2356_wen;
  logic [31:0] f2356_wdata;
  logic [0:0] f2356_clk;
  logic [0:0] f2356_rst;
  logic [31:0] f2356_rdata;
  sr_buffer_32_1 f2356(.wen(f2356_wen), .wdata(f2356_wdata), .clk(f2356_clk), .rst(f2356_rst), .rdata(f2356_rdata));
  assign f2356_clk = clk;
  assign f2356_rst = rst;
  // Bindings to f2356

  // f2358
  logic [0:0] f2358_wen;
  logic [31:0] f2358_wdata;
  logic [0:0] f2358_clk;
  logic [0:0] f2358_rst;
  logic [31:0] f2358_rdata;
  sr_buffer_32_1 f2358(.wen(f2358_wen), .wdata(f2358_wdata), .clk(f2358_clk), .rst(f2358_rst), .rdata(f2358_rdata));
  assign f2358_clk = clk;
  assign f2358_rst = rst;
  // Bindings to f2358

  // f2360
  logic [0:0] f2360_wen;
  logic [31:0] f2360_wdata;
  logic [0:0] f2360_clk;
  logic [0:0] f2360_rst;
  logic [31:0] f2360_rdata;
  sr_buffer_32_1 f2360(.wen(f2360_wen), .wdata(f2360_wdata), .clk(f2360_clk), .rst(f2360_rst), .rdata(f2360_rdata));
  assign f2360_clk = clk;
  assign f2360_rst = rst;
  // Bindings to f2360

  // f2362
  logic [0:0] f2362_wen;
  logic [31:0] f2362_wdata;
  logic [0:0] f2362_clk;
  logic [0:0] f2362_rst;
  logic [31:0] f2362_rdata;
  sr_buffer_32_1 f2362(.wen(f2362_wen), .wdata(f2362_wdata), .clk(f2362_clk), .rst(f2362_rst), .rdata(f2362_rdata));
  assign f2362_clk = clk;
  assign f2362_rst = rst;
  // Bindings to f2362

  // f2364
  logic [0:0] f2364_wen;
  logic [31:0] f2364_wdata;
  logic [0:0] f2364_clk;
  logic [0:0] f2364_rst;
  logic [31:0] f2364_rdata;
  sr_buffer_32_1 f2364(.wen(f2364_wen), .wdata(f2364_wdata), .clk(f2364_clk), .rst(f2364_rst), .rdata(f2364_rdata));
  assign f2364_clk = clk;
  assign f2364_rst = rst;
  // Bindings to f2364

  // f2366
  logic [0:0] f2366_wen;
  logic [31:0] f2366_wdata;
  logic [0:0] f2366_clk;
  logic [0:0] f2366_rst;
  logic [31:0] f2366_rdata;
  sr_buffer_32_1 f2366(.wen(f2366_wen), .wdata(f2366_wdata), .clk(f2366_clk), .rst(f2366_rst), .rdata(f2366_rdata));
  assign f2366_clk = clk;
  assign f2366_rst = rst;
  // Bindings to f2366

  // f2368
  logic [0:0] f2368_wen;
  logic [31:0] f2368_wdata;
  logic [0:0] f2368_clk;
  logic [0:0] f2368_rst;
  logic [31:0] f2368_rdata;
  sr_buffer_32_1 f2368(.wen(f2368_wen), .wdata(f2368_wdata), .clk(f2368_clk), .rst(f2368_rst), .rdata(f2368_rdata));
  assign f2368_clk = clk;
  assign f2368_rst = rst;
  // Bindings to f2368

  // f2370
  logic [0:0] f2370_wen;
  logic [31:0] f2370_wdata;
  logic [0:0] f2370_clk;
  logic [0:0] f2370_rst;
  logic [31:0] f2370_rdata;
  sr_buffer_32_1 f2370(.wen(f2370_wen), .wdata(f2370_wdata), .clk(f2370_clk), .rst(f2370_rst), .rdata(f2370_rdata));
  assign f2370_clk = clk;
  assign f2370_rst = rst;
  // Bindings to f2370

  // f2372
  logic [0:0] f2372_wen;
  logic [31:0] f2372_wdata;
  logic [0:0] f2372_clk;
  logic [0:0] f2372_rst;
  logic [31:0] f2372_rdata;
  sr_buffer_32_1 f2372(.wen(f2372_wen), .wdata(f2372_wdata), .clk(f2372_clk), .rst(f2372_rst), .rdata(f2372_rdata));
  assign f2372_clk = clk;
  assign f2372_rst = rst;
  // Bindings to f2372

  // f2374
  logic [0:0] f2374_wen;
  logic [31:0] f2374_wdata;
  logic [0:0] f2374_clk;
  logic [0:0] f2374_rst;
  logic [31:0] f2374_rdata;
  sr_buffer_32_1 f2374(.wen(f2374_wen), .wdata(f2374_wdata), .clk(f2374_clk), .rst(f2374_rst), .rdata(f2374_rdata));
  assign f2374_clk = clk;
  assign f2374_rst = rst;
  // Bindings to f2374

  // f2376
  logic [0:0] f2376_wen;
  logic [31:0] f2376_wdata;
  logic [0:0] f2376_clk;
  logic [0:0] f2376_rst;
  logic [31:0] f2376_rdata;
  sr_buffer_32_1 f2376(.wen(f2376_wen), .wdata(f2376_wdata), .clk(f2376_clk), .rst(f2376_rst), .rdata(f2376_rdata));
  assign f2376_clk = clk;
  assign f2376_rst = rst;
  // Bindings to f2376

  // f2378
  logic [0:0] f2378_wen;
  logic [31:0] f2378_wdata;
  logic [0:0] f2378_clk;
  logic [0:0] f2378_rst;
  logic [31:0] f2378_rdata;
  sr_buffer_32_1 f2378(.wen(f2378_wen), .wdata(f2378_wdata), .clk(f2378_clk), .rst(f2378_rst), .rdata(f2378_rdata));
  assign f2378_clk = clk;
  assign f2378_rst = rst;
  // Bindings to f2378

  // f2380
  logic [0:0] f2380_wen;
  logic [31:0] f2380_wdata;
  logic [0:0] f2380_clk;
  logic [0:0] f2380_rst;
  logic [31:0] f2380_rdata;
  sr_buffer_32_1 f2380(.wen(f2380_wen), .wdata(f2380_wdata), .clk(f2380_clk), .rst(f2380_rst), .rdata(f2380_rdata));
  assign f2380_clk = clk;
  assign f2380_rst = rst;
  // Bindings to f2380

  // f2382
  logic [0:0] f2382_wen;
  logic [31:0] f2382_wdata;
  logic [0:0] f2382_clk;
  logic [0:0] f2382_rst;
  logic [31:0] f2382_rdata;
  sr_buffer_32_1 f2382(.wen(f2382_wen), .wdata(f2382_wdata), .clk(f2382_clk), .rst(f2382_rst), .rdata(f2382_rdata));
  assign f2382_clk = clk;
  assign f2382_rst = rst;
  // Bindings to f2382

  // f2384
  logic [0:0] f2384_wen;
  logic [31:0] f2384_wdata;
  logic [0:0] f2384_clk;
  logic [0:0] f2384_rst;
  logic [31:0] f2384_rdata;
  sr_buffer_32_1 f2384(.wen(f2384_wen), .wdata(f2384_wdata), .clk(f2384_clk), .rst(f2384_rst), .rdata(f2384_rdata));
  assign f2384_clk = clk;
  assign f2384_rst = rst;
  // Bindings to f2384

  // f2386
  logic [0:0] f2386_wen;
  logic [31:0] f2386_wdata;
  logic [0:0] f2386_clk;
  logic [0:0] f2386_rst;
  logic [31:0] f2386_rdata;
  sr_buffer_32_1 f2386(.wen(f2386_wen), .wdata(f2386_wdata), .clk(f2386_clk), .rst(f2386_rst), .rdata(f2386_rdata));
  assign f2386_clk = clk;
  assign f2386_rst = rst;
  // Bindings to f2386

  // f2388
  logic [0:0] f2388_wen;
  logic [31:0] f2388_wdata;
  logic [0:0] f2388_clk;
  logic [0:0] f2388_rst;
  logic [31:0] f2388_rdata;
  sr_buffer_32_1 f2388(.wen(f2388_wen), .wdata(f2388_wdata), .clk(f2388_clk), .rst(f2388_rst), .rdata(f2388_rdata));
  assign f2388_clk = clk;
  assign f2388_rst = rst;
  // Bindings to f2388

  // f2390
  logic [0:0] f2390_wen;
  logic [31:0] f2390_wdata;
  logic [0:0] f2390_clk;
  logic [0:0] f2390_rst;
  logic [31:0] f2390_rdata;
  sr_buffer_32_1 f2390(.wen(f2390_wen), .wdata(f2390_wdata), .clk(f2390_clk), .rst(f2390_rst), .rdata(f2390_rdata));
  assign f2390_clk = clk;
  assign f2390_rst = rst;
  // Bindings to f2390

  // f2392
  logic [0:0] f2392_wen;
  logic [31:0] f2392_wdata;
  logic [0:0] f2392_clk;
  logic [0:0] f2392_rst;
  logic [31:0] f2392_rdata;
  sr_buffer_32_1 f2392(.wen(f2392_wen), .wdata(f2392_wdata), .clk(f2392_clk), .rst(f2392_rst), .rdata(f2392_rdata));
  assign f2392_clk = clk;
  assign f2392_rst = rst;
  // Bindings to f2392

  // f2394
  logic [0:0] f2394_wen;
  logic [31:0] f2394_wdata;
  logic [0:0] f2394_clk;
  logic [0:0] f2394_rst;
  logic [31:0] f2394_rdata;
  sr_buffer_32_1 f2394(.wen(f2394_wen), .wdata(f2394_wdata), .clk(f2394_clk), .rst(f2394_rst), .rdata(f2394_rdata));
  assign f2394_clk = clk;
  assign f2394_rst = rst;
  // Bindings to f2394

  // f2396
  logic [0:0] f2396_wen;
  logic [31:0] f2396_wdata;
  logic [0:0] f2396_clk;
  logic [0:0] f2396_rst;
  logic [31:0] f2396_rdata;
  sr_buffer_32_1 f2396(.wen(f2396_wen), .wdata(f2396_wdata), .clk(f2396_clk), .rst(f2396_rst), .rdata(f2396_rdata));
  assign f2396_clk = clk;
  assign f2396_rst = rst;
  // Bindings to f2396

  // f2398
  logic [0:0] f2398_wen;
  logic [31:0] f2398_wdata;
  logic [0:0] f2398_clk;
  logic [0:0] f2398_rst;
  logic [31:0] f2398_rdata;
  sr_buffer_32_1 f2398(.wen(f2398_wen), .wdata(f2398_wdata), .clk(f2398_clk), .rst(f2398_rst), .rdata(f2398_rdata));
  assign f2398_clk = clk;
  assign f2398_rst = rst;
  // Bindings to f2398

  // f2400
  logic [0:0] f2400_wen;
  logic [31:0] f2400_wdata;
  logic [0:0] f2400_clk;
  logic [0:0] f2400_rst;
  logic [31:0] f2400_rdata;
  sr_buffer_32_1 f2400(.wen(f2400_wen), .wdata(f2400_wdata), .clk(f2400_clk), .rst(f2400_rst), .rdata(f2400_rdata));
  assign f2400_clk = clk;
  assign f2400_rst = rst;
  // Bindings to f2400

  // f2402
  logic [0:0] f2402_wen;
  logic [31:0] f2402_wdata;
  logic [0:0] f2402_clk;
  logic [0:0] f2402_rst;
  logic [31:0] f2402_rdata;
  sr_buffer_32_1 f2402(.wen(f2402_wen), .wdata(f2402_wdata), .clk(f2402_clk), .rst(f2402_rst), .rdata(f2402_rdata));
  assign f2402_clk = clk;
  assign f2402_rst = rst;
  // Bindings to f2402

  // f2404
  logic [0:0] f2404_wen;
  logic [31:0] f2404_wdata;
  logic [0:0] f2404_clk;
  logic [0:0] f2404_rst;
  logic [31:0] f2404_rdata;
  sr_buffer_32_1 f2404(.wen(f2404_wen), .wdata(f2404_wdata), .clk(f2404_clk), .rst(f2404_rst), .rdata(f2404_rdata));
  assign f2404_clk = clk;
  assign f2404_rst = rst;
  // Bindings to f2404

  // f2406
  logic [0:0] f2406_wen;
  logic [31:0] f2406_wdata;
  logic [0:0] f2406_clk;
  logic [0:0] f2406_rst;
  logic [31:0] f2406_rdata;
  sr_buffer_32_1 f2406(.wen(f2406_wen), .wdata(f2406_wdata), .clk(f2406_clk), .rst(f2406_rst), .rdata(f2406_rdata));
  assign f2406_clk = clk;
  assign f2406_rst = rst;
  // Bindings to f2406

  // f2408
  logic [0:0] f2408_wen;
  logic [31:0] f2408_wdata;
  logic [0:0] f2408_clk;
  logic [0:0] f2408_rst;
  logic [31:0] f2408_rdata;
  sr_buffer_32_1 f2408(.wen(f2408_wen), .wdata(f2408_wdata), .clk(f2408_clk), .rst(f2408_rst), .rdata(f2408_rdata));
  assign f2408_clk = clk;
  assign f2408_rst = rst;
  // Bindings to f2408

  // f2410
  logic [0:0] f2410_wen;
  logic [31:0] f2410_wdata;
  logic [0:0] f2410_clk;
  logic [0:0] f2410_rst;
  logic [31:0] f2410_rdata;
  sr_buffer_32_1 f2410(.wen(f2410_wen), .wdata(f2410_wdata), .clk(f2410_clk), .rst(f2410_rst), .rdata(f2410_rdata));
  assign f2410_clk = clk;
  assign f2410_rst = rst;
  // Bindings to f2410

  // f2412
  logic [0:0] f2412_wen;
  logic [31:0] f2412_wdata;
  logic [0:0] f2412_clk;
  logic [0:0] f2412_rst;
  logic [31:0] f2412_rdata;
  sr_buffer_32_1 f2412(.wen(f2412_wen), .wdata(f2412_wdata), .clk(f2412_clk), .rst(f2412_rst), .rdata(f2412_rdata));
  assign f2412_clk = clk;
  assign f2412_rst = rst;
  // Bindings to f2412

  // f2414
  logic [0:0] f2414_wen;
  logic [31:0] f2414_wdata;
  logic [0:0] f2414_clk;
  logic [0:0] f2414_rst;
  logic [31:0] f2414_rdata;
  sr_buffer_32_1 f2414(.wen(f2414_wen), .wdata(f2414_wdata), .clk(f2414_clk), .rst(f2414_rst), .rdata(f2414_rdata));
  assign f2414_clk = clk;
  assign f2414_rst = rst;
  // Bindings to f2414

  // f2416
  logic [0:0] f2416_wen;
  logic [31:0] f2416_wdata;
  logic [0:0] f2416_clk;
  logic [0:0] f2416_rst;
  logic [31:0] f2416_rdata;
  sr_buffer_32_1 f2416(.wen(f2416_wen), .wdata(f2416_wdata), .clk(f2416_clk), .rst(f2416_rst), .rdata(f2416_rdata));
  assign f2416_clk = clk;
  assign f2416_rst = rst;
  // Bindings to f2416

  // f2418
  logic [0:0] f2418_wen;
  logic [31:0] f2418_wdata;
  logic [0:0] f2418_clk;
  logic [0:0] f2418_rst;
  logic [31:0] f2418_rdata;
  sr_buffer_32_1 f2418(.wen(f2418_wen), .wdata(f2418_wdata), .clk(f2418_clk), .rst(f2418_rst), .rdata(f2418_rdata));
  assign f2418_clk = clk;
  assign f2418_rst = rst;
  // Bindings to f2418

  // f2420
  logic [0:0] f2420_wen;
  logic [31:0] f2420_wdata;
  logic [0:0] f2420_clk;
  logic [0:0] f2420_rst;
  logic [31:0] f2420_rdata;
  sr_buffer_32_1 f2420(.wen(f2420_wen), .wdata(f2420_wdata), .clk(f2420_clk), .rst(f2420_rst), .rdata(f2420_rdata));
  assign f2420_clk = clk;
  assign f2420_rst = rst;
  // Bindings to f2420

  // f2422
  logic [0:0] f2422_wen;
  logic [31:0] f2422_wdata;
  logic [0:0] f2422_clk;
  logic [0:0] f2422_rst;
  logic [31:0] f2422_rdata;
  sr_buffer_32_1 f2422(.wen(f2422_wen), .wdata(f2422_wdata), .clk(f2422_clk), .rst(f2422_rst), .rdata(f2422_rdata));
  assign f2422_clk = clk;
  assign f2422_rst = rst;
  // Bindings to f2422

  // f2424
  logic [0:0] f2424_wen;
  logic [31:0] f2424_wdata;
  logic [0:0] f2424_clk;
  logic [0:0] f2424_rst;
  logic [31:0] f2424_rdata;
  sr_buffer_32_1 f2424(.wen(f2424_wen), .wdata(f2424_wdata), .clk(f2424_clk), .rst(f2424_rst), .rdata(f2424_rdata));
  assign f2424_clk = clk;
  assign f2424_rst = rst;
  // Bindings to f2424

  // f2426
  logic [0:0] f2426_wen;
  logic [31:0] f2426_wdata;
  logic [0:0] f2426_clk;
  logic [0:0] f2426_rst;
  logic [31:0] f2426_rdata;
  sr_buffer_32_1 f2426(.wen(f2426_wen), .wdata(f2426_wdata), .clk(f2426_clk), .rst(f2426_rst), .rdata(f2426_rdata));
  assign f2426_clk = clk;
  assign f2426_rst = rst;
  // Bindings to f2426

  // f2428
  logic [0:0] f2428_wen;
  logic [31:0] f2428_wdata;
  logic [0:0] f2428_clk;
  logic [0:0] f2428_rst;
  logic [31:0] f2428_rdata;
  sr_buffer_32_1 f2428(.wen(f2428_wen), .wdata(f2428_wdata), .clk(f2428_clk), .rst(f2428_rst), .rdata(f2428_rdata));
  assign f2428_clk = clk;
  assign f2428_rst = rst;
  // Bindings to f2428

  // f2430
  logic [0:0] f2430_wen;
  logic [31:0] f2430_wdata;
  logic [0:0] f2430_clk;
  logic [0:0] f2430_rst;
  logic [31:0] f2430_rdata;
  sr_buffer_32_1 f2430(.wen(f2430_wen), .wdata(f2430_wdata), .clk(f2430_clk), .rst(f2430_rst), .rdata(f2430_rdata));
  assign f2430_clk = clk;
  assign f2430_rst = rst;
  // Bindings to f2430

  // f2432
  logic [0:0] f2432_wen;
  logic [31:0] f2432_wdata;
  logic [0:0] f2432_clk;
  logic [0:0] f2432_rst;
  logic [31:0] f2432_rdata;
  sr_buffer_32_1 f2432(.wen(f2432_wen), .wdata(f2432_wdata), .clk(f2432_clk), .rst(f2432_rst), .rdata(f2432_rdata));
  assign f2432_clk = clk;
  assign f2432_rst = rst;
  // Bindings to f2432

  // f2434
  logic [0:0] f2434_wen;
  logic [31:0] f2434_wdata;
  logic [0:0] f2434_clk;
  logic [0:0] f2434_rst;
  logic [31:0] f2434_rdata;
  sr_buffer_32_1 f2434(.wen(f2434_wen), .wdata(f2434_wdata), .clk(f2434_clk), .rst(f2434_rst), .rdata(f2434_rdata));
  assign f2434_clk = clk;
  assign f2434_rst = rst;
  // Bindings to f2434

  // f2436
  logic [0:0] f2436_wen;
  logic [31:0] f2436_wdata;
  logic [0:0] f2436_clk;
  logic [0:0] f2436_rst;
  logic [31:0] f2436_rdata;
  sr_buffer_32_1 f2436(.wen(f2436_wen), .wdata(f2436_wdata), .clk(f2436_clk), .rst(f2436_rst), .rdata(f2436_rdata));
  assign f2436_clk = clk;
  assign f2436_rst = rst;
  // Bindings to f2436

  // f2438
  logic [0:0] f2438_wen;
  logic [31:0] f2438_wdata;
  logic [0:0] f2438_clk;
  logic [0:0] f2438_rst;
  logic [31:0] f2438_rdata;
  sr_buffer_32_1 f2438(.wen(f2438_wen), .wdata(f2438_wdata), .clk(f2438_clk), .rst(f2438_rst), .rdata(f2438_rdata));
  assign f2438_clk = clk;
  assign f2438_rst = rst;
  // Bindings to f2438

  // f2440
  logic [0:0] f2440_wen;
  logic [31:0] f2440_wdata;
  logic [0:0] f2440_clk;
  logic [0:0] f2440_rst;
  logic [31:0] f2440_rdata;
  sr_buffer_32_1 f2440(.wen(f2440_wen), .wdata(f2440_wdata), .clk(f2440_clk), .rst(f2440_rst), .rdata(f2440_rdata));
  assign f2440_clk = clk;
  assign f2440_rst = rst;
  // Bindings to f2440

  // f2442
  logic [0:0] f2442_wen;
  logic [31:0] f2442_wdata;
  logic [0:0] f2442_clk;
  logic [0:0] f2442_rst;
  logic [31:0] f2442_rdata;
  sr_buffer_32_1 f2442(.wen(f2442_wen), .wdata(f2442_wdata), .clk(f2442_clk), .rst(f2442_rst), .rdata(f2442_rdata));
  assign f2442_clk = clk;
  assign f2442_rst = rst;
  // Bindings to f2442

  // f2444
  logic [0:0] f2444_wen;
  logic [31:0] f2444_wdata;
  logic [0:0] f2444_clk;
  logic [0:0] f2444_rst;
  logic [31:0] f2444_rdata;
  sr_buffer_32_1 f2444(.wen(f2444_wen), .wdata(f2444_wdata), .clk(f2444_clk), .rst(f2444_rst), .rdata(f2444_rdata));
  assign f2444_clk = clk;
  assign f2444_rst = rst;
  // Bindings to f2444

  // f2446
  logic [0:0] f2446_wen;
  logic [31:0] f2446_wdata;
  logic [0:0] f2446_clk;
  logic [0:0] f2446_rst;
  logic [31:0] f2446_rdata;
  sr_buffer_32_1 f2446(.wen(f2446_wen), .wdata(f2446_wdata), .clk(f2446_clk), .rst(f2446_rst), .rdata(f2446_rdata));
  assign f2446_clk = clk;
  assign f2446_rst = rst;
  // Bindings to f2446

  // f2448
  logic [0:0] f2448_wen;
  logic [31:0] f2448_wdata;
  logic [0:0] f2448_clk;
  logic [0:0] f2448_rst;
  logic [31:0] f2448_rdata;
  sr_buffer_32_1 f2448(.wen(f2448_wen), .wdata(f2448_wdata), .clk(f2448_clk), .rst(f2448_rst), .rdata(f2448_rdata));
  assign f2448_clk = clk;
  assign f2448_rst = rst;
  // Bindings to f2448

  // f2450
  logic [0:0] f2450_wen;
  logic [31:0] f2450_wdata;
  logic [0:0] f2450_clk;
  logic [0:0] f2450_rst;
  logic [31:0] f2450_rdata;
  sr_buffer_32_1 f2450(.wen(f2450_wen), .wdata(f2450_wdata), .clk(f2450_clk), .rst(f2450_rst), .rdata(f2450_rdata));
  assign f2450_clk = clk;
  assign f2450_rst = rst;
  // Bindings to f2450

  // f2452
  logic [0:0] f2452_wen;
  logic [31:0] f2452_wdata;
  logic [0:0] f2452_clk;
  logic [0:0] f2452_rst;
  logic [31:0] f2452_rdata;
  sr_buffer_32_1 f2452(.wen(f2452_wen), .wdata(f2452_wdata), .clk(f2452_clk), .rst(f2452_rst), .rdata(f2452_rdata));
  assign f2452_clk = clk;
  assign f2452_rst = rst;
  // Bindings to f2452

  // f2454
  logic [0:0] f2454_wen;
  logic [31:0] f2454_wdata;
  logic [0:0] f2454_clk;
  logic [0:0] f2454_rst;
  logic [31:0] f2454_rdata;
  sr_buffer_32_1 f2454(.wen(f2454_wen), .wdata(f2454_wdata), .clk(f2454_clk), .rst(f2454_rst), .rdata(f2454_rdata));
  assign f2454_clk = clk;
  assign f2454_rst = rst;
  // Bindings to f2454

  // f2456
  logic [0:0] f2456_wen;
  logic [31:0] f2456_wdata;
  logic [0:0] f2456_clk;
  logic [0:0] f2456_rst;
  logic [31:0] f2456_rdata;
  sr_buffer_32_1 f2456(.wen(f2456_wen), .wdata(f2456_wdata), .clk(f2456_clk), .rst(f2456_rst), .rdata(f2456_rdata));
  assign f2456_clk = clk;
  assign f2456_rst = rst;
  // Bindings to f2456

  // f2458
  logic [0:0] f2458_wen;
  logic [31:0] f2458_wdata;
  logic [0:0] f2458_clk;
  logic [0:0] f2458_rst;
  logic [31:0] f2458_rdata;
  sr_buffer_32_1 f2458(.wen(f2458_wen), .wdata(f2458_wdata), .clk(f2458_clk), .rst(f2458_rst), .rdata(f2458_rdata));
  assign f2458_clk = clk;
  assign f2458_rst = rst;
  // Bindings to f2458

  // f2460
  logic [0:0] f2460_wen;
  logic [31:0] f2460_wdata;
  logic [0:0] f2460_clk;
  logic [0:0] f2460_rst;
  logic [31:0] f2460_rdata;
  sr_buffer_32_1 f2460(.wen(f2460_wen), .wdata(f2460_wdata), .clk(f2460_clk), .rst(f2460_rst), .rdata(f2460_rdata));
  assign f2460_clk = clk;
  assign f2460_rst = rst;
  // Bindings to f2460

  // f2462
  logic [0:0] f2462_wen;
  logic [31:0] f2462_wdata;
  logic [0:0] f2462_clk;
  logic [0:0] f2462_rst;
  logic [31:0] f2462_rdata;
  sr_buffer_32_1 f2462(.wen(f2462_wen), .wdata(f2462_wdata), .clk(f2462_clk), .rst(f2462_rst), .rdata(f2462_rdata));
  assign f2462_clk = clk;
  assign f2462_rst = rst;
  // Bindings to f2462

  // f2464
  logic [0:0] f2464_wen;
  logic [31:0] f2464_wdata;
  logic [0:0] f2464_clk;
  logic [0:0] f2464_rst;
  logic [31:0] f2464_rdata;
  sr_buffer_32_1 f2464(.wen(f2464_wen), .wdata(f2464_wdata), .clk(f2464_clk), .rst(f2464_rst), .rdata(f2464_rdata));
  assign f2464_clk = clk;
  assign f2464_rst = rst;
  // Bindings to f2464

  // f2466
  logic [0:0] f2466_wen;
  logic [31:0] f2466_wdata;
  logic [0:0] f2466_clk;
  logic [0:0] f2466_rst;
  logic [31:0] f2466_rdata;
  sr_buffer_32_1 f2466(.wen(f2466_wen), .wdata(f2466_wdata), .clk(f2466_clk), .rst(f2466_rst), .rdata(f2466_rdata));
  assign f2466_clk = clk;
  assign f2466_rst = rst;
  // Bindings to f2466

  // f2468
  logic [0:0] f2468_wen;
  logic [31:0] f2468_wdata;
  logic [0:0] f2468_clk;
  logic [0:0] f2468_rst;
  logic [31:0] f2468_rdata;
  sr_buffer_32_1 f2468(.wen(f2468_wen), .wdata(f2468_wdata), .clk(f2468_clk), .rst(f2468_rst), .rdata(f2468_rdata));
  assign f2468_clk = clk;
  assign f2468_rst = rst;
  // Bindings to f2468

  // f2470
  logic [0:0] f2470_wen;
  logic [31:0] f2470_wdata;
  logic [0:0] f2470_clk;
  logic [0:0] f2470_rst;
  logic [31:0] f2470_rdata;
  sr_buffer_32_1 f2470(.wen(f2470_wen), .wdata(f2470_wdata), .clk(f2470_clk), .rst(f2470_rst), .rdata(f2470_rdata));
  assign f2470_clk = clk;
  assign f2470_rst = rst;
  // Bindings to f2470

  // f2472
  logic [0:0] f2472_wen;
  logic [31:0] f2472_wdata;
  logic [0:0] f2472_clk;
  logic [0:0] f2472_rst;
  logic [31:0] f2472_rdata;
  sr_buffer_32_1 f2472(.wen(f2472_wen), .wdata(f2472_wdata), .clk(f2472_clk), .rst(f2472_rst), .rdata(f2472_rdata));
  assign f2472_clk = clk;
  assign f2472_rst = rst;
  // Bindings to f2472

  // f2474
  logic [0:0] f2474_wen;
  logic [31:0] f2474_wdata;
  logic [0:0] f2474_clk;
  logic [0:0] f2474_rst;
  logic [31:0] f2474_rdata;
  sr_buffer_32_1 f2474(.wen(f2474_wen), .wdata(f2474_wdata), .clk(f2474_clk), .rst(f2474_rst), .rdata(f2474_rdata));
  assign f2474_clk = clk;
  assign f2474_rst = rst;
  // Bindings to f2474

  // f2476
  logic [0:0] f2476_wen;
  logic [31:0] f2476_wdata;
  logic [0:0] f2476_clk;
  logic [0:0] f2476_rst;
  logic [31:0] f2476_rdata;
  sr_buffer_32_1 f2476(.wen(f2476_wen), .wdata(f2476_wdata), .clk(f2476_clk), .rst(f2476_rst), .rdata(f2476_rdata));
  assign f2476_clk = clk;
  assign f2476_rst = rst;
  // Bindings to f2476

  // f2478
  logic [0:0] f2478_wen;
  logic [31:0] f2478_wdata;
  logic [0:0] f2478_clk;
  logic [0:0] f2478_rst;
  logic [31:0] f2478_rdata;
  sr_buffer_32_1 f2478(.wen(f2478_wen), .wdata(f2478_wdata), .clk(f2478_clk), .rst(f2478_rst), .rdata(f2478_rdata));
  assign f2478_clk = clk;
  assign f2478_rst = rst;
  // Bindings to f2478

  // f2480
  logic [0:0] f2480_wen;
  logic [31:0] f2480_wdata;
  logic [0:0] f2480_clk;
  logic [0:0] f2480_rst;
  logic [31:0] f2480_rdata;
  sr_buffer_32_1 f2480(.wen(f2480_wen), .wdata(f2480_wdata), .clk(f2480_clk), .rst(f2480_rst), .rdata(f2480_rdata));
  assign f2480_clk = clk;
  assign f2480_rst = rst;
  // Bindings to f2480

  // f2482
  logic [0:0] f2482_wen;
  logic [31:0] f2482_wdata;
  logic [0:0] f2482_clk;
  logic [0:0] f2482_rst;
  logic [31:0] f2482_rdata;
  sr_buffer_32_1 f2482(.wen(f2482_wen), .wdata(f2482_wdata), .clk(f2482_clk), .rst(f2482_rst), .rdata(f2482_rdata));
  assign f2482_clk = clk;
  assign f2482_rst = rst;
  // Bindings to f2482

  // f2484
  logic [0:0] f2484_wen;
  logic [31:0] f2484_wdata;
  logic [0:0] f2484_clk;
  logic [0:0] f2484_rst;
  logic [31:0] f2484_rdata;
  sr_buffer_32_1 f2484(.wen(f2484_wen), .wdata(f2484_wdata), .clk(f2484_clk), .rst(f2484_rst), .rdata(f2484_rdata));
  assign f2484_clk = clk;
  assign f2484_rst = rst;
  // Bindings to f2484

  // f2486
  logic [0:0] f2486_wen;
  logic [31:0] f2486_wdata;
  logic [0:0] f2486_clk;
  logic [0:0] f2486_rst;
  logic [31:0] f2486_rdata;
  sr_buffer_32_1 f2486(.wen(f2486_wen), .wdata(f2486_wdata), .clk(f2486_clk), .rst(f2486_rst), .rdata(f2486_rdata));
  assign f2486_clk = clk;
  assign f2486_rst = rst;
  // Bindings to f2486

  // f2488
  logic [0:0] f2488_wen;
  logic [31:0] f2488_wdata;
  logic [0:0] f2488_clk;
  logic [0:0] f2488_rst;
  logic [31:0] f2488_rdata;
  sr_buffer_32_1 f2488(.wen(f2488_wen), .wdata(f2488_wdata), .clk(f2488_clk), .rst(f2488_rst), .rdata(f2488_rdata));
  assign f2488_clk = clk;
  assign f2488_rst = rst;
  // Bindings to f2488

  // f2490
  logic [0:0] f2490_wen;
  logic [31:0] f2490_wdata;
  logic [0:0] f2490_clk;
  logic [0:0] f2490_rst;
  logic [31:0] f2490_rdata;
  sr_buffer_32_1 f2490(.wen(f2490_wen), .wdata(f2490_wdata), .clk(f2490_clk), .rst(f2490_rst), .rdata(f2490_rdata));
  assign f2490_clk = clk;
  assign f2490_rst = rst;
  // Bindings to f2490

  // f2492
  logic [0:0] f2492_wen;
  logic [31:0] f2492_wdata;
  logic [0:0] f2492_clk;
  logic [0:0] f2492_rst;
  logic [31:0] f2492_rdata;
  sr_buffer_32_1 f2492(.wen(f2492_wen), .wdata(f2492_wdata), .clk(f2492_clk), .rst(f2492_rst), .rdata(f2492_rdata));
  assign f2492_clk = clk;
  assign f2492_rst = rst;
  // Bindings to f2492



endmodule


module bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_3790 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f314
  logic [0:0] f314_wen;
  logic [31:0] f314_wdata;
  logic [0:0] f314_clk;
  logic [0:0] f314_rst;
  logic [31:0] f314_rdata;
  sr_buffer_32_1 f314(.wen(f314_wen), .wdata(f314_wdata), .clk(f314_clk), .rst(f314_rst), .rdata(f314_rdata));
  assign f314_clk = clk;
  assign f314_rst = rst;
  // Bindings to f314

  // f316
  logic [0:0] f316_wen;
  logic [31:0] f316_wdata;
  logic [0:0] f316_clk;
  logic [0:0] f316_rst;
  logic [31:0] f316_rdata;
  sr_buffer_32_1 f316(.wen(f316_wen), .wdata(f316_wdata), .clk(f316_clk), .rst(f316_rst), .rdata(f316_rdata));
  assign f316_clk = clk;
  assign f316_rst = rst;
  // Bindings to f316

  // f318
  logic [0:0] f318_wen;
  logic [31:0] f318_wdata;
  logic [0:0] f318_clk;
  logic [0:0] f318_rst;
  logic [31:0] f318_rdata;
  sr_buffer_32_1 f318(.wen(f318_wen), .wdata(f318_wdata), .clk(f318_clk), .rst(f318_rst), .rdata(f318_rdata));
  assign f318_clk = clk;
  assign f318_rst = rst;
  // Bindings to f318

  // f320
  logic [0:0] f320_wen;
  logic [31:0] f320_wdata;
  logic [0:0] f320_clk;
  logic [0:0] f320_rst;
  logic [31:0] f320_rdata;
  sr_buffer_32_1 f320(.wen(f320_wen), .wdata(f320_wdata), .clk(f320_clk), .rst(f320_rst), .rdata(f320_rdata));
  assign f320_clk = clk;
  assign f320_rst = rst;
  // Bindings to f320

  // f322
  logic [0:0] f322_wen;
  logic [31:0] f322_wdata;
  logic [0:0] f322_clk;
  logic [0:0] f322_rst;
  logic [31:0] f322_rdata;
  sr_buffer_32_1 f322(.wen(f322_wen), .wdata(f322_wdata), .clk(f322_clk), .rst(f322_rst), .rdata(f322_rdata));
  assign f322_clk = clk;
  assign f322_rst = rst;
  // Bindings to f322

  // f324
  logic [0:0] f324_wen;
  logic [31:0] f324_wdata;
  logic [0:0] f324_clk;
  logic [0:0] f324_rst;
  logic [31:0] f324_rdata;
  sr_buffer_32_1 f324(.wen(f324_wen), .wdata(f324_wdata), .clk(f324_clk), .rst(f324_rst), .rdata(f324_rdata));
  assign f324_clk = clk;
  assign f324_rst = rst;
  // Bindings to f324

  // f326
  logic [0:0] f326_wen;
  logic [31:0] f326_wdata;
  logic [0:0] f326_clk;
  logic [0:0] f326_rst;
  logic [31:0] f326_rdata;
  sr_buffer_32_1 f326(.wen(f326_wen), .wdata(f326_wdata), .clk(f326_clk), .rst(f326_rst), .rdata(f326_rdata));
  assign f326_clk = clk;
  assign f326_rst = rst;
  // Bindings to f326

  // f328
  logic [0:0] f328_wen;
  logic [31:0] f328_wdata;
  logic [0:0] f328_clk;
  logic [0:0] f328_rst;
  logic [31:0] f328_rdata;
  sr_buffer_32_1 f328(.wen(f328_wen), .wdata(f328_wdata), .clk(f328_clk), .rst(f328_rst), .rdata(f328_rdata));
  assign f328_clk = clk;
  assign f328_rst = rst;
  // Bindings to f328

  // f330
  logic [0:0] f330_wen;
  logic [31:0] f330_wdata;
  logic [0:0] f330_clk;
  logic [0:0] f330_rst;
  logic [31:0] f330_rdata;
  sr_buffer_32_1 f330(.wen(f330_wen), .wdata(f330_wdata), .clk(f330_clk), .rst(f330_rst), .rdata(f330_rdata));
  assign f330_clk = clk;
  assign f330_rst = rst;
  // Bindings to f330

  // f332
  logic [0:0] f332_wen;
  logic [31:0] f332_wdata;
  logic [0:0] f332_clk;
  logic [0:0] f332_rst;
  logic [31:0] f332_rdata;
  sr_buffer_32_1 f332(.wen(f332_wen), .wdata(f332_wdata), .clk(f332_clk), .rst(f332_rst), .rdata(f332_rdata));
  assign f332_clk = clk;
  assign f332_rst = rst;
  // Bindings to f332

  // f334
  logic [0:0] f334_wen;
  logic [31:0] f334_wdata;
  logic [0:0] f334_clk;
  logic [0:0] f334_rst;
  logic [31:0] f334_rdata;
  sr_buffer_32_1 f334(.wen(f334_wen), .wdata(f334_wdata), .clk(f334_clk), .rst(f334_rst), .rdata(f334_rdata));
  assign f334_clk = clk;
  assign f334_rst = rst;
  // Bindings to f334

  // f336
  logic [0:0] f336_wen;
  logic [31:0] f336_wdata;
  logic [0:0] f336_clk;
  logic [0:0] f336_rst;
  logic [31:0] f336_rdata;
  sr_buffer_32_1 f336(.wen(f336_wen), .wdata(f336_wdata), .clk(f336_clk), .rst(f336_rst), .rdata(f336_rdata));
  assign f336_clk = clk;
  assign f336_rst = rst;
  // Bindings to f336

  // f338
  logic [0:0] f338_wen;
  logic [31:0] f338_wdata;
  logic [0:0] f338_clk;
  logic [0:0] f338_rst;
  logic [31:0] f338_rdata;
  sr_buffer_32_1 f338(.wen(f338_wen), .wdata(f338_wdata), .clk(f338_clk), .rst(f338_rst), .rdata(f338_rdata));
  assign f338_clk = clk;
  assign f338_rst = rst;
  // Bindings to f338

  // f340
  logic [0:0] f340_wen;
  logic [31:0] f340_wdata;
  logic [0:0] f340_clk;
  logic [0:0] f340_rst;
  logic [31:0] f340_rdata;
  sr_buffer_32_1 f340(.wen(f340_wen), .wdata(f340_wdata), .clk(f340_clk), .rst(f340_rst), .rdata(f340_rdata));
  assign f340_clk = clk;
  assign f340_rst = rst;
  // Bindings to f340

  // f342
  logic [0:0] f342_wen;
  logic [31:0] f342_wdata;
  logic [0:0] f342_clk;
  logic [0:0] f342_rst;
  logic [31:0] f342_rdata;
  sr_buffer_32_1 f342(.wen(f342_wen), .wdata(f342_wdata), .clk(f342_clk), .rst(f342_rst), .rdata(f342_rdata));
  assign f342_clk = clk;
  assign f342_rst = rst;
  // Bindings to f342

  // f344
  logic [0:0] f344_wen;
  logic [31:0] f344_wdata;
  logic [0:0] f344_clk;
  logic [0:0] f344_rst;
  logic [31:0] f344_rdata;
  sr_buffer_32_1 f344(.wen(f344_wen), .wdata(f344_wdata), .clk(f344_clk), .rst(f344_rst), .rdata(f344_rdata));
  assign f344_clk = clk;
  assign f344_rst = rst;
  // Bindings to f344

  // f346
  logic [0:0] f346_wen;
  logic [31:0] f346_wdata;
  logic [0:0] f346_clk;
  logic [0:0] f346_rst;
  logic [31:0] f346_rdata;
  sr_buffer_32_1 f346(.wen(f346_wen), .wdata(f346_wdata), .clk(f346_clk), .rst(f346_rst), .rdata(f346_rdata));
  assign f346_clk = clk;
  assign f346_rst = rst;
  // Bindings to f346

  // f348
  logic [0:0] f348_wen;
  logic [31:0] f348_wdata;
  logic [0:0] f348_clk;
  logic [0:0] f348_rst;
  logic [31:0] f348_rdata;
  sr_buffer_32_1 f348(.wen(f348_wen), .wdata(f348_wdata), .clk(f348_clk), .rst(f348_rst), .rdata(f348_rdata));
  assign f348_clk = clk;
  assign f348_rst = rst;
  // Bindings to f348

  // f350
  logic [0:0] f350_wen;
  logic [31:0] f350_wdata;
  logic [0:0] f350_clk;
  logic [0:0] f350_rst;
  logic [31:0] f350_rdata;
  sr_buffer_32_1 f350(.wen(f350_wen), .wdata(f350_wdata), .clk(f350_clk), .rst(f350_rst), .rdata(f350_rdata));
  assign f350_clk = clk;
  assign f350_rst = rst;
  // Bindings to f350

  // f352
  logic [0:0] f352_wen;
  logic [31:0] f352_wdata;
  logic [0:0] f352_clk;
  logic [0:0] f352_rst;
  logic [31:0] f352_rdata;
  sr_buffer_32_1 f352(.wen(f352_wen), .wdata(f352_wdata), .clk(f352_clk), .rst(f352_rst), .rdata(f352_rdata));
  assign f352_clk = clk;
  assign f352_rst = rst;
  // Bindings to f352

  // f354
  logic [0:0] f354_wen;
  logic [31:0] f354_wdata;
  logic [0:0] f354_clk;
  logic [0:0] f354_rst;
  logic [31:0] f354_rdata;
  sr_buffer_32_1 f354(.wen(f354_wen), .wdata(f354_wdata), .clk(f354_clk), .rst(f354_rst), .rdata(f354_rdata));
  assign f354_clk = clk;
  assign f354_rst = rst;
  // Bindings to f354

  // f356
  logic [0:0] f356_wen;
  logic [31:0] f356_wdata;
  logic [0:0] f356_clk;
  logic [0:0] f356_rst;
  logic [31:0] f356_rdata;
  sr_buffer_32_1 f356(.wen(f356_wen), .wdata(f356_wdata), .clk(f356_clk), .rst(f356_rst), .rdata(f356_rdata));
  assign f356_clk = clk;
  assign f356_rst = rst;
  // Bindings to f356

  // f358
  logic [0:0] f358_wen;
  logic [31:0] f358_wdata;
  logic [0:0] f358_clk;
  logic [0:0] f358_rst;
  logic [31:0] f358_rdata;
  sr_buffer_32_1 f358(.wen(f358_wen), .wdata(f358_wdata), .clk(f358_clk), .rst(f358_rst), .rdata(f358_rdata));
  assign f358_clk = clk;
  assign f358_rst = rst;
  // Bindings to f358

  // f360
  logic [0:0] f360_wen;
  logic [31:0] f360_wdata;
  logic [0:0] f360_clk;
  logic [0:0] f360_rst;
  logic [31:0] f360_rdata;
  sr_buffer_32_1 f360(.wen(f360_wen), .wdata(f360_wdata), .clk(f360_clk), .rst(f360_rst), .rdata(f360_rdata));
  assign f360_clk = clk;
  assign f360_rst = rst;
  // Bindings to f360

  // f362
  logic [0:0] f362_wen;
  logic [31:0] f362_wdata;
  logic [0:0] f362_clk;
  logic [0:0] f362_rst;
  logic [31:0] f362_rdata;
  sr_buffer_32_1 f362(.wen(f362_wen), .wdata(f362_wdata), .clk(f362_clk), .rst(f362_rst), .rdata(f362_rdata));
  assign f362_clk = clk;
  assign f362_rst = rst;
  // Bindings to f362

  // f364
  logic [0:0] f364_wen;
  logic [31:0] f364_wdata;
  logic [0:0] f364_clk;
  logic [0:0] f364_rst;
  logic [31:0] f364_rdata;
  sr_buffer_32_1 f364(.wen(f364_wen), .wdata(f364_wdata), .clk(f364_clk), .rst(f364_rst), .rdata(f364_rdata));
  assign f364_clk = clk;
  assign f364_rst = rst;
  // Bindings to f364

  // f366
  logic [0:0] f366_wen;
  logic [31:0] f366_wdata;
  logic [0:0] f366_clk;
  logic [0:0] f366_rst;
  logic [31:0] f366_rdata;
  sr_buffer_32_1 f366(.wen(f366_wen), .wdata(f366_wdata), .clk(f366_clk), .rst(f366_rst), .rdata(f366_rdata));
  assign f366_clk = clk;
  assign f366_rst = rst;
  // Bindings to f366

  // f368
  logic [0:0] f368_wen;
  logic [31:0] f368_wdata;
  logic [0:0] f368_clk;
  logic [0:0] f368_rst;
  logic [31:0] f368_rdata;
  sr_buffer_32_1 f368(.wen(f368_wen), .wdata(f368_wdata), .clk(f368_clk), .rst(f368_rst), .rdata(f368_rdata));
  assign f368_clk = clk;
  assign f368_rst = rst;
  // Bindings to f368

  // f370
  logic [0:0] f370_wen;
  logic [31:0] f370_wdata;
  logic [0:0] f370_clk;
  logic [0:0] f370_rst;
  logic [31:0] f370_rdata;
  sr_buffer_32_1 f370(.wen(f370_wen), .wdata(f370_wdata), .clk(f370_clk), .rst(f370_rst), .rdata(f370_rdata));
  assign f370_clk = clk;
  assign f370_rst = rst;
  // Bindings to f370

  // f372
  logic [0:0] f372_wen;
  logic [31:0] f372_wdata;
  logic [0:0] f372_clk;
  logic [0:0] f372_rst;
  logic [31:0] f372_rdata;
  sr_buffer_32_1 f372(.wen(f372_wen), .wdata(f372_wdata), .clk(f372_clk), .rst(f372_rst), .rdata(f372_rdata));
  assign f372_clk = clk;
  assign f372_rst = rst;
  // Bindings to f372

  // f374
  logic [0:0] f374_wen;
  logic [31:0] f374_wdata;
  logic [0:0] f374_clk;
  logic [0:0] f374_rst;
  logic [31:0] f374_rdata;
  sr_buffer_32_1 f374(.wen(f374_wen), .wdata(f374_wdata), .clk(f374_clk), .rst(f374_rst), .rdata(f374_rdata));
  assign f374_clk = clk;
  assign f374_rst = rst;
  // Bindings to f374

  // f376
  logic [0:0] f376_wen;
  logic [31:0] f376_wdata;
  logic [0:0] f376_clk;
  logic [0:0] f376_rst;
  logic [31:0] f376_rdata;
  sr_buffer_32_1 f376(.wen(f376_wen), .wdata(f376_wdata), .clk(f376_clk), .rst(f376_rst), .rdata(f376_rdata));
  assign f376_clk = clk;
  assign f376_rst = rst;
  // Bindings to f376

  // f378
  logic [0:0] f378_wen;
  logic [31:0] f378_wdata;
  logic [0:0] f378_clk;
  logic [0:0] f378_rst;
  logic [31:0] f378_rdata;
  sr_buffer_32_1 f378(.wen(f378_wen), .wdata(f378_wdata), .clk(f378_clk), .rst(f378_rst), .rdata(f378_rdata));
  assign f378_clk = clk;
  assign f378_rst = rst;
  // Bindings to f378

  // f380
  logic [0:0] f380_wen;
  logic [31:0] f380_wdata;
  logic [0:0] f380_clk;
  logic [0:0] f380_rst;
  logic [31:0] f380_rdata;
  sr_buffer_32_1 f380(.wen(f380_wen), .wdata(f380_wdata), .clk(f380_clk), .rst(f380_rst), .rdata(f380_rdata));
  assign f380_clk = clk;
  assign f380_rst = rst;
  // Bindings to f380

  // f382
  logic [0:0] f382_wen;
  logic [31:0] f382_wdata;
  logic [0:0] f382_clk;
  logic [0:0] f382_rst;
  logic [31:0] f382_rdata;
  sr_buffer_32_1 f382(.wen(f382_wen), .wdata(f382_wdata), .clk(f382_clk), .rst(f382_rst), .rdata(f382_rdata));
  assign f382_clk = clk;
  assign f382_rst = rst;
  // Bindings to f382

  // f384
  logic [0:0] f384_wen;
  logic [31:0] f384_wdata;
  logic [0:0] f384_clk;
  logic [0:0] f384_rst;
  logic [31:0] f384_rdata;
  sr_buffer_32_1 f384(.wen(f384_wen), .wdata(f384_wdata), .clk(f384_clk), .rst(f384_rst), .rdata(f384_rdata));
  assign f384_clk = clk;
  assign f384_rst = rst;
  // Bindings to f384

  // f386
  logic [0:0] f386_wen;
  logic [31:0] f386_wdata;
  logic [0:0] f386_clk;
  logic [0:0] f386_rst;
  logic [31:0] f386_rdata;
  sr_buffer_32_1 f386(.wen(f386_wen), .wdata(f386_wdata), .clk(f386_clk), .rst(f386_rst), .rdata(f386_rdata));
  assign f386_clk = clk;
  assign f386_rst = rst;
  // Bindings to f386

  // f388
  logic [0:0] f388_wen;
  logic [31:0] f388_wdata;
  logic [0:0] f388_clk;
  logic [0:0] f388_rst;
  logic [31:0] f388_rdata;
  sr_buffer_32_1 f388(.wen(f388_wen), .wdata(f388_wdata), .clk(f388_clk), .rst(f388_rst), .rdata(f388_rdata));
  assign f388_clk = clk;
  assign f388_rst = rst;
  // Bindings to f388

  // f390
  logic [0:0] f390_wen;
  logic [31:0] f390_wdata;
  logic [0:0] f390_clk;
  logic [0:0] f390_rst;
  logic [31:0] f390_rdata;
  sr_buffer_32_1 f390(.wen(f390_wen), .wdata(f390_wdata), .clk(f390_clk), .rst(f390_rst), .rdata(f390_rdata));
  assign f390_clk = clk;
  assign f390_rst = rst;
  // Bindings to f390

  // f392
  logic [0:0] f392_wen;
  logic [31:0] f392_wdata;
  logic [0:0] f392_clk;
  logic [0:0] f392_rst;
  logic [31:0] f392_rdata;
  sr_buffer_32_1 f392(.wen(f392_wen), .wdata(f392_wdata), .clk(f392_clk), .rst(f392_rst), .rdata(f392_rdata));
  assign f392_clk = clk;
  assign f392_rst = rst;
  // Bindings to f392

  // f394
  logic [0:0] f394_wen;
  logic [31:0] f394_wdata;
  logic [0:0] f394_clk;
  logic [0:0] f394_rst;
  logic [31:0] f394_rdata;
  sr_buffer_32_1 f394(.wen(f394_wen), .wdata(f394_wdata), .clk(f394_clk), .rst(f394_rst), .rdata(f394_rdata));
  assign f394_clk = clk;
  assign f394_rst = rst;
  // Bindings to f394

  // f396
  logic [0:0] f396_wen;
  logic [31:0] f396_wdata;
  logic [0:0] f396_clk;
  logic [0:0] f396_rst;
  logic [31:0] f396_rdata;
  sr_buffer_32_1 f396(.wen(f396_wen), .wdata(f396_wdata), .clk(f396_clk), .rst(f396_rst), .rdata(f396_rdata));
  assign f396_clk = clk;
  assign f396_rst = rst;
  // Bindings to f396

  // f398
  logic [0:0] f398_wen;
  logic [31:0] f398_wdata;
  logic [0:0] f398_clk;
  logic [0:0] f398_rst;
  logic [31:0] f398_rdata;
  sr_buffer_32_1 f398(.wen(f398_wen), .wdata(f398_wdata), .clk(f398_clk), .rst(f398_rst), .rdata(f398_rdata));
  assign f398_clk = clk;
  assign f398_rst = rst;
  // Bindings to f398

  // f400
  logic [0:0] f400_wen;
  logic [31:0] f400_wdata;
  logic [0:0] f400_clk;
  logic [0:0] f400_rst;
  logic [31:0] f400_rdata;
  sr_buffer_32_1 f400(.wen(f400_wen), .wdata(f400_wdata), .clk(f400_clk), .rst(f400_rst), .rdata(f400_rdata));
  assign f400_clk = clk;
  assign f400_rst = rst;
  // Bindings to f400

  // f402
  logic [0:0] f402_wen;
  logic [31:0] f402_wdata;
  logic [0:0] f402_clk;
  logic [0:0] f402_rst;
  logic [31:0] f402_rdata;
  sr_buffer_32_1 f402(.wen(f402_wen), .wdata(f402_wdata), .clk(f402_clk), .rst(f402_rst), .rdata(f402_rdata));
  assign f402_clk = clk;
  assign f402_rst = rst;
  // Bindings to f402

  // f404
  logic [0:0] f404_wen;
  logic [31:0] f404_wdata;
  logic [0:0] f404_clk;
  logic [0:0] f404_rst;
  logic [31:0] f404_rdata;
  sr_buffer_32_1 f404(.wen(f404_wen), .wdata(f404_wdata), .clk(f404_clk), .rst(f404_rst), .rdata(f404_rdata));
  assign f404_clk = clk;
  assign f404_rst = rst;
  // Bindings to f404

  // f406
  logic [0:0] f406_wen;
  logic [31:0] f406_wdata;
  logic [0:0] f406_clk;
  logic [0:0] f406_rst;
  logic [31:0] f406_rdata;
  sr_buffer_32_1 f406(.wen(f406_wen), .wdata(f406_wdata), .clk(f406_clk), .rst(f406_rst), .rdata(f406_rdata));
  assign f406_clk = clk;
  assign f406_rst = rst;
  // Bindings to f406

  // f408
  logic [0:0] f408_wen;
  logic [31:0] f408_wdata;
  logic [0:0] f408_clk;
  logic [0:0] f408_rst;
  logic [31:0] f408_rdata;
  sr_buffer_32_1 f408(.wen(f408_wen), .wdata(f408_wdata), .clk(f408_clk), .rst(f408_rst), .rdata(f408_rdata));
  assign f408_clk = clk;
  assign f408_rst = rst;
  // Bindings to f408

  // f410
  logic [0:0] f410_wen;
  logic [31:0] f410_wdata;
  logic [0:0] f410_clk;
  logic [0:0] f410_rst;
  logic [31:0] f410_rdata;
  sr_buffer_32_1 f410(.wen(f410_wen), .wdata(f410_wdata), .clk(f410_clk), .rst(f410_rst), .rdata(f410_rdata));
  assign f410_clk = clk;
  assign f410_rst = rst;
  // Bindings to f410

  // f412
  logic [0:0] f412_wen;
  logic [31:0] f412_wdata;
  logic [0:0] f412_clk;
  logic [0:0] f412_rst;
  logic [31:0] f412_rdata;
  sr_buffer_32_1 f412(.wen(f412_wen), .wdata(f412_wdata), .clk(f412_clk), .rst(f412_rst), .rdata(f412_rdata));
  assign f412_clk = clk;
  assign f412_rst = rst;
  // Bindings to f412

  // f414
  logic [0:0] f414_wen;
  logic [31:0] f414_wdata;
  logic [0:0] f414_clk;
  logic [0:0] f414_rst;
  logic [31:0] f414_rdata;
  sr_buffer_32_1 f414(.wen(f414_wen), .wdata(f414_wdata), .clk(f414_clk), .rst(f414_rst), .rdata(f414_rdata));
  assign f414_clk = clk;
  assign f414_rst = rst;
  // Bindings to f414

  // f416
  logic [0:0] f416_wen;
  logic [31:0] f416_wdata;
  logic [0:0] f416_clk;
  logic [0:0] f416_rst;
  logic [31:0] f416_rdata;
  sr_buffer_32_1 f416(.wen(f416_wen), .wdata(f416_wdata), .clk(f416_clk), .rst(f416_rst), .rdata(f416_rdata));
  assign f416_clk = clk;
  assign f416_rst = rst;
  // Bindings to f416

  // f418
  logic [0:0] f418_wen;
  logic [31:0] f418_wdata;
  logic [0:0] f418_clk;
  logic [0:0] f418_rst;
  logic [31:0] f418_rdata;
  sr_buffer_32_1 f418(.wen(f418_wen), .wdata(f418_wdata), .clk(f418_clk), .rst(f418_rst), .rdata(f418_rdata));
  assign f418_clk = clk;
  assign f418_rst = rst;
  // Bindings to f418

  // f420
  logic [0:0] f420_wen;
  logic [31:0] f420_wdata;
  logic [0:0] f420_clk;
  logic [0:0] f420_rst;
  logic [31:0] f420_rdata;
  sr_buffer_32_1 f420(.wen(f420_wen), .wdata(f420_wdata), .clk(f420_clk), .rst(f420_rst), .rdata(f420_rdata));
  assign f420_clk = clk;
  assign f420_rst = rst;
  // Bindings to f420

  // f422
  logic [0:0] f422_wen;
  logic [31:0] f422_wdata;
  logic [0:0] f422_clk;
  logic [0:0] f422_rst;
  logic [31:0] f422_rdata;
  sr_buffer_32_1 f422(.wen(f422_wen), .wdata(f422_wdata), .clk(f422_clk), .rst(f422_rst), .rdata(f422_rdata));
  assign f422_clk = clk;
  assign f422_rst = rst;
  // Bindings to f422

  // f424
  logic [0:0] f424_wen;
  logic [31:0] f424_wdata;
  logic [0:0] f424_clk;
  logic [0:0] f424_rst;
  logic [31:0] f424_rdata;
  sr_buffer_32_1 f424(.wen(f424_wen), .wdata(f424_wdata), .clk(f424_clk), .rst(f424_rst), .rdata(f424_rdata));
  assign f424_clk = clk;
  assign f424_rst = rst;
  // Bindings to f424

  // f426
  logic [0:0] f426_wen;
  logic [31:0] f426_wdata;
  logic [0:0] f426_clk;
  logic [0:0] f426_rst;
  logic [31:0] f426_rdata;
  sr_buffer_32_1 f426(.wen(f426_wen), .wdata(f426_wdata), .clk(f426_clk), .rst(f426_rst), .rdata(f426_rdata));
  assign f426_clk = clk;
  assign f426_rst = rst;
  // Bindings to f426

  // f428
  logic [0:0] f428_wen;
  logic [31:0] f428_wdata;
  logic [0:0] f428_clk;
  logic [0:0] f428_rst;
  logic [31:0] f428_rdata;
  sr_buffer_32_1 f428(.wen(f428_wen), .wdata(f428_wdata), .clk(f428_clk), .rst(f428_rst), .rdata(f428_rdata));
  assign f428_clk = clk;
  assign f428_rst = rst;
  // Bindings to f428

  // f430
  logic [0:0] f430_wen;
  logic [31:0] f430_wdata;
  logic [0:0] f430_clk;
  logic [0:0] f430_rst;
  logic [31:0] f430_rdata;
  sr_buffer_32_1 f430(.wen(f430_wen), .wdata(f430_wdata), .clk(f430_clk), .rst(f430_rst), .rdata(f430_rdata));
  assign f430_clk = clk;
  assign f430_rst = rst;
  // Bindings to f430

  // f432
  logic [0:0] f432_wen;
  logic [31:0] f432_wdata;
  logic [0:0] f432_clk;
  logic [0:0] f432_rst;
  logic [31:0] f432_rdata;
  sr_buffer_32_1 f432(.wen(f432_wen), .wdata(f432_wdata), .clk(f432_clk), .rst(f432_rst), .rdata(f432_rdata));
  assign f432_clk = clk;
  assign f432_rst = rst;
  // Bindings to f432

  // f434
  logic [0:0] f434_wen;
  logic [31:0] f434_wdata;
  logic [0:0] f434_clk;
  logic [0:0] f434_rst;
  logic [31:0] f434_rdata;
  sr_buffer_32_1 f434(.wen(f434_wen), .wdata(f434_wdata), .clk(f434_clk), .rst(f434_rst), .rdata(f434_rdata));
  assign f434_clk = clk;
  assign f434_rst = rst;
  // Bindings to f434

  // f436
  logic [0:0] f436_wen;
  logic [31:0] f436_wdata;
  logic [0:0] f436_clk;
  logic [0:0] f436_rst;
  logic [31:0] f436_rdata;
  sr_buffer_32_1 f436(.wen(f436_wen), .wdata(f436_wdata), .clk(f436_clk), .rst(f436_rst), .rdata(f436_rdata));
  assign f436_clk = clk;
  assign f436_rst = rst;
  // Bindings to f436

  // f438
  logic [0:0] f438_wen;
  logic [31:0] f438_wdata;
  logic [0:0] f438_clk;
  logic [0:0] f438_rst;
  logic [31:0] f438_rdata;
  sr_buffer_32_1 f438(.wen(f438_wen), .wdata(f438_wdata), .clk(f438_clk), .rst(f438_rst), .rdata(f438_rdata));
  assign f438_clk = clk;
  assign f438_rst = rst;
  // Bindings to f438

  // f440
  logic [0:0] f440_wen;
  logic [31:0] f440_wdata;
  logic [0:0] f440_clk;
  logic [0:0] f440_rst;
  logic [31:0] f440_rdata;
  sr_buffer_32_1 f440(.wen(f440_wen), .wdata(f440_wdata), .clk(f440_clk), .rst(f440_rst), .rdata(f440_rdata));
  assign f440_clk = clk;
  assign f440_rst = rst;
  // Bindings to f440

  // f442
  logic [0:0] f442_wen;
  logic [31:0] f442_wdata;
  logic [0:0] f442_clk;
  logic [0:0] f442_rst;
  logic [31:0] f442_rdata;
  sr_buffer_32_1 f442(.wen(f442_wen), .wdata(f442_wdata), .clk(f442_clk), .rst(f442_rst), .rdata(f442_rdata));
  assign f442_clk = clk;
  assign f442_rst = rst;
  // Bindings to f442

  // f444
  logic [0:0] f444_wen;
  logic [31:0] f444_wdata;
  logic [0:0] f444_clk;
  logic [0:0] f444_rst;
  logic [31:0] f444_rdata;
  sr_buffer_32_1 f444(.wen(f444_wen), .wdata(f444_wdata), .clk(f444_clk), .rst(f444_rst), .rdata(f444_rdata));
  assign f444_clk = clk;
  assign f444_rst = rst;
  // Bindings to f444

  // f446
  logic [0:0] f446_wen;
  logic [31:0] f446_wdata;
  logic [0:0] f446_clk;
  logic [0:0] f446_rst;
  logic [31:0] f446_rdata;
  sr_buffer_32_1 f446(.wen(f446_wen), .wdata(f446_wdata), .clk(f446_clk), .rst(f446_rst), .rdata(f446_rdata));
  assign f446_clk = clk;
  assign f446_rst = rst;
  // Bindings to f446

  // f448
  logic [0:0] f448_wen;
  logic [31:0] f448_wdata;
  logic [0:0] f448_clk;
  logic [0:0] f448_rst;
  logic [31:0] f448_rdata;
  sr_buffer_32_1 f448(.wen(f448_wen), .wdata(f448_wdata), .clk(f448_clk), .rst(f448_rst), .rdata(f448_rdata));
  assign f448_clk = clk;
  assign f448_rst = rst;
  // Bindings to f448

  // f450
  logic [0:0] f450_wen;
  logic [31:0] f450_wdata;
  logic [0:0] f450_clk;
  logic [0:0] f450_rst;
  logic [31:0] f450_rdata;
  sr_buffer_32_1 f450(.wen(f450_wen), .wdata(f450_wdata), .clk(f450_clk), .rst(f450_rst), .rdata(f450_rdata));
  assign f450_clk = clk;
  assign f450_rst = rst;
  // Bindings to f450

  // f452
  logic [0:0] f452_wen;
  logic [31:0] f452_wdata;
  logic [0:0] f452_clk;
  logic [0:0] f452_rst;
  logic [31:0] f452_rdata;
  sr_buffer_32_1 f452(.wen(f452_wen), .wdata(f452_wdata), .clk(f452_clk), .rst(f452_rst), .rdata(f452_rdata));
  assign f452_clk = clk;
  assign f452_rst = rst;
  // Bindings to f452

  // f454
  logic [0:0] f454_wen;
  logic [31:0] f454_wdata;
  logic [0:0] f454_clk;
  logic [0:0] f454_rst;
  logic [31:0] f454_rdata;
  sr_buffer_32_1 f454(.wen(f454_wen), .wdata(f454_wdata), .clk(f454_clk), .rst(f454_rst), .rdata(f454_rdata));
  assign f454_clk = clk;
  assign f454_rst = rst;
  // Bindings to f454

  // f456
  logic [0:0] f456_wen;
  logic [31:0] f456_wdata;
  logic [0:0] f456_clk;
  logic [0:0] f456_rst;
  logic [31:0] f456_rdata;
  sr_buffer_32_1 f456(.wen(f456_wen), .wdata(f456_wdata), .clk(f456_clk), .rst(f456_rst), .rdata(f456_rdata));
  assign f456_clk = clk;
  assign f456_rst = rst;
  // Bindings to f456

  // f458
  logic [0:0] f458_wen;
  logic [31:0] f458_wdata;
  logic [0:0] f458_clk;
  logic [0:0] f458_rst;
  logic [31:0] f458_rdata;
  sr_buffer_32_1 f458(.wen(f458_wen), .wdata(f458_wdata), .clk(f458_clk), .rst(f458_rst), .rdata(f458_rdata));
  assign f458_clk = clk;
  assign f458_rst = rst;
  // Bindings to f458

  // f460
  logic [0:0] f460_wen;
  logic [31:0] f460_wdata;
  logic [0:0] f460_clk;
  logic [0:0] f460_rst;
  logic [31:0] f460_rdata;
  sr_buffer_32_1 f460(.wen(f460_wen), .wdata(f460_wdata), .clk(f460_clk), .rst(f460_rst), .rdata(f460_rdata));
  assign f460_clk = clk;
  assign f460_rst = rst;
  // Bindings to f460

  // f462
  logic [0:0] f462_wen;
  logic [31:0] f462_wdata;
  logic [0:0] f462_clk;
  logic [0:0] f462_rst;
  logic [31:0] f462_rdata;
  sr_buffer_32_1 f462(.wen(f462_wen), .wdata(f462_wdata), .clk(f462_clk), .rst(f462_rst), .rdata(f462_rdata));
  assign f462_clk = clk;
  assign f462_rst = rst;
  // Bindings to f462

  // f464
  logic [0:0] f464_wen;
  logic [31:0] f464_wdata;
  logic [0:0] f464_clk;
  logic [0:0] f464_rst;
  logic [31:0] f464_rdata;
  sr_buffer_32_1 f464(.wen(f464_wen), .wdata(f464_wdata), .clk(f464_clk), .rst(f464_rst), .rdata(f464_rdata));
  assign f464_clk = clk;
  assign f464_rst = rst;
  // Bindings to f464

  // f466
  logic [0:0] f466_wen;
  logic [31:0] f466_wdata;
  logic [0:0] f466_clk;
  logic [0:0] f466_rst;
  logic [31:0] f466_rdata;
  sr_buffer_32_1 f466(.wen(f466_wen), .wdata(f466_wdata), .clk(f466_clk), .rst(f466_rst), .rdata(f466_rdata));
  assign f466_clk = clk;
  assign f466_rst = rst;
  // Bindings to f466

  // f468
  logic [0:0] f468_wen;
  logic [31:0] f468_wdata;
  logic [0:0] f468_clk;
  logic [0:0] f468_rst;
  logic [31:0] f468_rdata;
  sr_buffer_32_1 f468(.wen(f468_wen), .wdata(f468_wdata), .clk(f468_clk), .rst(f468_rst), .rdata(f468_rdata));
  assign f468_clk = clk;
  assign f468_rst = rst;
  // Bindings to f468

  // f470
  logic [0:0] f470_wen;
  logic [31:0] f470_wdata;
  logic [0:0] f470_clk;
  logic [0:0] f470_rst;
  logic [31:0] f470_rdata;
  sr_buffer_32_1 f470(.wen(f470_wen), .wdata(f470_wdata), .clk(f470_clk), .rst(f470_rst), .rdata(f470_rdata));
  assign f470_clk = clk;
  assign f470_rst = rst;
  // Bindings to f470

  // f472
  logic [0:0] f472_wen;
  logic [31:0] f472_wdata;
  logic [0:0] f472_clk;
  logic [0:0] f472_rst;
  logic [31:0] f472_rdata;
  sr_buffer_32_1 f472(.wen(f472_wen), .wdata(f472_wdata), .clk(f472_clk), .rst(f472_rst), .rdata(f472_rdata));
  assign f472_clk = clk;
  assign f472_rst = rst;
  // Bindings to f472

  // f474
  logic [0:0] f474_wen;
  logic [31:0] f474_wdata;
  logic [0:0] f474_clk;
  logic [0:0] f474_rst;
  logic [31:0] f474_rdata;
  sr_buffer_32_1 f474(.wen(f474_wen), .wdata(f474_wdata), .clk(f474_clk), .rst(f474_rst), .rdata(f474_rdata));
  assign f474_clk = clk;
  assign f474_rst = rst;
  // Bindings to f474

  // f476
  logic [0:0] f476_wen;
  logic [31:0] f476_wdata;
  logic [0:0] f476_clk;
  logic [0:0] f476_rst;
  logic [31:0] f476_rdata;
  sr_buffer_32_1 f476(.wen(f476_wen), .wdata(f476_wdata), .clk(f476_clk), .rst(f476_rst), .rdata(f476_rdata));
  assign f476_clk = clk;
  assign f476_rst = rst;
  // Bindings to f476

  // f478
  logic [0:0] f478_wen;
  logic [31:0] f478_wdata;
  logic [0:0] f478_clk;
  logic [0:0] f478_rst;
  logic [31:0] f478_rdata;
  sr_buffer_32_1 f478(.wen(f478_wen), .wdata(f478_wdata), .clk(f478_clk), .rst(f478_rst), .rdata(f478_rdata));
  assign f478_clk = clk;
  assign f478_rst = rst;
  // Bindings to f478

  // f480
  logic [0:0] f480_wen;
  logic [31:0] f480_wdata;
  logic [0:0] f480_clk;
  logic [0:0] f480_rst;
  logic [31:0] f480_rdata;
  sr_buffer_32_1 f480(.wen(f480_wen), .wdata(f480_wdata), .clk(f480_clk), .rst(f480_rst), .rdata(f480_rdata));
  assign f480_clk = clk;
  assign f480_rst = rst;
  // Bindings to f480

  // f482
  logic [0:0] f482_wen;
  logic [31:0] f482_wdata;
  logic [0:0] f482_clk;
  logic [0:0] f482_rst;
  logic [31:0] f482_rdata;
  sr_buffer_32_1 f482(.wen(f482_wen), .wdata(f482_wdata), .clk(f482_clk), .rst(f482_rst), .rdata(f482_rdata));
  assign f482_clk = clk;
  assign f482_rst = rst;
  // Bindings to f482

  // f484
  logic [0:0] f484_wen;
  logic [31:0] f484_wdata;
  logic [0:0] f484_clk;
  logic [0:0] f484_rst;
  logic [31:0] f484_rdata;
  sr_buffer_32_1 f484(.wen(f484_wen), .wdata(f484_wdata), .clk(f484_clk), .rst(f484_rst), .rdata(f484_rdata));
  assign f484_clk = clk;
  assign f484_rst = rst;
  // Bindings to f484

  // f486
  logic [0:0] f486_wen;
  logic [31:0] f486_wdata;
  logic [0:0] f486_clk;
  logic [0:0] f486_rst;
  logic [31:0] f486_rdata;
  sr_buffer_32_1 f486(.wen(f486_wen), .wdata(f486_wdata), .clk(f486_clk), .rst(f486_rst), .rdata(f486_rdata));
  assign f486_clk = clk;
  assign f486_rst = rst;
  // Bindings to f486

  // f488
  logic [0:0] f488_wen;
  logic [31:0] f488_wdata;
  logic [0:0] f488_clk;
  logic [0:0] f488_rst;
  logic [31:0] f488_rdata;
  sr_buffer_32_1 f488(.wen(f488_wen), .wdata(f488_wdata), .clk(f488_clk), .rst(f488_rst), .rdata(f488_rdata));
  assign f488_clk = clk;
  assign f488_rst = rst;
  // Bindings to f488

  // f490
  logic [0:0] f490_wen;
  logic [31:0] f490_wdata;
  logic [0:0] f490_clk;
  logic [0:0] f490_rst;
  logic [31:0] f490_rdata;
  sr_buffer_32_1 f490(.wen(f490_wen), .wdata(f490_wdata), .clk(f490_clk), .rst(f490_rst), .rdata(f490_rdata));
  assign f490_clk = clk;
  assign f490_rst = rst;
  // Bindings to f490

  // f492
  logic [0:0] f492_wen;
  logic [31:0] f492_wdata;
  logic [0:0] f492_clk;
  logic [0:0] f492_rst;
  logic [31:0] f492_rdata;
  sr_buffer_32_1 f492(.wen(f492_wen), .wdata(f492_wdata), .clk(f492_clk), .rst(f492_rst), .rdata(f492_rdata));
  assign f492_clk = clk;
  assign f492_rst = rst;
  // Bindings to f492

  // f494
  logic [0:0] f494_wen;
  logic [31:0] f494_wdata;
  logic [0:0] f494_clk;
  logic [0:0] f494_rst;
  logic [31:0] f494_rdata;
  sr_buffer_32_1 f494(.wen(f494_wen), .wdata(f494_wdata), .clk(f494_clk), .rst(f494_rst), .rdata(f494_rdata));
  assign f494_clk = clk;
  assign f494_rst = rst;
  // Bindings to f494

  // f496
  logic [0:0] f496_wen;
  logic [31:0] f496_wdata;
  logic [0:0] f496_clk;
  logic [0:0] f496_rst;
  logic [31:0] f496_rdata;
  sr_buffer_32_1 f496(.wen(f496_wen), .wdata(f496_wdata), .clk(f496_clk), .rst(f496_rst), .rdata(f496_rdata));
  assign f496_clk = clk;
  assign f496_rst = rst;
  // Bindings to f496

  // f498
  logic [0:0] f498_wen;
  logic [31:0] f498_wdata;
  logic [0:0] f498_clk;
  logic [0:0] f498_rst;
  logic [31:0] f498_rdata;
  sr_buffer_32_1 f498(.wen(f498_wen), .wdata(f498_wdata), .clk(f498_clk), .rst(f498_rst), .rdata(f498_rdata));
  assign f498_clk = clk;
  assign f498_rst = rst;
  // Bindings to f498

  // f500
  logic [0:0] f500_wen;
  logic [31:0] f500_wdata;
  logic [0:0] f500_clk;
  logic [0:0] f500_rst;
  logic [31:0] f500_rdata;
  sr_buffer_32_1 f500(.wen(f500_wen), .wdata(f500_wdata), .clk(f500_clk), .rst(f500_rst), .rdata(f500_rdata));
  assign f500_clk = clk;
  assign f500_rst = rst;
  // Bindings to f500

  // f502
  logic [0:0] f502_wen;
  logic [31:0] f502_wdata;
  logic [0:0] f502_clk;
  logic [0:0] f502_rst;
  logic [31:0] f502_rdata;
  sr_buffer_32_1 f502(.wen(f502_wen), .wdata(f502_wdata), .clk(f502_clk), .rst(f502_rst), .rdata(f502_rdata));
  assign f502_clk = clk;
  assign f502_rst = rst;
  // Bindings to f502

  // f504
  logic [0:0] f504_wen;
  logic [31:0] f504_wdata;
  logic [0:0] f504_clk;
  logic [0:0] f504_rst;
  logic [31:0] f504_rdata;
  sr_buffer_32_1 f504(.wen(f504_wen), .wdata(f504_wdata), .clk(f504_clk), .rst(f504_rst), .rdata(f504_rdata));
  assign f504_clk = clk;
  assign f504_rst = rst;
  // Bindings to f504

  // f506
  logic [0:0] f506_wen;
  logic [31:0] f506_wdata;
  logic [0:0] f506_clk;
  logic [0:0] f506_rst;
  logic [31:0] f506_rdata;
  sr_buffer_32_1 f506(.wen(f506_wen), .wdata(f506_wdata), .clk(f506_clk), .rst(f506_rst), .rdata(f506_rdata));
  assign f506_clk = clk;
  assign f506_rst = rst;
  // Bindings to f506

  // f508
  logic [0:0] f508_wen;
  logic [31:0] f508_wdata;
  logic [0:0] f508_clk;
  logic [0:0] f508_rst;
  logic [31:0] f508_rdata;
  sr_buffer_32_1 f508(.wen(f508_wen), .wdata(f508_wdata), .clk(f508_clk), .rst(f508_rst), .rdata(f508_rdata));
  assign f508_clk = clk;
  assign f508_rst = rst;
  // Bindings to f508

  // f510
  logic [0:0] f510_wen;
  logic [31:0] f510_wdata;
  logic [0:0] f510_clk;
  logic [0:0] f510_rst;
  logic [31:0] f510_rdata;
  sr_buffer_32_1 f510(.wen(f510_wen), .wdata(f510_wdata), .clk(f510_clk), .rst(f510_rst), .rdata(f510_rdata));
  assign f510_clk = clk;
  assign f510_rst = rst;
  // Bindings to f510

  // f512
  logic [0:0] f512_wen;
  logic [31:0] f512_wdata;
  logic [0:0] f512_clk;
  logic [0:0] f512_rst;
  logic [31:0] f512_rdata;
  sr_buffer_32_1 f512(.wen(f512_wen), .wdata(f512_wdata), .clk(f512_clk), .rst(f512_rst), .rdata(f512_rdata));
  assign f512_clk = clk;
  assign f512_rst = rst;
  // Bindings to f512

  // f514
  logic [0:0] f514_wen;
  logic [31:0] f514_wdata;
  logic [0:0] f514_clk;
  logic [0:0] f514_rst;
  logic [31:0] f514_rdata;
  sr_buffer_32_1 f514(.wen(f514_wen), .wdata(f514_wdata), .clk(f514_clk), .rst(f514_rst), .rdata(f514_rdata));
  assign f514_clk = clk;
  assign f514_rst = rst;
  // Bindings to f514

  // f516
  logic [0:0] f516_wen;
  logic [31:0] f516_wdata;
  logic [0:0] f516_clk;
  logic [0:0] f516_rst;
  logic [31:0] f516_rdata;
  sr_buffer_32_1 f516(.wen(f516_wen), .wdata(f516_wdata), .clk(f516_clk), .rst(f516_rst), .rdata(f516_rdata));
  assign f516_clk = clk;
  assign f516_rst = rst;
  // Bindings to f516

  // f518
  logic [0:0] f518_wen;
  logic [31:0] f518_wdata;
  logic [0:0] f518_clk;
  logic [0:0] f518_rst;
  logic [31:0] f518_rdata;
  sr_buffer_32_1 f518(.wen(f518_wen), .wdata(f518_wdata), .clk(f518_clk), .rst(f518_rst), .rdata(f518_rdata));
  assign f518_clk = clk;
  assign f518_rst = rst;
  // Bindings to f518

  // f520
  logic [0:0] f520_wen;
  logic [31:0] f520_wdata;
  logic [0:0] f520_clk;
  logic [0:0] f520_rst;
  logic [31:0] f520_rdata;
  sr_buffer_32_1 f520(.wen(f520_wen), .wdata(f520_wdata), .clk(f520_clk), .rst(f520_rst), .rdata(f520_rdata));
  assign f520_clk = clk;
  assign f520_rst = rst;
  // Bindings to f520

  // f522
  logic [0:0] f522_wen;
  logic [31:0] f522_wdata;
  logic [0:0] f522_clk;
  logic [0:0] f522_rst;
  logic [31:0] f522_rdata;
  sr_buffer_32_1 f522(.wen(f522_wen), .wdata(f522_wdata), .clk(f522_clk), .rst(f522_rst), .rdata(f522_rdata));
  assign f522_clk = clk;
  assign f522_rst = rst;
  // Bindings to f522

  // f524
  logic [0:0] f524_wen;
  logic [31:0] f524_wdata;
  logic [0:0] f524_clk;
  logic [0:0] f524_rst;
  logic [31:0] f524_rdata;
  sr_buffer_32_1 f524(.wen(f524_wen), .wdata(f524_wdata), .clk(f524_clk), .rst(f524_rst), .rdata(f524_rdata));
  assign f524_clk = clk;
  assign f524_rst = rst;
  // Bindings to f524

  // f526
  logic [0:0] f526_wen;
  logic [31:0] f526_wdata;
  logic [0:0] f526_clk;
  logic [0:0] f526_rst;
  logic [31:0] f526_rdata;
  sr_buffer_32_1 f526(.wen(f526_wen), .wdata(f526_wdata), .clk(f526_clk), .rst(f526_rst), .rdata(f526_rdata));
  assign f526_clk = clk;
  assign f526_rst = rst;
  // Bindings to f526

  // f528
  logic [0:0] f528_wen;
  logic [31:0] f528_wdata;
  logic [0:0] f528_clk;
  logic [0:0] f528_rst;
  logic [31:0] f528_rdata;
  sr_buffer_32_1 f528(.wen(f528_wen), .wdata(f528_wdata), .clk(f528_clk), .rst(f528_rst), .rdata(f528_rdata));
  assign f528_clk = clk;
  assign f528_rst = rst;
  // Bindings to f528

  // f530
  logic [0:0] f530_wen;
  logic [31:0] f530_wdata;
  logic [0:0] f530_clk;
  logic [0:0] f530_rst;
  logic [31:0] f530_rdata;
  sr_buffer_32_1 f530(.wen(f530_wen), .wdata(f530_wdata), .clk(f530_clk), .rst(f530_rst), .rdata(f530_rdata));
  assign f530_clk = clk;
  assign f530_rst = rst;
  // Bindings to f530

  // f532
  logic [0:0] f532_wen;
  logic [31:0] f532_wdata;
  logic [0:0] f532_clk;
  logic [0:0] f532_rst;
  logic [31:0] f532_rdata;
  sr_buffer_32_1 f532(.wen(f532_wen), .wdata(f532_wdata), .clk(f532_clk), .rst(f532_rst), .rdata(f532_rdata));
  assign f532_clk = clk;
  assign f532_rst = rst;
  // Bindings to f532

  // f534
  logic [0:0] f534_wen;
  logic [31:0] f534_wdata;
  logic [0:0] f534_clk;
  logic [0:0] f534_rst;
  logic [31:0] f534_rdata;
  sr_buffer_32_1 f534(.wen(f534_wen), .wdata(f534_wdata), .clk(f534_clk), .rst(f534_rst), .rdata(f534_rdata));
  assign f534_clk = clk;
  assign f534_rst = rst;
  // Bindings to f534

  // f536
  logic [0:0] f536_wen;
  logic [31:0] f536_wdata;
  logic [0:0] f536_clk;
  logic [0:0] f536_rst;
  logic [31:0] f536_rdata;
  sr_buffer_32_1 f536(.wen(f536_wen), .wdata(f536_wdata), .clk(f536_clk), .rst(f536_rst), .rdata(f536_rdata));
  assign f536_clk = clk;
  assign f536_rst = rst;
  // Bindings to f536

  // f538
  logic [0:0] f538_wen;
  logic [31:0] f538_wdata;
  logic [0:0] f538_clk;
  logic [0:0] f538_rst;
  logic [31:0] f538_rdata;
  sr_buffer_32_1 f538(.wen(f538_wen), .wdata(f538_wdata), .clk(f538_clk), .rst(f538_rst), .rdata(f538_rdata));
  assign f538_clk = clk;
  assign f538_rst = rst;
  // Bindings to f538

  // f540
  logic [0:0] f540_wen;
  logic [31:0] f540_wdata;
  logic [0:0] f540_clk;
  logic [0:0] f540_rst;
  logic [31:0] f540_rdata;
  sr_buffer_32_1 f540(.wen(f540_wen), .wdata(f540_wdata), .clk(f540_clk), .rst(f540_rst), .rdata(f540_rdata));
  assign f540_clk = clk;
  assign f540_rst = rst;
  // Bindings to f540

  // f542
  logic [0:0] f542_wen;
  logic [31:0] f542_wdata;
  logic [0:0] f542_clk;
  logic [0:0] f542_rst;
  logic [31:0] f542_rdata;
  sr_buffer_32_1 f542(.wen(f542_wen), .wdata(f542_wdata), .clk(f542_clk), .rst(f542_rst), .rdata(f542_rdata));
  assign f542_clk = clk;
  assign f542_rst = rst;
  // Bindings to f542

  // f544
  logic [0:0] f544_wen;
  logic [31:0] f544_wdata;
  logic [0:0] f544_clk;
  logic [0:0] f544_rst;
  logic [31:0] f544_rdata;
  sr_buffer_32_1 f544(.wen(f544_wen), .wdata(f544_wdata), .clk(f544_clk), .rst(f544_rst), .rdata(f544_rdata));
  assign f544_clk = clk;
  assign f544_rst = rst;
  // Bindings to f544

  // f546
  logic [0:0] f546_wen;
  logic [31:0] f546_wdata;
  logic [0:0] f546_clk;
  logic [0:0] f546_rst;
  logic [31:0] f546_rdata;
  sr_buffer_32_1 f546(.wen(f546_wen), .wdata(f546_wdata), .clk(f546_clk), .rst(f546_rst), .rdata(f546_rdata));
  assign f546_clk = clk;
  assign f546_rst = rst;
  // Bindings to f546

  // f548
  logic [0:0] f548_wen;
  logic [31:0] f548_wdata;
  logic [0:0] f548_clk;
  logic [0:0] f548_rst;
  logic [31:0] f548_rdata;
  sr_buffer_32_1 f548(.wen(f548_wen), .wdata(f548_wdata), .clk(f548_clk), .rst(f548_rst), .rdata(f548_rdata));
  assign f548_clk = clk;
  assign f548_rst = rst;
  // Bindings to f548

  // f550
  logic [0:0] f550_wen;
  logic [31:0] f550_wdata;
  logic [0:0] f550_clk;
  logic [0:0] f550_rst;
  logic [31:0] f550_rdata;
  sr_buffer_32_1 f550(.wen(f550_wen), .wdata(f550_wdata), .clk(f550_clk), .rst(f550_rst), .rdata(f550_rdata));
  assign f550_clk = clk;
  assign f550_rst = rst;
  // Bindings to f550

  // f552
  logic [0:0] f552_wen;
  logic [31:0] f552_wdata;
  logic [0:0] f552_clk;
  logic [0:0] f552_rst;
  logic [31:0] f552_rdata;
  sr_buffer_32_1 f552(.wen(f552_wen), .wdata(f552_wdata), .clk(f552_clk), .rst(f552_rst), .rdata(f552_rdata));
  assign f552_clk = clk;
  assign f552_rst = rst;
  // Bindings to f552

  // f554
  logic [0:0] f554_wen;
  logic [31:0] f554_wdata;
  logic [0:0] f554_clk;
  logic [0:0] f554_rst;
  logic [31:0] f554_rdata;
  sr_buffer_32_1 f554(.wen(f554_wen), .wdata(f554_wdata), .clk(f554_clk), .rst(f554_rst), .rdata(f554_rdata));
  assign f554_clk = clk;
  assign f554_rst = rst;
  // Bindings to f554

  // f556
  logic [0:0] f556_wen;
  logic [31:0] f556_wdata;
  logic [0:0] f556_clk;
  logic [0:0] f556_rst;
  logic [31:0] f556_rdata;
  sr_buffer_32_1 f556(.wen(f556_wen), .wdata(f556_wdata), .clk(f556_clk), .rst(f556_rst), .rdata(f556_rdata));
  assign f556_clk = clk;
  assign f556_rst = rst;
  // Bindings to f556

  // f558
  logic [0:0] f558_wen;
  logic [31:0] f558_wdata;
  logic [0:0] f558_clk;
  logic [0:0] f558_rst;
  logic [31:0] f558_rdata;
  sr_buffer_32_1 f558(.wen(f558_wen), .wdata(f558_wdata), .clk(f558_clk), .rst(f558_rst), .rdata(f558_rdata));
  assign f558_clk = clk;
  assign f558_rst = rst;
  // Bindings to f558

  // f560
  logic [0:0] f560_wen;
  logic [31:0] f560_wdata;
  logic [0:0] f560_clk;
  logic [0:0] f560_rst;
  logic [31:0] f560_rdata;
  sr_buffer_32_1 f560(.wen(f560_wen), .wdata(f560_wdata), .clk(f560_clk), .rst(f560_rst), .rdata(f560_rdata));
  assign f560_clk = clk;
  assign f560_rst = rst;
  // Bindings to f560

  // f562
  logic [0:0] f562_wen;
  logic [31:0] f562_wdata;
  logic [0:0] f562_clk;
  logic [0:0] f562_rst;
  logic [31:0] f562_rdata;
  sr_buffer_32_1 f562(.wen(f562_wen), .wdata(f562_wdata), .clk(f562_clk), .rst(f562_rst), .rdata(f562_rdata));
  assign f562_clk = clk;
  assign f562_rst = rst;
  // Bindings to f562

  // f564
  logic [0:0] f564_wen;
  logic [31:0] f564_wdata;
  logic [0:0] f564_clk;
  logic [0:0] f564_rst;
  logic [31:0] f564_rdata;
  sr_buffer_32_1 f564(.wen(f564_wen), .wdata(f564_wdata), .clk(f564_clk), .rst(f564_rst), .rdata(f564_rdata));
  assign f564_clk = clk;
  assign f564_rst = rst;
  // Bindings to f564

  // f566
  logic [0:0] f566_wen;
  logic [31:0] f566_wdata;
  logic [0:0] f566_clk;
  logic [0:0] f566_rst;
  logic [31:0] f566_rdata;
  sr_buffer_32_1 f566(.wen(f566_wen), .wdata(f566_wdata), .clk(f566_clk), .rst(f566_rst), .rdata(f566_rdata));
  assign f566_clk = clk;
  assign f566_rst = rst;
  // Bindings to f566

  // f568
  logic [0:0] f568_wen;
  logic [31:0] f568_wdata;
  logic [0:0] f568_clk;
  logic [0:0] f568_rst;
  logic [31:0] f568_rdata;
  sr_buffer_32_1 f568(.wen(f568_wen), .wdata(f568_wdata), .clk(f568_clk), .rst(f568_rst), .rdata(f568_rdata));
  assign f568_clk = clk;
  assign f568_rst = rst;
  // Bindings to f568

  // f570
  logic [0:0] f570_wen;
  logic [31:0] f570_wdata;
  logic [0:0] f570_clk;
  logic [0:0] f570_rst;
  logic [31:0] f570_rdata;
  sr_buffer_32_1 f570(.wen(f570_wen), .wdata(f570_wdata), .clk(f570_clk), .rst(f570_rst), .rdata(f570_rdata));
  assign f570_clk = clk;
  assign f570_rst = rst;
  // Bindings to f570

  // f572
  logic [0:0] f572_wen;
  logic [31:0] f572_wdata;
  logic [0:0] f572_clk;
  logic [0:0] f572_rst;
  logic [31:0] f572_rdata;
  sr_buffer_32_1 f572(.wen(f572_wen), .wdata(f572_wdata), .clk(f572_clk), .rst(f572_rst), .rdata(f572_rdata));
  assign f572_clk = clk;
  assign f572_rst = rst;
  // Bindings to f572

  // f574
  logic [0:0] f574_wen;
  logic [31:0] f574_wdata;
  logic [0:0] f574_clk;
  logic [0:0] f574_rst;
  logic [31:0] f574_rdata;
  sr_buffer_32_1 f574(.wen(f574_wen), .wdata(f574_wdata), .clk(f574_clk), .rst(f574_rst), .rdata(f574_rdata));
  assign f574_clk = clk;
  assign f574_rst = rst;
  // Bindings to f574

  // f576
  logic [0:0] f576_wen;
  logic [31:0] f576_wdata;
  logic [0:0] f576_clk;
  logic [0:0] f576_rst;
  logic [31:0] f576_rdata;
  sr_buffer_32_1 f576(.wen(f576_wen), .wdata(f576_wdata), .clk(f576_clk), .rst(f576_rst), .rdata(f576_rdata));
  assign f576_clk = clk;
  assign f576_rst = rst;
  // Bindings to f576

  // f578
  logic [0:0] f578_wen;
  logic [31:0] f578_wdata;
  logic [0:0] f578_clk;
  logic [0:0] f578_rst;
  logic [31:0] f578_rdata;
  sr_buffer_32_1 f578(.wen(f578_wen), .wdata(f578_wdata), .clk(f578_clk), .rst(f578_rst), .rdata(f578_rdata));
  assign f578_clk = clk;
  assign f578_rst = rst;
  // Bindings to f578

  // f580
  logic [0:0] f580_wen;
  logic [31:0] f580_wdata;
  logic [0:0] f580_clk;
  logic [0:0] f580_rst;
  logic [31:0] f580_rdata;
  sr_buffer_32_1 f580(.wen(f580_wen), .wdata(f580_wdata), .clk(f580_clk), .rst(f580_rst), .rdata(f580_rdata));
  assign f580_clk = clk;
  assign f580_rst = rst;
  // Bindings to f580

  // f582
  logic [0:0] f582_wen;
  logic [31:0] f582_wdata;
  logic [0:0] f582_clk;
  logic [0:0] f582_rst;
  logic [31:0] f582_rdata;
  sr_buffer_32_1 f582(.wen(f582_wen), .wdata(f582_wdata), .clk(f582_clk), .rst(f582_rst), .rdata(f582_rdata));
  assign f582_clk = clk;
  assign f582_rst = rst;
  // Bindings to f582

  // f584
  logic [0:0] f584_wen;
  logic [31:0] f584_wdata;
  logic [0:0] f584_clk;
  logic [0:0] f584_rst;
  logic [31:0] f584_rdata;
  sr_buffer_32_1 f584(.wen(f584_wen), .wdata(f584_wdata), .clk(f584_clk), .rst(f584_rst), .rdata(f584_rdata));
  assign f584_clk = clk;
  assign f584_rst = rst;
  // Bindings to f584

  // f586
  logic [0:0] f586_wen;
  logic [31:0] f586_wdata;
  logic [0:0] f586_clk;
  logic [0:0] f586_rst;
  logic [31:0] f586_rdata;
  sr_buffer_32_1 f586(.wen(f586_wen), .wdata(f586_wdata), .clk(f586_clk), .rst(f586_rst), .rdata(f586_rdata));
  assign f586_clk = clk;
  assign f586_rst = rst;
  // Bindings to f586

  // f588
  logic [0:0] f588_wen;
  logic [31:0] f588_wdata;
  logic [0:0] f588_clk;
  logic [0:0] f588_rst;
  logic [31:0] f588_rdata;
  sr_buffer_32_1 f588(.wen(f588_wen), .wdata(f588_wdata), .clk(f588_clk), .rst(f588_rst), .rdata(f588_rdata));
  assign f588_clk = clk;
  assign f588_rst = rst;
  // Bindings to f588

  // f590
  logic [0:0] f590_wen;
  logic [31:0] f590_wdata;
  logic [0:0] f590_clk;
  logic [0:0] f590_rst;
  logic [31:0] f590_rdata;
  sr_buffer_32_1 f590(.wen(f590_wen), .wdata(f590_wdata), .clk(f590_clk), .rst(f590_rst), .rdata(f590_rdata));
  assign f590_clk = clk;
  assign f590_rst = rst;
  // Bindings to f590

  // f592
  logic [0:0] f592_wen;
  logic [31:0] f592_wdata;
  logic [0:0] f592_clk;
  logic [0:0] f592_rst;
  logic [31:0] f592_rdata;
  sr_buffer_32_1 f592(.wen(f592_wen), .wdata(f592_wdata), .clk(f592_clk), .rst(f592_rst), .rdata(f592_rdata));
  assign f592_clk = clk;
  assign f592_rst = rst;
  // Bindings to f592

  // f594
  logic [0:0] f594_wen;
  logic [31:0] f594_wdata;
  logic [0:0] f594_clk;
  logic [0:0] f594_rst;
  logic [31:0] f594_rdata;
  sr_buffer_32_1 f594(.wen(f594_wen), .wdata(f594_wdata), .clk(f594_clk), .rst(f594_rst), .rdata(f594_rdata));
  assign f594_clk = clk;
  assign f594_rst = rst;
  // Bindings to f594

  // f596
  logic [0:0] f596_wen;
  logic [31:0] f596_wdata;
  logic [0:0] f596_clk;
  logic [0:0] f596_rst;
  logic [31:0] f596_rdata;
  sr_buffer_32_1 f596(.wen(f596_wen), .wdata(f596_wdata), .clk(f596_clk), .rst(f596_rst), .rdata(f596_rdata));
  assign f596_clk = clk;
  assign f596_rst = rst;
  // Bindings to f596

  // f598
  logic [0:0] f598_wen;
  logic [31:0] f598_wdata;
  logic [0:0] f598_clk;
  logic [0:0] f598_rst;
  logic [31:0] f598_rdata;
  sr_buffer_32_1 f598(.wen(f598_wen), .wdata(f598_wdata), .clk(f598_clk), .rst(f598_rst), .rdata(f598_rdata));
  assign f598_clk = clk;
  assign f598_rst = rst;
  // Bindings to f598

  // f600
  logic [0:0] f600_wen;
  logic [31:0] f600_wdata;
  logic [0:0] f600_clk;
  logic [0:0] f600_rst;
  logic [31:0] f600_rdata;
  sr_buffer_32_1 f600(.wen(f600_wen), .wdata(f600_wdata), .clk(f600_clk), .rst(f600_rst), .rdata(f600_rdata));
  assign f600_clk = clk;
  assign f600_rst = rst;
  // Bindings to f600

  // f602
  logic [0:0] f602_wen;
  logic [31:0] f602_wdata;
  logic [0:0] f602_clk;
  logic [0:0] f602_rst;
  logic [31:0] f602_rdata;
  sr_buffer_32_1 f602(.wen(f602_wen), .wdata(f602_wdata), .clk(f602_clk), .rst(f602_rst), .rdata(f602_rdata));
  assign f602_clk = clk;
  assign f602_rst = rst;
  // Bindings to f602

  // f604
  logic [0:0] f604_wen;
  logic [31:0] f604_wdata;
  logic [0:0] f604_clk;
  logic [0:0] f604_rst;
  logic [31:0] f604_rdata;
  sr_buffer_32_1 f604(.wen(f604_wen), .wdata(f604_wdata), .clk(f604_clk), .rst(f604_rst), .rdata(f604_rdata));
  assign f604_clk = clk;
  assign f604_rst = rst;
  // Bindings to f604

  // f606
  logic [0:0] f606_wen;
  logic [31:0] f606_wdata;
  logic [0:0] f606_clk;
  logic [0:0] f606_rst;
  logic [31:0] f606_rdata;
  sr_buffer_32_1 f606(.wen(f606_wen), .wdata(f606_wdata), .clk(f606_clk), .rst(f606_rst), .rdata(f606_rdata));
  assign f606_clk = clk;
  assign f606_rst = rst;
  // Bindings to f606

  // f608
  logic [0:0] f608_wen;
  logic [31:0] f608_wdata;
  logic [0:0] f608_clk;
  logic [0:0] f608_rst;
  logic [31:0] f608_rdata;
  sr_buffer_32_1 f608(.wen(f608_wen), .wdata(f608_wdata), .clk(f608_clk), .rst(f608_rst), .rdata(f608_rdata));
  assign f608_clk = clk;
  assign f608_rst = rst;
  // Bindings to f608

  // f610
  logic [0:0] f610_wen;
  logic [31:0] f610_wdata;
  logic [0:0] f610_clk;
  logic [0:0] f610_rst;
  logic [31:0] f610_rdata;
  sr_buffer_32_1 f610(.wen(f610_wen), .wdata(f610_wdata), .clk(f610_clk), .rst(f610_rst), .rdata(f610_rdata));
  assign f610_clk = clk;
  assign f610_rst = rst;
  // Bindings to f610

  // f612
  logic [0:0] f612_wen;
  logic [31:0] f612_wdata;
  logic [0:0] f612_clk;
  logic [0:0] f612_rst;
  logic [31:0] f612_rdata;
  sr_buffer_32_1 f612(.wen(f612_wen), .wdata(f612_wdata), .clk(f612_clk), .rst(f612_rst), .rdata(f612_rdata));
  assign f612_clk = clk;
  assign f612_rst = rst;
  // Bindings to f612

  // f614
  logic [0:0] f614_wen;
  logic [31:0] f614_wdata;
  logic [0:0] f614_clk;
  logic [0:0] f614_rst;
  logic [31:0] f614_rdata;
  sr_buffer_32_1 f614(.wen(f614_wen), .wdata(f614_wdata), .clk(f614_clk), .rst(f614_rst), .rdata(f614_rdata));
  assign f614_clk = clk;
  assign f614_rst = rst;
  // Bindings to f614

  // f616
  logic [0:0] f616_wen;
  logic [31:0] f616_wdata;
  logic [0:0] f616_clk;
  logic [0:0] f616_rst;
  logic [31:0] f616_rdata;
  sr_buffer_32_1 f616(.wen(f616_wen), .wdata(f616_wdata), .clk(f616_clk), .rst(f616_rst), .rdata(f616_rdata));
  assign f616_clk = clk;
  assign f616_rst = rst;
  // Bindings to f616

  // f618
  logic [0:0] f618_wen;
  logic [31:0] f618_wdata;
  logic [0:0] f618_clk;
  logic [0:0] f618_rst;
  logic [31:0] f618_rdata;
  sr_buffer_32_1 f618(.wen(f618_wen), .wdata(f618_wdata), .clk(f618_clk), .rst(f618_rst), .rdata(f618_rdata));
  assign f618_clk = clk;
  assign f618_rst = rst;
  // Bindings to f618

  // f620
  logic [0:0] f620_wen;
  logic [31:0] f620_wdata;
  logic [0:0] f620_clk;
  logic [0:0] f620_rst;
  logic [31:0] f620_rdata;
  sr_buffer_32_1 f620(.wen(f620_wen), .wdata(f620_wdata), .clk(f620_clk), .rst(f620_rst), .rdata(f620_rdata));
  assign f620_clk = clk;
  assign f620_rst = rst;
  // Bindings to f620

  // f622
  logic [0:0] f622_wen;
  logic [31:0] f622_wdata;
  logic [0:0] f622_clk;
  logic [0:0] f622_rst;
  logic [31:0] f622_rdata;
  sr_buffer_32_1 f622(.wen(f622_wen), .wdata(f622_wdata), .clk(f622_clk), .rst(f622_rst), .rdata(f622_rdata));
  assign f622_clk = clk;
  assign f622_rst = rst;
  // Bindings to f622

  // f624
  logic [0:0] f624_wen;
  logic [31:0] f624_wdata;
  logic [0:0] f624_clk;
  logic [0:0] f624_rst;
  logic [31:0] f624_rdata;
  sr_buffer_32_1 f624(.wen(f624_wen), .wdata(f624_wdata), .clk(f624_clk), .rst(f624_rst), .rdata(f624_rdata));
  assign f624_clk = clk;
  assign f624_rst = rst;
  // Bindings to f624

  // f626
  logic [0:0] f626_wen;
  logic [31:0] f626_wdata;
  logic [0:0] f626_clk;
  logic [0:0] f626_rst;
  logic [31:0] f626_rdata;
  sr_buffer_32_1 f626(.wen(f626_wen), .wdata(f626_wdata), .clk(f626_clk), .rst(f626_rst), .rdata(f626_rdata));
  assign f626_clk = clk;
  assign f626_rst = rst;
  // Bindings to f626

  // f628
  logic [0:0] f628_wen;
  logic [31:0] f628_wdata;
  logic [0:0] f628_clk;
  logic [0:0] f628_rst;
  logic [31:0] f628_rdata;
  sr_buffer_32_1 f628(.wen(f628_wen), .wdata(f628_wdata), .clk(f628_clk), .rst(f628_rst), .rdata(f628_rdata));
  assign f628_clk = clk;
  assign f628_rst = rst;
  // Bindings to f628

  // f630
  logic [0:0] f630_wen;
  logic [31:0] f630_wdata;
  logic [0:0] f630_clk;
  logic [0:0] f630_rst;
  logic [31:0] f630_rdata;
  sr_buffer_32_1 f630(.wen(f630_wen), .wdata(f630_wdata), .clk(f630_clk), .rst(f630_rst), .rdata(f630_rdata));
  assign f630_clk = clk;
  assign f630_rst = rst;
  // Bindings to f630

  // f632
  logic [0:0] f632_wen;
  logic [31:0] f632_wdata;
  logic [0:0] f632_clk;
  logic [0:0] f632_rst;
  logic [31:0] f632_rdata;
  sr_buffer_32_1 f632(.wen(f632_wen), .wdata(f632_wdata), .clk(f632_clk), .rst(f632_rst), .rdata(f632_rdata));
  assign f632_clk = clk;
  assign f632_rst = rst;
  // Bindings to f632

  // f634
  logic [0:0] f634_wen;
  logic [31:0] f634_wdata;
  logic [0:0] f634_clk;
  logic [0:0] f634_rst;
  logic [31:0] f634_rdata;
  sr_buffer_32_1 f634(.wen(f634_wen), .wdata(f634_wdata), .clk(f634_clk), .rst(f634_rst), .rdata(f634_rdata));
  assign f634_clk = clk;
  assign f634_rst = rst;
  // Bindings to f634

  // f636
  logic [0:0] f636_wen;
  logic [31:0] f636_wdata;
  logic [0:0] f636_clk;
  logic [0:0] f636_rst;
  logic [31:0] f636_rdata;
  sr_buffer_32_1 f636(.wen(f636_wen), .wdata(f636_wdata), .clk(f636_clk), .rst(f636_rst), .rdata(f636_rdata));
  assign f636_clk = clk;
  assign f636_rst = rst;
  // Bindings to f636

  // f638
  logic [0:0] f638_wen;
  logic [31:0] f638_wdata;
  logic [0:0] f638_clk;
  logic [0:0] f638_rst;
  logic [31:0] f638_rdata;
  sr_buffer_32_1 f638(.wen(f638_wen), .wdata(f638_wdata), .clk(f638_clk), .rst(f638_rst), .rdata(f638_rdata));
  assign f638_clk = clk;
  assign f638_rst = rst;
  // Bindings to f638

  // f640
  logic [0:0] f640_wen;
  logic [31:0] f640_wdata;
  logic [0:0] f640_clk;
  logic [0:0] f640_rst;
  logic [31:0] f640_rdata;
  sr_buffer_32_1 f640(.wen(f640_wen), .wdata(f640_wdata), .clk(f640_clk), .rst(f640_rst), .rdata(f640_rdata));
  assign f640_clk = clk;
  assign f640_rst = rst;
  // Bindings to f640

  // f642
  logic [0:0] f642_wen;
  logic [31:0] f642_wdata;
  logic [0:0] f642_clk;
  logic [0:0] f642_rst;
  logic [31:0] f642_rdata;
  sr_buffer_32_1 f642(.wen(f642_wen), .wdata(f642_wdata), .clk(f642_clk), .rst(f642_rst), .rdata(f642_rdata));
  assign f642_clk = clk;
  assign f642_rst = rst;
  // Bindings to f642

  // f644
  logic [0:0] f644_wen;
  logic [31:0] f644_wdata;
  logic [0:0] f644_clk;
  logic [0:0] f644_rst;
  logic [31:0] f644_rdata;
  sr_buffer_32_1 f644(.wen(f644_wen), .wdata(f644_wdata), .clk(f644_clk), .rst(f644_rst), .rdata(f644_rdata));
  assign f644_clk = clk;
  assign f644_rst = rst;
  // Bindings to f644

  // f646
  logic [0:0] f646_wen;
  logic [31:0] f646_wdata;
  logic [0:0] f646_clk;
  logic [0:0] f646_rst;
  logic [31:0] f646_rdata;
  sr_buffer_32_1 f646(.wen(f646_wen), .wdata(f646_wdata), .clk(f646_clk), .rst(f646_rst), .rdata(f646_rdata));
  assign f646_clk = clk;
  assign f646_rst = rst;
  // Bindings to f646

  // f648
  logic [0:0] f648_wen;
  logic [31:0] f648_wdata;
  logic [0:0] f648_clk;
  logic [0:0] f648_rst;
  logic [31:0] f648_rdata;
  sr_buffer_32_1 f648(.wen(f648_wen), .wdata(f648_wdata), .clk(f648_clk), .rst(f648_rst), .rdata(f648_rdata));
  assign f648_clk = clk;
  assign f648_rst = rst;
  // Bindings to f648

  // f650
  logic [0:0] f650_wen;
  logic [31:0] f650_wdata;
  logic [0:0] f650_clk;
  logic [0:0] f650_rst;
  logic [31:0] f650_rdata;
  sr_buffer_32_1 f650(.wen(f650_wen), .wdata(f650_wdata), .clk(f650_clk), .rst(f650_rst), .rdata(f650_rdata));
  assign f650_clk = clk;
  assign f650_rst = rst;
  // Bindings to f650

  // f652
  logic [0:0] f652_wen;
  logic [31:0] f652_wdata;
  logic [0:0] f652_clk;
  logic [0:0] f652_rst;
  logic [31:0] f652_rdata;
  sr_buffer_32_1 f652(.wen(f652_wen), .wdata(f652_wdata), .clk(f652_clk), .rst(f652_rst), .rdata(f652_rdata));
  assign f652_clk = clk;
  assign f652_rst = rst;
  // Bindings to f652

  // f654
  logic [0:0] f654_wen;
  logic [31:0] f654_wdata;
  logic [0:0] f654_clk;
  logic [0:0] f654_rst;
  logic [31:0] f654_rdata;
  sr_buffer_32_1 f654(.wen(f654_wen), .wdata(f654_wdata), .clk(f654_clk), .rst(f654_rst), .rdata(f654_rdata));
  assign f654_clk = clk;
  assign f654_rst = rst;
  // Bindings to f654

  // f656
  logic [0:0] f656_wen;
  logic [31:0] f656_wdata;
  logic [0:0] f656_clk;
  logic [0:0] f656_rst;
  logic [31:0] f656_rdata;
  sr_buffer_32_1 f656(.wen(f656_wen), .wdata(f656_wdata), .clk(f656_clk), .rst(f656_rst), .rdata(f656_rdata));
  assign f656_clk = clk;
  assign f656_rst = rst;
  // Bindings to f656

  // f658
  logic [0:0] f658_wen;
  logic [31:0] f658_wdata;
  logic [0:0] f658_clk;
  logic [0:0] f658_rst;
  logic [31:0] f658_rdata;
  sr_buffer_32_1 f658(.wen(f658_wen), .wdata(f658_wdata), .clk(f658_clk), .rst(f658_rst), .rdata(f658_rdata));
  assign f658_clk = clk;
  assign f658_rst = rst;
  // Bindings to f658

  // f660
  logic [0:0] f660_wen;
  logic [31:0] f660_wdata;
  logic [0:0] f660_clk;
  logic [0:0] f660_rst;
  logic [31:0] f660_rdata;
  sr_buffer_32_1 f660(.wen(f660_wen), .wdata(f660_wdata), .clk(f660_clk), .rst(f660_rst), .rdata(f660_rdata));
  assign f660_clk = clk;
  assign f660_rst = rst;
  // Bindings to f660

  // f662
  logic [0:0] f662_wen;
  logic [31:0] f662_wdata;
  logic [0:0] f662_clk;
  logic [0:0] f662_rst;
  logic [31:0] f662_rdata;
  sr_buffer_32_1 f662(.wen(f662_wen), .wdata(f662_wdata), .clk(f662_clk), .rst(f662_rst), .rdata(f662_rdata));
  assign f662_clk = clk;
  assign f662_rst = rst;
  // Bindings to f662

  // f664
  logic [0:0] f664_wen;
  logic [31:0] f664_wdata;
  logic [0:0] f664_clk;
  logic [0:0] f664_rst;
  logic [31:0] f664_rdata;
  sr_buffer_32_1 f664(.wen(f664_wen), .wdata(f664_wdata), .clk(f664_clk), .rst(f664_rst), .rdata(f664_rdata));
  assign f664_clk = clk;
  assign f664_rst = rst;
  // Bindings to f664

  // f666
  logic [0:0] f666_wen;
  logic [31:0] f666_wdata;
  logic [0:0] f666_clk;
  logic [0:0] f666_rst;
  logic [31:0] f666_rdata;
  sr_buffer_32_1 f666(.wen(f666_wen), .wdata(f666_wdata), .clk(f666_clk), .rst(f666_rst), .rdata(f666_rdata));
  assign f666_clk = clk;
  assign f666_rst = rst;
  // Bindings to f666

  // f668
  logic [0:0] f668_wen;
  logic [31:0] f668_wdata;
  logic [0:0] f668_clk;
  logic [0:0] f668_rst;
  logic [31:0] f668_rdata;
  sr_buffer_32_1 f668(.wen(f668_wen), .wdata(f668_wdata), .clk(f668_clk), .rst(f668_rst), .rdata(f668_rdata));
  assign f668_clk = clk;
  assign f668_rst = rst;
  // Bindings to f668

  // f670
  logic [0:0] f670_wen;
  logic [31:0] f670_wdata;
  logic [0:0] f670_clk;
  logic [0:0] f670_rst;
  logic [31:0] f670_rdata;
  sr_buffer_32_1 f670(.wen(f670_wen), .wdata(f670_wdata), .clk(f670_clk), .rst(f670_rst), .rdata(f670_rdata));
  assign f670_clk = clk;
  assign f670_rst = rst;
  // Bindings to f670

  // f672
  logic [0:0] f672_wen;
  logic [31:0] f672_wdata;
  logic [0:0] f672_clk;
  logic [0:0] f672_rst;
  logic [31:0] f672_rdata;
  sr_buffer_32_1 f672(.wen(f672_wen), .wdata(f672_wdata), .clk(f672_clk), .rst(f672_rst), .rdata(f672_rdata));
  assign f672_clk = clk;
  assign f672_rst = rst;
  // Bindings to f672

  // f674
  logic [0:0] f674_wen;
  logic [31:0] f674_wdata;
  logic [0:0] f674_clk;
  logic [0:0] f674_rst;
  logic [31:0] f674_rdata;
  sr_buffer_32_1 f674(.wen(f674_wen), .wdata(f674_wdata), .clk(f674_clk), .rst(f674_rst), .rdata(f674_rdata));
  assign f674_clk = clk;
  assign f674_rst = rst;
  // Bindings to f674

  // f676
  logic [0:0] f676_wen;
  logic [31:0] f676_wdata;
  logic [0:0] f676_clk;
  logic [0:0] f676_rst;
  logic [31:0] f676_rdata;
  sr_buffer_32_1 f676(.wen(f676_wen), .wdata(f676_wdata), .clk(f676_clk), .rst(f676_rst), .rdata(f676_rdata));
  assign f676_clk = clk;
  assign f676_rst = rst;
  // Bindings to f676

  // f678
  logic [0:0] f678_wen;
  logic [31:0] f678_wdata;
  logic [0:0] f678_clk;
  logic [0:0] f678_rst;
  logic [31:0] f678_rdata;
  sr_buffer_32_1 f678(.wen(f678_wen), .wdata(f678_wdata), .clk(f678_clk), .rst(f678_rst), .rdata(f678_rdata));
  assign f678_clk = clk;
  assign f678_rst = rst;
  // Bindings to f678

  // f680
  logic [0:0] f680_wen;
  logic [31:0] f680_wdata;
  logic [0:0] f680_clk;
  logic [0:0] f680_rst;
  logic [31:0] f680_rdata;
  sr_buffer_32_1 f680(.wen(f680_wen), .wdata(f680_wdata), .clk(f680_clk), .rst(f680_rst), .rdata(f680_rdata));
  assign f680_clk = clk;
  assign f680_rst = rst;
  // Bindings to f680

  // f682
  logic [0:0] f682_wen;
  logic [31:0] f682_wdata;
  logic [0:0] f682_clk;
  logic [0:0] f682_rst;
  logic [31:0] f682_rdata;
  sr_buffer_32_1 f682(.wen(f682_wen), .wdata(f682_wdata), .clk(f682_clk), .rst(f682_rst), .rdata(f682_rdata));
  assign f682_clk = clk;
  assign f682_rst = rst;
  // Bindings to f682

  // f684
  logic [0:0] f684_wen;
  logic [31:0] f684_wdata;
  logic [0:0] f684_clk;
  logic [0:0] f684_rst;
  logic [31:0] f684_rdata;
  sr_buffer_32_1 f684(.wen(f684_wen), .wdata(f684_wdata), .clk(f684_clk), .rst(f684_rst), .rdata(f684_rdata));
  assign f684_clk = clk;
  assign f684_rst = rst;
  // Bindings to f684

  // f686
  logic [0:0] f686_wen;
  logic [31:0] f686_wdata;
  logic [0:0] f686_clk;
  logic [0:0] f686_rst;
  logic [31:0] f686_rdata;
  sr_buffer_32_1 f686(.wen(f686_wen), .wdata(f686_wdata), .clk(f686_clk), .rst(f686_rst), .rdata(f686_rdata));
  assign f686_clk = clk;
  assign f686_rst = rst;
  // Bindings to f686

  // f688
  logic [0:0] f688_wen;
  logic [31:0] f688_wdata;
  logic [0:0] f688_clk;
  logic [0:0] f688_rst;
  logic [31:0] f688_rdata;
  sr_buffer_32_1 f688(.wen(f688_wen), .wdata(f688_wdata), .clk(f688_clk), .rst(f688_rst), .rdata(f688_rdata));
  assign f688_clk = clk;
  assign f688_rst = rst;
  // Bindings to f688

  // f690
  logic [0:0] f690_wen;
  logic [31:0] f690_wdata;
  logic [0:0] f690_clk;
  logic [0:0] f690_rst;
  logic [31:0] f690_rdata;
  sr_buffer_32_1 f690(.wen(f690_wen), .wdata(f690_wdata), .clk(f690_clk), .rst(f690_rst), .rdata(f690_rdata));
  assign f690_clk = clk;
  assign f690_rst = rst;
  // Bindings to f690

  // f692
  logic [0:0] f692_wen;
  logic [31:0] f692_wdata;
  logic [0:0] f692_clk;
  logic [0:0] f692_rst;
  logic [31:0] f692_rdata;
  sr_buffer_32_1 f692(.wen(f692_wen), .wdata(f692_wdata), .clk(f692_clk), .rst(f692_rst), .rdata(f692_rdata));
  assign f692_clk = clk;
  assign f692_rst = rst;
  // Bindings to f692

  // f694
  logic [0:0] f694_wen;
  logic [31:0] f694_wdata;
  logic [0:0] f694_clk;
  logic [0:0] f694_rst;
  logic [31:0] f694_rdata;
  sr_buffer_32_1 f694(.wen(f694_wen), .wdata(f694_wdata), .clk(f694_clk), .rst(f694_rst), .rdata(f694_rdata));
  assign f694_clk = clk;
  assign f694_rst = rst;
  // Bindings to f694

  // f696
  logic [0:0] f696_wen;
  logic [31:0] f696_wdata;
  logic [0:0] f696_clk;
  logic [0:0] f696_rst;
  logic [31:0] f696_rdata;
  sr_buffer_32_1 f696(.wen(f696_wen), .wdata(f696_wdata), .clk(f696_clk), .rst(f696_rst), .rdata(f696_rdata));
  assign f696_clk = clk;
  assign f696_rst = rst;
  // Bindings to f696

  // f698
  logic [0:0] f698_wen;
  logic [31:0] f698_wdata;
  logic [0:0] f698_clk;
  logic [0:0] f698_rst;
  logic [31:0] f698_rdata;
  sr_buffer_32_1 f698(.wen(f698_wen), .wdata(f698_wdata), .clk(f698_clk), .rst(f698_rst), .rdata(f698_rdata));
  assign f698_clk = clk;
  assign f698_rst = rst;
  // Bindings to f698

  // f700
  logic [0:0] f700_wen;
  logic [31:0] f700_wdata;
  logic [0:0] f700_clk;
  logic [0:0] f700_rst;
  logic [31:0] f700_rdata;
  sr_buffer_32_1 f700(.wen(f700_wen), .wdata(f700_wdata), .clk(f700_clk), .rst(f700_rst), .rdata(f700_rdata));
  assign f700_clk = clk;
  assign f700_rst = rst;
  // Bindings to f700

  // f702
  logic [0:0] f702_wen;
  logic [31:0] f702_wdata;
  logic [0:0] f702_clk;
  logic [0:0] f702_rst;
  logic [31:0] f702_rdata;
  sr_buffer_32_1 f702(.wen(f702_wen), .wdata(f702_wdata), .clk(f702_clk), .rst(f702_rst), .rdata(f702_rdata));
  assign f702_clk = clk;
  assign f702_rst = rst;
  // Bindings to f702

  // f768
  logic [0:0] f768_wen;
  logic [31:0] f768_wdata;
  logic [0:0] f768_clk;
  logic [0:0] f768_rst;
  logic [31:0] f768_rdata;
  sr_buffer_32_1 f768(.wen(f768_wen), .wdata(f768_wdata), .clk(f768_clk), .rst(f768_rst), .rdata(f768_rdata));
  assign f768_clk = clk;
  assign f768_rst = rst;
  // Bindings to f768

  // f766
  logic [0:0] f766_wen;
  logic [31:0] f766_wdata;
  logic [0:0] f766_clk;
  logic [0:0] f766_rst;
  logic [31:0] f766_rdata;
  sr_buffer_32_1 f766(.wen(f766_wen), .wdata(f766_wdata), .clk(f766_clk), .rst(f766_rst), .rdata(f766_rdata));
  assign f766_clk = clk;
  assign f766_rst = rst;
  // Bindings to f766

  // f756
  logic [0:0] f756_wen;
  logic [31:0] f756_wdata;
  logic [0:0] f756_clk;
  logic [0:0] f756_rst;
  logic [31:0] f756_rdata;
  sr_buffer_32_1 f756(.wen(f756_wen), .wdata(f756_wdata), .clk(f756_clk), .rst(f756_rst), .rdata(f756_rdata));
  assign f756_clk = clk;
  assign f756_rst = rst;
  // Bindings to f756

  // f764
  logic [0:0] f764_wen;
  logic [31:0] f764_wdata;
  logic [0:0] f764_clk;
  logic [0:0] f764_rst;
  logic [31:0] f764_rdata;
  sr_buffer_32_1 f764(.wen(f764_wen), .wdata(f764_wdata), .clk(f764_clk), .rst(f764_rst), .rdata(f764_rdata));
  assign f764_clk = clk;
  assign f764_rst = rst;
  // Bindings to f764

  // f752
  logic [0:0] f752_wen;
  logic [31:0] f752_wdata;
  logic [0:0] f752_clk;
  logic [0:0] f752_rst;
  logic [31:0] f752_rdata;
  sr_buffer_32_1 f752(.wen(f752_wen), .wdata(f752_wdata), .clk(f752_clk), .rst(f752_rst), .rdata(f752_rdata));
  assign f752_clk = clk;
  assign f752_rst = rst;
  // Bindings to f752

  // f750
  logic [0:0] f750_wen;
  logic [31:0] f750_wdata;
  logic [0:0] f750_clk;
  logic [0:0] f750_rst;
  logic [31:0] f750_rdata;
  sr_buffer_32_1 f750(.wen(f750_wen), .wdata(f750_wdata), .clk(f750_clk), .rst(f750_rst), .rdata(f750_rdata));
  assign f750_clk = clk;
  assign f750_rst = rst;
  // Bindings to f750

  // f744
  logic [0:0] f744_wen;
  logic [31:0] f744_wdata;
  logic [0:0] f744_clk;
  logic [0:0] f744_rst;
  logic [31:0] f744_rdata;
  sr_buffer_32_1 f744(.wen(f744_wen), .wdata(f744_wdata), .clk(f744_clk), .rst(f744_rst), .rdata(f744_rdata));
  assign f744_clk = clk;
  assign f744_rst = rst;
  // Bindings to f744

  // f748
  logic [0:0] f748_wen;
  logic [31:0] f748_wdata;
  logic [0:0] f748_clk;
  logic [0:0] f748_rst;
  logic [31:0] f748_rdata;
  sr_buffer_32_1 f748(.wen(f748_wen), .wdata(f748_wdata), .clk(f748_clk), .rst(f748_rst), .rdata(f748_rdata));
  assign f748_clk = clk;
  assign f748_rst = rst;
  // Bindings to f748

  // f808
  logic [0:0] f808_wen;
  logic [31:0] f808_wdata;
  logic [0:0] f808_clk;
  logic [0:0] f808_rst;
  logic [31:0] f808_rdata;
  sr_buffer_32_1 f808(.wen(f808_wen), .wdata(f808_wdata), .clk(f808_clk), .rst(f808_rst), .rdata(f808_rdata));
  assign f808_clk = clk;
  assign f808_rst = rst;
  // Bindings to f808

  // f816
  logic [0:0] f816_wen;
  logic [31:0] f816_wdata;
  logic [0:0] f816_clk;
  logic [0:0] f816_rst;
  logic [31:0] f816_rdata;
  sr_buffer_32_1 f816(.wen(f816_wen), .wdata(f816_wdata), .clk(f816_clk), .rst(f816_rst), .rdata(f816_rdata));
  assign f816_clk = clk;
  assign f816_rst = rst;
  // Bindings to f816

  // f790
  logic [0:0] f790_wen;
  logic [31:0] f790_wdata;
  logic [0:0] f790_clk;
  logic [0:0] f790_rst;
  logic [31:0] f790_rdata;
  sr_buffer_32_1 f790(.wen(f790_wen), .wdata(f790_wdata), .clk(f790_clk), .rst(f790_rst), .rdata(f790_rdata));
  assign f790_clk = clk;
  assign f790_rst = rst;
  // Bindings to f790

  // f788
  logic [0:0] f788_wen;
  logic [31:0] f788_wdata;
  logic [0:0] f788_clk;
  logic [0:0] f788_rst;
  logic [31:0] f788_rdata;
  sr_buffer_32_1 f788(.wen(f788_wen), .wdata(f788_wdata), .clk(f788_clk), .rst(f788_rst), .rdata(f788_rdata));
  assign f788_clk = clk;
  assign f788_rst = rst;
  // Bindings to f788

  // f786
  logic [0:0] f786_wen;
  logic [31:0] f786_wdata;
  logic [0:0] f786_clk;
  logic [0:0] f786_rst;
  logic [31:0] f786_rdata;
  sr_buffer_32_1 f786(.wen(f786_wen), .wdata(f786_wdata), .clk(f786_clk), .rst(f786_rst), .rdata(f786_rdata));
  assign f786_clk = clk;
  assign f786_rst = rst;
  // Bindings to f786

  // f782
  logic [0:0] f782_wen;
  logic [31:0] f782_wdata;
  logic [0:0] f782_clk;
  logic [0:0] f782_rst;
  logic [31:0] f782_rdata;
  sr_buffer_32_1 f782(.wen(f782_wen), .wdata(f782_wdata), .clk(f782_clk), .rst(f782_rst), .rdata(f782_rdata));
  assign f782_clk = clk;
  assign f782_rst = rst;
  // Bindings to f782

  // f784
  logic [0:0] f784_wen;
  logic [31:0] f784_wdata;
  logic [0:0] f784_clk;
  logic [0:0] f784_rst;
  logic [31:0] f784_rdata;
  sr_buffer_32_1 f784(.wen(f784_wen), .wdata(f784_wdata), .clk(f784_clk), .rst(f784_rst), .rdata(f784_rdata));
  assign f784_clk = clk;
  assign f784_rst = rst;
  // Bindings to f784

  // f780
  logic [0:0] f780_wen;
  logic [31:0] f780_wdata;
  logic [0:0] f780_clk;
  logic [0:0] f780_rst;
  logic [31:0] f780_rdata;
  sr_buffer_32_1 f780(.wen(f780_wen), .wdata(f780_wdata), .clk(f780_clk), .rst(f780_rst), .rdata(f780_rdata));
  assign f780_clk = clk;
  assign f780_rst = rst;
  // Bindings to f780

  // f778
  logic [0:0] f778_wen;
  logic [31:0] f778_wdata;
  logic [0:0] f778_clk;
  logic [0:0] f778_rst;
  logic [31:0] f778_rdata;
  sr_buffer_32_1 f778(.wen(f778_wen), .wdata(f778_wdata), .clk(f778_clk), .rst(f778_rst), .rdata(f778_rdata));
  assign f778_clk = clk;
  assign f778_rst = rst;
  // Bindings to f778

  // f776
  logic [0:0] f776_wen;
  logic [31:0] f776_wdata;
  logic [0:0] f776_clk;
  logic [0:0] f776_rst;
  logic [31:0] f776_rdata;
  sr_buffer_32_1 f776(.wen(f776_wen), .wdata(f776_wdata), .clk(f776_clk), .rst(f776_rst), .rdata(f776_rdata));
  assign f776_clk = clk;
  assign f776_rst = rst;
  // Bindings to f776

  // f774
  logic [0:0] f774_wen;
  logic [31:0] f774_wdata;
  logic [0:0] f774_clk;
  logic [0:0] f774_rst;
  logic [31:0] f774_rdata;
  sr_buffer_32_1 f774(.wen(f774_wen), .wdata(f774_wdata), .clk(f774_clk), .rst(f774_rst), .rdata(f774_rdata));
  assign f774_clk = clk;
  assign f774_rst = rst;
  // Bindings to f774

  // f770
  logic [0:0] f770_wen;
  logic [31:0] f770_wdata;
  logic [0:0] f770_clk;
  logic [0:0] f770_rst;
  logic [31:0] f770_rdata;
  sr_buffer_32_1 f770(.wen(f770_wen), .wdata(f770_wdata), .clk(f770_clk), .rst(f770_rst), .rdata(f770_rdata));
  assign f770_clk = clk;
  assign f770_rst = rst;
  // Bindings to f770

  // f772
  logic [0:0] f772_wen;
  logic [31:0] f772_wdata;
  logic [0:0] f772_clk;
  logic [0:0] f772_rst;
  logic [31:0] f772_rdata;
  sr_buffer_32_1 f772(.wen(f772_wen), .wdata(f772_wdata), .clk(f772_clk), .rst(f772_rst), .rdata(f772_rdata));
  assign f772_clk = clk;
  assign f772_rst = rst;
  // Bindings to f772

  // f830
  logic [0:0] f830_wen;
  logic [31:0] f830_wdata;
  logic [0:0] f830_clk;
  logic [0:0] f830_rst;
  logic [31:0] f830_rdata;
  sr_buffer_32_1 f830(.wen(f830_wen), .wdata(f830_wdata), .clk(f830_clk), .rst(f830_rst), .rdata(f830_rdata));
  assign f830_clk = clk;
  assign f830_rst = rst;
  // Bindings to f830

  // f828
  logic [0:0] f828_wen;
  logic [31:0] f828_wdata;
  logic [0:0] f828_clk;
  logic [0:0] f828_rst;
  logic [31:0] f828_rdata;
  sr_buffer_32_1 f828(.wen(f828_wen), .wdata(f828_wdata), .clk(f828_clk), .rst(f828_rst), .rdata(f828_rdata));
  assign f828_clk = clk;
  assign f828_rst = rst;
  // Bindings to f828

  // f796
  logic [0:0] f796_wen;
  logic [31:0] f796_wdata;
  logic [0:0] f796_clk;
  logic [0:0] f796_rst;
  logic [31:0] f796_rdata;
  sr_buffer_32_1 f796(.wen(f796_wen), .wdata(f796_wdata), .clk(f796_clk), .rst(f796_rst), .rdata(f796_rdata));
  assign f796_clk = clk;
  assign f796_rst = rst;
  // Bindings to f796

  // f826
  logic [0:0] f826_wen;
  logic [31:0] f826_wdata;
  logic [0:0] f826_clk;
  logic [0:0] f826_rst;
  logic [31:0] f826_rdata;
  sr_buffer_32_1 f826(.wen(f826_wen), .wdata(f826_wdata), .clk(f826_clk), .rst(f826_rst), .rdata(f826_rdata));
  assign f826_clk = clk;
  assign f826_rst = rst;
  // Bindings to f826

  // f824
  logic [0:0] f824_wen;
  logic [31:0] f824_wdata;
  logic [0:0] f824_clk;
  logic [0:0] f824_rst;
  logic [31:0] f824_rdata;
  sr_buffer_32_1 f824(.wen(f824_wen), .wdata(f824_wdata), .clk(f824_clk), .rst(f824_rst), .rdata(f824_rdata));
  assign f824_clk = clk;
  assign f824_rst = rst;
  // Bindings to f824

  // f822
  logic [0:0] f822_wen;
  logic [31:0] f822_wdata;
  logic [0:0] f822_clk;
  logic [0:0] f822_rst;
  logic [31:0] f822_rdata;
  sr_buffer_32_1 f822(.wen(f822_wen), .wdata(f822_wdata), .clk(f822_clk), .rst(f822_rst), .rdata(f822_rdata));
  assign f822_clk = clk;
  assign f822_rst = rst;
  // Bindings to f822

  // f820
  logic [0:0] f820_wen;
  logic [31:0] f820_wdata;
  logic [0:0] f820_clk;
  logic [0:0] f820_rst;
  logic [31:0] f820_rdata;
  sr_buffer_32_1 f820(.wen(f820_wen), .wdata(f820_wdata), .clk(f820_clk), .rst(f820_rst), .rdata(f820_rdata));
  assign f820_clk = clk;
  assign f820_rst = rst;
  // Bindings to f820

  // f818
  logic [0:0] f818_wen;
  logic [31:0] f818_wdata;
  logic [0:0] f818_clk;
  logic [0:0] f818_rst;
  logic [31:0] f818_rdata;
  sr_buffer_32_1 f818(.wen(f818_wen), .wdata(f818_wdata), .clk(f818_clk), .rst(f818_rst), .rdata(f818_rdata));
  assign f818_clk = clk;
  assign f818_rst = rst;
  // Bindings to f818

  // f762
  logic [0:0] f762_wen;
  logic [31:0] f762_wdata;
  logic [0:0] f762_clk;
  logic [0:0] f762_rst;
  logic [31:0] f762_rdata;
  sr_buffer_32_1 f762(.wen(f762_wen), .wdata(f762_wdata), .clk(f762_clk), .rst(f762_rst), .rdata(f762_rdata));
  assign f762_clk = clk;
  assign f762_rst = rst;
  // Bindings to f762

  // f758
  logic [0:0] f758_wen;
  logic [31:0] f758_wdata;
  logic [0:0] f758_clk;
  logic [0:0] f758_rst;
  logic [31:0] f758_rdata;
  sr_buffer_32_1 f758(.wen(f758_wen), .wdata(f758_wdata), .clk(f758_clk), .rst(f758_rst), .rdata(f758_rdata));
  assign f758_clk = clk;
  assign f758_rst = rst;
  // Bindings to f758

  // f760
  logic [0:0] f760_wen;
  logic [31:0] f760_wdata;
  logic [0:0] f760_clk;
  logic [0:0] f760_rst;
  logic [31:0] f760_rdata;
  sr_buffer_32_1 f760(.wen(f760_wen), .wdata(f760_wdata), .clk(f760_clk), .rst(f760_rst), .rdata(f760_rdata));
  assign f760_clk = clk;
  assign f760_rst = rst;
  // Bindings to f760

  // f900
  logic [0:0] f900_wen;
  logic [31:0] f900_wdata;
  logic [0:0] f900_clk;
  logic [0:0] f900_rst;
  logic [31:0] f900_rdata;
  sr_buffer_32_1 f900(.wen(f900_wen), .wdata(f900_wdata), .clk(f900_clk), .rst(f900_rst), .rdata(f900_rdata));
  assign f900_clk = clk;
  assign f900_rst = rst;
  // Bindings to f900

  // f890
  logic [0:0] f890_wen;
  logic [31:0] f890_wdata;
  logic [0:0] f890_clk;
  logic [0:0] f890_rst;
  logic [31:0] f890_rdata;
  sr_buffer_32_1 f890(.wen(f890_wen), .wdata(f890_wdata), .clk(f890_clk), .rst(f890_rst), .rdata(f890_rdata));
  assign f890_clk = clk;
  assign f890_rst = rst;
  // Bindings to f890

  // f802
  logic [0:0] f802_wen;
  logic [31:0] f802_wdata;
  logic [0:0] f802_clk;
  logic [0:0] f802_rst;
  logic [31:0] f802_rdata;
  sr_buffer_32_1 f802(.wen(f802_wen), .wdata(f802_wdata), .clk(f802_clk), .rst(f802_rst), .rdata(f802_rdata));
  assign f802_clk = clk;
  assign f802_rst = rst;
  // Bindings to f802

  // f804
  logic [0:0] f804_wen;
  logic [31:0] f804_wdata;
  logic [0:0] f804_clk;
  logic [0:0] f804_rst;
  logic [31:0] f804_rdata;
  sr_buffer_32_1 f804(.wen(f804_wen), .wdata(f804_wdata), .clk(f804_clk), .rst(f804_rst), .rdata(f804_rdata));
  assign f804_clk = clk;
  assign f804_rst = rst;
  // Bindings to f804

  // f800
  logic [0:0] f800_wen;
  logic [31:0] f800_wdata;
  logic [0:0] f800_clk;
  logic [0:0] f800_rst;
  logic [31:0] f800_rdata;
  sr_buffer_32_1 f800(.wen(f800_wen), .wdata(f800_wdata), .clk(f800_clk), .rst(f800_rst), .rdata(f800_rdata));
  assign f800_clk = clk;
  assign f800_rst = rst;
  // Bindings to f800

  // f798
  logic [0:0] f798_wen;
  logic [31:0] f798_wdata;
  logic [0:0] f798_clk;
  logic [0:0] f798_rst;
  logic [31:0] f798_rdata;
  sr_buffer_32_1 f798(.wen(f798_wen), .wdata(f798_wdata), .clk(f798_clk), .rst(f798_rst), .rdata(f798_rdata));
  assign f798_clk = clk;
  assign f798_rst = rst;
  // Bindings to f798

  // f754
  logic [0:0] f754_wen;
  logic [31:0] f754_wdata;
  logic [0:0] f754_clk;
  logic [0:0] f754_rst;
  logic [31:0] f754_rdata;
  sr_buffer_32_1 f754(.wen(f754_wen), .wdata(f754_wdata), .clk(f754_clk), .rst(f754_rst), .rdata(f754_rdata));
  assign f754_clk = clk;
  assign f754_rst = rst;
  // Bindings to f754

  // f792
  logic [0:0] f792_wen;
  logic [31:0] f792_wdata;
  logic [0:0] f792_clk;
  logic [0:0] f792_rst;
  logic [31:0] f792_rdata;
  sr_buffer_32_1 f792(.wen(f792_wen), .wdata(f792_wdata), .clk(f792_clk), .rst(f792_rst), .rdata(f792_rdata));
  assign f792_clk = clk;
  assign f792_rst = rst;
  // Bindings to f792

  // f794
  logic [0:0] f794_wen;
  logic [31:0] f794_wdata;
  logic [0:0] f794_clk;
  logic [0:0] f794_rst;
  logic [31:0] f794_rdata;
  sr_buffer_32_1 f794(.wen(f794_wen), .wdata(f794_wdata), .clk(f794_clk), .rst(f794_rst), .rdata(f794_rdata));
  assign f794_clk = clk;
  assign f794_rst = rst;
  // Bindings to f794

  // f836
  logic [0:0] f836_wen;
  logic [31:0] f836_wdata;
  logic [0:0] f836_clk;
  logic [0:0] f836_rst;
  logic [31:0] f836_rdata;
  sr_buffer_32_1 f836(.wen(f836_wen), .wdata(f836_wdata), .clk(f836_clk), .rst(f836_rst), .rdata(f836_rdata));
  assign f836_clk = clk;
  assign f836_rst = rst;
  // Bindings to f836

  // f834
  logic [0:0] f834_wen;
  logic [31:0] f834_wdata;
  logic [0:0] f834_clk;
  logic [0:0] f834_rst;
  logic [31:0] f834_rdata;
  sr_buffer_32_1 f834(.wen(f834_wen), .wdata(f834_wdata), .clk(f834_clk), .rst(f834_rst), .rdata(f834_rdata));
  assign f834_clk = clk;
  assign f834_rst = rst;
  // Bindings to f834

  // f832
  logic [0:0] f832_wen;
  logic [31:0] f832_wdata;
  logic [0:0] f832_clk;
  logic [0:0] f832_rst;
  logic [31:0] f832_rdata;
  sr_buffer_32_1 f832(.wen(f832_wen), .wdata(f832_wdata), .clk(f832_clk), .rst(f832_rst), .rdata(f832_rdata));
  assign f832_clk = clk;
  assign f832_rst = rst;
  // Bindings to f832

  // f872
  logic [0:0] f872_wen;
  logic [31:0] f872_wdata;
  logic [0:0] f872_clk;
  logic [0:0] f872_rst;
  logic [31:0] f872_rdata;
  sr_buffer_32_1 f872(.wen(f872_wen), .wdata(f872_wdata), .clk(f872_clk), .rst(f872_rst), .rdata(f872_rdata));
  assign f872_clk = clk;
  assign f872_rst = rst;
  // Bindings to f872

  // f866
  logic [0:0] f866_wen;
  logic [31:0] f866_wdata;
  logic [0:0] f866_clk;
  logic [0:0] f866_rst;
  logic [31:0] f866_rdata;
  sr_buffer_32_1 f866(.wen(f866_wen), .wdata(f866_wdata), .clk(f866_clk), .rst(f866_rst), .rdata(f866_rdata));
  assign f866_clk = clk;
  assign f866_rst = rst;
  // Bindings to f866

  // f814
  logic [0:0] f814_wen;
  logic [31:0] f814_wdata;
  logic [0:0] f814_clk;
  logic [0:0] f814_rst;
  logic [31:0] f814_rdata;
  sr_buffer_32_1 f814(.wen(f814_wen), .wdata(f814_wdata), .clk(f814_clk), .rst(f814_rst), .rdata(f814_rdata));
  assign f814_clk = clk;
  assign f814_rst = rst;
  // Bindings to f814

  // f810
  logic [0:0] f810_wen;
  logic [31:0] f810_wdata;
  logic [0:0] f810_clk;
  logic [0:0] f810_rst;
  logic [31:0] f810_rdata;
  sr_buffer_32_1 f810(.wen(f810_wen), .wdata(f810_wdata), .clk(f810_clk), .rst(f810_rst), .rdata(f810_rdata));
  assign f810_clk = clk;
  assign f810_rst = rst;
  // Bindings to f810

  // f812
  logic [0:0] f812_wen;
  logic [31:0] f812_wdata;
  logic [0:0] f812_clk;
  logic [0:0] f812_rst;
  logic [31:0] f812_rdata;
  sr_buffer_32_1 f812(.wen(f812_wen), .wdata(f812_wdata), .clk(f812_clk), .rst(f812_rst), .rdata(f812_rdata));
  assign f812_clk = clk;
  assign f812_rst = rst;
  // Bindings to f812

  // f806
  logic [0:0] f806_wen;
  logic [31:0] f806_wdata;
  logic [0:0] f806_clk;
  logic [0:0] f806_rst;
  logic [31:0] f806_rdata;
  sr_buffer_32_1 f806(.wen(f806_wen), .wdata(f806_wdata), .clk(f806_clk), .rst(f806_rst), .rdata(f806_rdata));
  assign f806_clk = clk;
  assign f806_rst = rst;
  // Bindings to f806

  // f746
  logic [0:0] f746_wen;
  logic [31:0] f746_wdata;
  logic [0:0] f746_clk;
  logic [0:0] f746_rst;
  logic [31:0] f746_rdata;
  sr_buffer_32_1 f746(.wen(f746_wen), .wdata(f746_wdata), .clk(f746_clk), .rst(f746_rst), .rdata(f746_rdata));
  assign f746_clk = clk;
  assign f746_rst = rst;
  // Bindings to f746

  // f742
  logic [0:0] f742_wen;
  logic [31:0] f742_wdata;
  logic [0:0] f742_clk;
  logic [0:0] f742_rst;
  logic [31:0] f742_rdata;
  sr_buffer_32_1 f742(.wen(f742_wen), .wdata(f742_wdata), .clk(f742_clk), .rst(f742_rst), .rdata(f742_rdata));
  assign f742_clk = clk;
  assign f742_rst = rst;
  // Bindings to f742

  // f740
  logic [0:0] f740_wen;
  logic [31:0] f740_wdata;
  logic [0:0] f740_clk;
  logic [0:0] f740_rst;
  logic [31:0] f740_rdata;
  sr_buffer_32_1 f740(.wen(f740_wen), .wdata(f740_wdata), .clk(f740_clk), .rst(f740_rst), .rdata(f740_rdata));
  assign f740_clk = clk;
  assign f740_rst = rst;
  // Bindings to f740

  // f734
  logic [0:0] f734_wen;
  logic [31:0] f734_wdata;
  logic [0:0] f734_clk;
  logic [0:0] f734_rst;
  logic [31:0] f734_rdata;
  sr_buffer_32_1 f734(.wen(f734_wen), .wdata(f734_wdata), .clk(f734_clk), .rst(f734_rst), .rdata(f734_rdata));
  assign f734_clk = clk;
  assign f734_rst = rst;
  // Bindings to f734

  // f738
  logic [0:0] f738_wen;
  logic [31:0] f738_wdata;
  logic [0:0] f738_clk;
  logic [0:0] f738_rst;
  logic [31:0] f738_rdata;
  sr_buffer_32_1 f738(.wen(f738_wen), .wdata(f738_wdata), .clk(f738_clk), .rst(f738_rst), .rdata(f738_rdata));
  assign f738_clk = clk;
  assign f738_rst = rst;
  // Bindings to f738

  // f736
  logic [0:0] f736_wen;
  logic [31:0] f736_wdata;
  logic [0:0] f736_clk;
  logic [0:0] f736_rst;
  logic [31:0] f736_rdata;
  sr_buffer_32_1 f736(.wen(f736_wen), .wdata(f736_wdata), .clk(f736_clk), .rst(f736_rst), .rdata(f736_rdata));
  assign f736_clk = clk;
  assign f736_rst = rst;
  // Bindings to f736

  // f732
  logic [0:0] f732_wen;
  logic [31:0] f732_wdata;
  logic [0:0] f732_clk;
  logic [0:0] f732_rst;
  logic [31:0] f732_rdata;
  sr_buffer_32_1 f732(.wen(f732_wen), .wdata(f732_wdata), .clk(f732_clk), .rst(f732_rst), .rdata(f732_rdata));
  assign f732_clk = clk;
  assign f732_rst = rst;
  // Bindings to f732

  // f730
  logic [0:0] f730_wen;
  logic [31:0] f730_wdata;
  logic [0:0] f730_clk;
  logic [0:0] f730_rst;
  logic [31:0] f730_rdata;
  sr_buffer_32_1 f730(.wen(f730_wen), .wdata(f730_wdata), .clk(f730_clk), .rst(f730_rst), .rdata(f730_rdata));
  assign f730_clk = clk;
  assign f730_rst = rst;
  // Bindings to f730

  // f728
  logic [0:0] f728_wen;
  logic [31:0] f728_wdata;
  logic [0:0] f728_clk;
  logic [0:0] f728_rst;
  logic [31:0] f728_rdata;
  sr_buffer_32_1 f728(.wen(f728_wen), .wdata(f728_wdata), .clk(f728_clk), .rst(f728_rst), .rdata(f728_rdata));
  assign f728_clk = clk;
  assign f728_rst = rst;
  // Bindings to f728

  // f722
  logic [0:0] f722_wen;
  logic [31:0] f722_wdata;
  logic [0:0] f722_clk;
  logic [0:0] f722_rst;
  logic [31:0] f722_rdata;
  sr_buffer_32_1 f722(.wen(f722_wen), .wdata(f722_wdata), .clk(f722_clk), .rst(f722_rst), .rdata(f722_rdata));
  assign f722_clk = clk;
  assign f722_rst = rst;
  // Bindings to f722

  // f726
  logic [0:0] f726_wen;
  logic [31:0] f726_wdata;
  logic [0:0] f726_clk;
  logic [0:0] f726_rst;
  logic [31:0] f726_rdata;
  sr_buffer_32_1 f726(.wen(f726_wen), .wdata(f726_wdata), .clk(f726_clk), .rst(f726_rst), .rdata(f726_rdata));
  assign f726_clk = clk;
  assign f726_rst = rst;
  // Bindings to f726

  // f724
  logic [0:0] f724_wen;
  logic [31:0] f724_wdata;
  logic [0:0] f724_clk;
  logic [0:0] f724_rst;
  logic [31:0] f724_rdata;
  sr_buffer_32_1 f724(.wen(f724_wen), .wdata(f724_wdata), .clk(f724_clk), .rst(f724_rst), .rdata(f724_rdata));
  assign f724_clk = clk;
  assign f724_rst = rst;
  // Bindings to f724

  // f720
  logic [0:0] f720_wen;
  logic [31:0] f720_wdata;
  logic [0:0] f720_clk;
  logic [0:0] f720_rst;
  logic [31:0] f720_rdata;
  sr_buffer_32_1 f720(.wen(f720_wen), .wdata(f720_wdata), .clk(f720_clk), .rst(f720_rst), .rdata(f720_rdata));
  assign f720_clk = clk;
  assign f720_rst = rst;
  // Bindings to f720

  // f712
  logic [0:0] f712_wen;
  logic [31:0] f712_wdata;
  logic [0:0] f712_clk;
  logic [0:0] f712_rst;
  logic [31:0] f712_rdata;
  sr_buffer_32_1 f712(.wen(f712_wen), .wdata(f712_wdata), .clk(f712_clk), .rst(f712_rst), .rdata(f712_rdata));
  assign f712_clk = clk;
  assign f712_rst = rst;
  // Bindings to f712

  // f718
  logic [0:0] f718_wen;
  logic [31:0] f718_wdata;
  logic [0:0] f718_clk;
  logic [0:0] f718_rst;
  logic [31:0] f718_rdata;
  sr_buffer_32_1 f718(.wen(f718_wen), .wdata(f718_wdata), .clk(f718_clk), .rst(f718_rst), .rdata(f718_rdata));
  assign f718_clk = clk;
  assign f718_rst = rst;
  // Bindings to f718

  // f716
  logic [0:0] f716_wen;
  logic [31:0] f716_wdata;
  logic [0:0] f716_clk;
  logic [0:0] f716_rst;
  logic [31:0] f716_rdata;
  sr_buffer_32_1 f716(.wen(f716_wen), .wdata(f716_wdata), .clk(f716_clk), .rst(f716_rst), .rdata(f716_rdata));
  assign f716_clk = clk;
  assign f716_rst = rst;
  // Bindings to f716

  // f714
  logic [0:0] f714_wen;
  logic [31:0] f714_wdata;
  logic [0:0] f714_clk;
  logic [0:0] f714_rst;
  logic [31:0] f714_rdata;
  sr_buffer_32_1 f714(.wen(f714_wen), .wdata(f714_wdata), .clk(f714_clk), .rst(f714_rst), .rdata(f714_rdata));
  assign f714_clk = clk;
  assign f714_rst = rst;
  // Bindings to f714

  // f710
  logic [0:0] f710_wen;
  logic [31:0] f710_wdata;
  logic [0:0] f710_clk;
  logic [0:0] f710_rst;
  logic [31:0] f710_rdata;
  sr_buffer_32_1 f710(.wen(f710_wen), .wdata(f710_wdata), .clk(f710_clk), .rst(f710_rst), .rdata(f710_rdata));
  assign f710_clk = clk;
  assign f710_rst = rst;
  // Bindings to f710

  // f704
  logic [0:0] f704_wen;
  logic [31:0] f704_wdata;
  logic [0:0] f704_clk;
  logic [0:0] f704_rst;
  logic [31:0] f704_rdata;
  sr_buffer_32_1 f704(.wen(f704_wen), .wdata(f704_wdata), .clk(f704_clk), .rst(f704_rst), .rdata(f704_rdata));
  assign f704_clk = clk;
  assign f704_rst = rst;
  // Bindings to f704

  // f708
  logic [0:0] f708_wen;
  logic [31:0] f708_wdata;
  logic [0:0] f708_clk;
  logic [0:0] f708_rst;
  logic [31:0] f708_rdata;
  sr_buffer_32_1 f708(.wen(f708_wen), .wdata(f708_wdata), .clk(f708_clk), .rst(f708_rst), .rdata(f708_rdata));
  assign f708_clk = clk;
  assign f708_rst = rst;
  // Bindings to f708

  // f706
  logic [0:0] f706_wen;
  logic [31:0] f706_wdata;
  logic [0:0] f706_clk;
  logic [0:0] f706_rst;
  logic [31:0] f706_rdata;
  sr_buffer_32_1 f706(.wen(f706_wen), .wdata(f706_wdata), .clk(f706_clk), .rst(f706_rst), .rdata(f706_rdata));
  assign f706_clk = clk;
  assign f706_rst = rst;
  // Bindings to f706

  // f1226
  logic [0:0] f1226_wen;
  logic [31:0] f1226_wdata;
  logic [0:0] f1226_clk;
  logic [0:0] f1226_rst;
  logic [31:0] f1226_rdata;
  sr_buffer_32_1 f1226(.wen(f1226_wen), .wdata(f1226_wdata), .clk(f1226_clk), .rst(f1226_rst), .rdata(f1226_rdata));
  assign f1226_clk = clk;
  assign f1226_rst = rst;
  // Bindings to f1226

  // f1248
  logic [0:0] f1248_wen;
  logic [31:0] f1248_wdata;
  logic [0:0] f1248_clk;
  logic [0:0] f1248_rst;
  logic [31:0] f1248_rdata;
  sr_buffer_32_1 f1248(.wen(f1248_wen), .wdata(f1248_wdata), .clk(f1248_clk), .rst(f1248_rst), .rdata(f1248_rdata));
  assign f1248_clk = clk;
  assign f1248_rst = rst;
  // Bindings to f1248

  // f1252
  logic [0:0] f1252_wen;
  logic [31:0] f1252_wdata;
  logic [0:0] f1252_clk;
  logic [0:0] f1252_rst;
  logic [31:0] f1252_rdata;
  sr_buffer_32_1 f1252(.wen(f1252_wen), .wdata(f1252_wdata), .clk(f1252_clk), .rst(f1252_rst), .rdata(f1252_rdata));
  assign f1252_clk = clk;
  assign f1252_rst = rst;
  // Bindings to f1252

  // f1250
  logic [0:0] f1250_wen;
  logic [31:0] f1250_wdata;
  logic [0:0] f1250_clk;
  logic [0:0] f1250_rst;
  logic [31:0] f1250_rdata;
  sr_buffer_32_1 f1250(.wen(f1250_wen), .wdata(f1250_wdata), .clk(f1250_clk), .rst(f1250_rst), .rdata(f1250_rdata));
  assign f1250_clk = clk;
  assign f1250_rst = rst;
  // Bindings to f1250

  // f1228
  logic [0:0] f1228_wen;
  logic [31:0] f1228_wdata;
  logic [0:0] f1228_clk;
  logic [0:0] f1228_rst;
  logic [31:0] f1228_rdata;
  sr_buffer_32_1 f1228(.wen(f1228_wen), .wdata(f1228_wdata), .clk(f1228_clk), .rst(f1228_rst), .rdata(f1228_rdata));
  assign f1228_clk = clk;
  assign f1228_rst = rst;
  // Bindings to f1228

  // f1246
  logic [0:0] f1246_wen;
  logic [31:0] f1246_wdata;
  logic [0:0] f1246_clk;
  logic [0:0] f1246_rst;
  logic [31:0] f1246_rdata;
  sr_buffer_32_1 f1246(.wen(f1246_wen), .wdata(f1246_wdata), .clk(f1246_clk), .rst(f1246_rst), .rdata(f1246_rdata));
  assign f1246_clk = clk;
  assign f1246_rst = rst;
  // Bindings to f1246

  // f1242
  logic [0:0] f1242_wen;
  logic [31:0] f1242_wdata;
  logic [0:0] f1242_clk;
  logic [0:0] f1242_rst;
  logic [31:0] f1242_rdata;
  sr_buffer_32_1 f1242(.wen(f1242_wen), .wdata(f1242_wdata), .clk(f1242_clk), .rst(f1242_rst), .rdata(f1242_rdata));
  assign f1242_clk = clk;
  assign f1242_rst = rst;
  // Bindings to f1242

  // f1244
  logic [0:0] f1244_wen;
  logic [31:0] f1244_wdata;
  logic [0:0] f1244_clk;
  logic [0:0] f1244_rst;
  logic [31:0] f1244_rdata;
  sr_buffer_32_1 f1244(.wen(f1244_wen), .wdata(f1244_wdata), .clk(f1244_clk), .rst(f1244_rst), .rdata(f1244_rdata));
  assign f1244_clk = clk;
  assign f1244_rst = rst;
  // Bindings to f1244

  // f1240
  logic [0:0] f1240_wen;
  logic [31:0] f1240_wdata;
  logic [0:0] f1240_clk;
  logic [0:0] f1240_rst;
  logic [31:0] f1240_rdata;
  sr_buffer_32_1 f1240(.wen(f1240_wen), .wdata(f1240_wdata), .clk(f1240_clk), .rst(f1240_rst), .rdata(f1240_rdata));
  assign f1240_clk = clk;
  assign f1240_rst = rst;
  // Bindings to f1240

  // f1238
  logic [0:0] f1238_wen;
  logic [31:0] f1238_wdata;
  logic [0:0] f1238_clk;
  logic [0:0] f1238_rst;
  logic [31:0] f1238_rdata;
  sr_buffer_32_1 f1238(.wen(f1238_wen), .wdata(f1238_wdata), .clk(f1238_clk), .rst(f1238_rst), .rdata(f1238_rdata));
  assign f1238_clk = clk;
  assign f1238_rst = rst;
  // Bindings to f1238

  // f1236
  logic [0:0] f1236_wen;
  logic [31:0] f1236_wdata;
  logic [0:0] f1236_clk;
  logic [0:0] f1236_rst;
  logic [31:0] f1236_rdata;
  sr_buffer_32_1 f1236(.wen(f1236_wen), .wdata(f1236_wdata), .clk(f1236_clk), .rst(f1236_rst), .rdata(f1236_rdata));
  assign f1236_clk = clk;
  assign f1236_rst = rst;
  // Bindings to f1236

  // f1234
  logic [0:0] f1234_wen;
  logic [31:0] f1234_wdata;
  logic [0:0] f1234_clk;
  logic [0:0] f1234_rst;
  logic [31:0] f1234_rdata;
  sr_buffer_32_1 f1234(.wen(f1234_wen), .wdata(f1234_wdata), .clk(f1234_clk), .rst(f1234_rst), .rdata(f1234_rdata));
  assign f1234_clk = clk;
  assign f1234_rst = rst;
  // Bindings to f1234

  // f1230
  logic [0:0] f1230_wen;
  logic [31:0] f1230_wdata;
  logic [0:0] f1230_clk;
  logic [0:0] f1230_rst;
  logic [31:0] f1230_rdata;
  sr_buffer_32_1 f1230(.wen(f1230_wen), .wdata(f1230_wdata), .clk(f1230_clk), .rst(f1230_rst), .rdata(f1230_rdata));
  assign f1230_clk = clk;
  assign f1230_rst = rst;
  // Bindings to f1230

  // f1232
  logic [0:0] f1232_wen;
  logic [31:0] f1232_wdata;
  logic [0:0] f1232_clk;
  logic [0:0] f1232_rst;
  logic [31:0] f1232_rdata;
  sr_buffer_32_1 f1232(.wen(f1232_wen), .wdata(f1232_wdata), .clk(f1232_clk), .rst(f1232_rst), .rdata(f1232_rdata));
  assign f1232_clk = clk;
  assign f1232_rst = rst;
  // Bindings to f1232

  // f1224
  logic [0:0] f1224_wen;
  logic [31:0] f1224_wdata;
  logic [0:0] f1224_clk;
  logic [0:0] f1224_rst;
  logic [31:0] f1224_rdata;
  sr_buffer_32_1 f1224(.wen(f1224_wen), .wdata(f1224_wdata), .clk(f1224_clk), .rst(f1224_rst), .rdata(f1224_rdata));
  assign f1224_clk = clk;
  assign f1224_rst = rst;
  // Bindings to f1224

  // f1222
  logic [0:0] f1222_wen;
  logic [31:0] f1222_wdata;
  logic [0:0] f1222_clk;
  logic [0:0] f1222_rst;
  logic [31:0] f1222_rdata;
  sr_buffer_32_1 f1222(.wen(f1222_wen), .wdata(f1222_wdata), .clk(f1222_clk), .rst(f1222_rst), .rdata(f1222_rdata));
  assign f1222_clk = clk;
  assign f1222_rst = rst;
  // Bindings to f1222

  // f1220
  logic [0:0] f1220_wen;
  logic [31:0] f1220_wdata;
  logic [0:0] f1220_clk;
  logic [0:0] f1220_rst;
  logic [31:0] f1220_rdata;
  sr_buffer_32_1 f1220(.wen(f1220_wen), .wdata(f1220_wdata), .clk(f1220_clk), .rst(f1220_rst), .rdata(f1220_rdata));
  assign f1220_clk = clk;
  assign f1220_rst = rst;
  // Bindings to f1220

  // f1218
  logic [0:0] f1218_wen;
  logic [31:0] f1218_wdata;
  logic [0:0] f1218_clk;
  logic [0:0] f1218_rst;
  logic [31:0] f1218_rdata;
  sr_buffer_32_1 f1218(.wen(f1218_wen), .wdata(f1218_wdata), .clk(f1218_clk), .rst(f1218_rst), .rdata(f1218_rdata));
  assign f1218_clk = clk;
  assign f1218_rst = rst;
  // Bindings to f1218

  // f1204
  logic [0:0] f1204_wen;
  logic [31:0] f1204_wdata;
  logic [0:0] f1204_clk;
  logic [0:0] f1204_rst;
  logic [31:0] f1204_rdata;
  sr_buffer_32_1 f1204(.wen(f1204_wen), .wdata(f1204_wdata), .clk(f1204_clk), .rst(f1204_rst), .rdata(f1204_rdata));
  assign f1204_clk = clk;
  assign f1204_rst = rst;
  // Bindings to f1204

  // f1216
  logic [0:0] f1216_wen;
  logic [31:0] f1216_wdata;
  logic [0:0] f1216_clk;
  logic [0:0] f1216_rst;
  logic [31:0] f1216_rdata;
  sr_buffer_32_1 f1216(.wen(f1216_wen), .wdata(f1216_wdata), .clk(f1216_clk), .rst(f1216_rst), .rdata(f1216_rdata));
  assign f1216_clk = clk;
  assign f1216_rst = rst;
  // Bindings to f1216

  // f1214
  logic [0:0] f1214_wen;
  logic [31:0] f1214_wdata;
  logic [0:0] f1214_clk;
  logic [0:0] f1214_rst;
  logic [31:0] f1214_rdata;
  sr_buffer_32_1 f1214(.wen(f1214_wen), .wdata(f1214_wdata), .clk(f1214_clk), .rst(f1214_rst), .rdata(f1214_rdata));
  assign f1214_clk = clk;
  assign f1214_rst = rst;
  // Bindings to f1214

  // f1212
  logic [0:0] f1212_wen;
  logic [31:0] f1212_wdata;
  logic [0:0] f1212_clk;
  logic [0:0] f1212_rst;
  logic [31:0] f1212_rdata;
  sr_buffer_32_1 f1212(.wen(f1212_wen), .wdata(f1212_wdata), .clk(f1212_clk), .rst(f1212_rst), .rdata(f1212_rdata));
  assign f1212_clk = clk;
  assign f1212_rst = rst;
  // Bindings to f1212

  // f1210
  logic [0:0] f1210_wen;
  logic [31:0] f1210_wdata;
  logic [0:0] f1210_clk;
  logic [0:0] f1210_rst;
  logic [31:0] f1210_rdata;
  sr_buffer_32_1 f1210(.wen(f1210_wen), .wdata(f1210_wdata), .clk(f1210_clk), .rst(f1210_rst), .rdata(f1210_rdata));
  assign f1210_clk = clk;
  assign f1210_rst = rst;
  // Bindings to f1210

  // f1208
  logic [0:0] f1208_wen;
  logic [31:0] f1208_wdata;
  logic [0:0] f1208_clk;
  logic [0:0] f1208_rst;
  logic [31:0] f1208_rdata;
  sr_buffer_32_1 f1208(.wen(f1208_wen), .wdata(f1208_wdata), .clk(f1208_clk), .rst(f1208_rst), .rdata(f1208_rdata));
  assign f1208_clk = clk;
  assign f1208_rst = rst;
  // Bindings to f1208

  // f1206
  logic [0:0] f1206_wen;
  logic [31:0] f1206_wdata;
  logic [0:0] f1206_clk;
  logic [0:0] f1206_rst;
  logic [31:0] f1206_rdata;
  sr_buffer_32_1 f1206(.wen(f1206_wen), .wdata(f1206_wdata), .clk(f1206_clk), .rst(f1206_rst), .rdata(f1206_rdata));
  assign f1206_clk = clk;
  assign f1206_rst = rst;
  // Bindings to f1206

  // f1202
  logic [0:0] f1202_wen;
  logic [31:0] f1202_wdata;
  logic [0:0] f1202_clk;
  logic [0:0] f1202_rst;
  logic [31:0] f1202_rdata;
  sr_buffer_32_1 f1202(.wen(f1202_wen), .wdata(f1202_wdata), .clk(f1202_clk), .rst(f1202_rst), .rdata(f1202_rdata));
  assign f1202_clk = clk;
  assign f1202_rst = rst;
  // Bindings to f1202

  // f1200
  logic [0:0] f1200_wen;
  logic [31:0] f1200_wdata;
  logic [0:0] f1200_clk;
  logic [0:0] f1200_rst;
  logic [31:0] f1200_rdata;
  sr_buffer_32_1 f1200(.wen(f1200_wen), .wdata(f1200_wdata), .clk(f1200_clk), .rst(f1200_rst), .rdata(f1200_rdata));
  assign f1200_clk = clk;
  assign f1200_rst = rst;
  // Bindings to f1200

  // f1198
  logic [0:0] f1198_wen;
  logic [31:0] f1198_wdata;
  logic [0:0] f1198_clk;
  logic [0:0] f1198_rst;
  logic [31:0] f1198_rdata;
  sr_buffer_32_1 f1198(.wen(f1198_wen), .wdata(f1198_wdata), .clk(f1198_clk), .rst(f1198_rst), .rdata(f1198_rdata));
  assign f1198_clk = clk;
  assign f1198_rst = rst;
  // Bindings to f1198

  // f1194
  logic [0:0] f1194_wen;
  logic [31:0] f1194_wdata;
  logic [0:0] f1194_clk;
  logic [0:0] f1194_rst;
  logic [31:0] f1194_rdata;
  sr_buffer_32_1 f1194(.wen(f1194_wen), .wdata(f1194_wdata), .clk(f1194_clk), .rst(f1194_rst), .rdata(f1194_rdata));
  assign f1194_clk = clk;
  assign f1194_rst = rst;
  // Bindings to f1194

  // f1196
  logic [0:0] f1196_wen;
  logic [31:0] f1196_wdata;
  logic [0:0] f1196_clk;
  logic [0:0] f1196_rst;
  logic [31:0] f1196_rdata;
  sr_buffer_32_1 f1196(.wen(f1196_wen), .wdata(f1196_wdata), .clk(f1196_clk), .rst(f1196_rst), .rdata(f1196_rdata));
  assign f1196_clk = clk;
  assign f1196_rst = rst;
  // Bindings to f1196

  // f1192
  logic [0:0] f1192_wen;
  logic [31:0] f1192_wdata;
  logic [0:0] f1192_clk;
  logic [0:0] f1192_rst;
  logic [31:0] f1192_rdata;
  sr_buffer_32_1 f1192(.wen(f1192_wen), .wdata(f1192_wdata), .clk(f1192_clk), .rst(f1192_rst), .rdata(f1192_rdata));
  assign f1192_clk = clk;
  assign f1192_rst = rst;
  // Bindings to f1192

  // f1190
  logic [0:0] f1190_wen;
  logic [31:0] f1190_wdata;
  logic [0:0] f1190_clk;
  logic [0:0] f1190_rst;
  logic [31:0] f1190_rdata;
  sr_buffer_32_1 f1190(.wen(f1190_wen), .wdata(f1190_wdata), .clk(f1190_clk), .rst(f1190_rst), .rdata(f1190_rdata));
  assign f1190_clk = clk;
  assign f1190_rst = rst;
  // Bindings to f1190

  // f1180
  logic [0:0] f1180_wen;
  logic [31:0] f1180_wdata;
  logic [0:0] f1180_clk;
  logic [0:0] f1180_rst;
  logic [31:0] f1180_rdata;
  sr_buffer_32_1 f1180(.wen(f1180_wen), .wdata(f1180_wdata), .clk(f1180_clk), .rst(f1180_rst), .rdata(f1180_rdata));
  assign f1180_clk = clk;
  assign f1180_rst = rst;
  // Bindings to f1180

  // f1188
  logic [0:0] f1188_wen;
  logic [31:0] f1188_wdata;
  logic [0:0] f1188_clk;
  logic [0:0] f1188_rst;
  logic [31:0] f1188_rdata;
  sr_buffer_32_1 f1188(.wen(f1188_wen), .wdata(f1188_wdata), .clk(f1188_clk), .rst(f1188_rst), .rdata(f1188_rdata));
  assign f1188_clk = clk;
  assign f1188_rst = rst;
  // Bindings to f1188

  // f1186
  logic [0:0] f1186_wen;
  logic [31:0] f1186_wdata;
  logic [0:0] f1186_clk;
  logic [0:0] f1186_rst;
  logic [31:0] f1186_rdata;
  sr_buffer_32_1 f1186(.wen(f1186_wen), .wdata(f1186_wdata), .clk(f1186_clk), .rst(f1186_rst), .rdata(f1186_rdata));
  assign f1186_clk = clk;
  assign f1186_rst = rst;
  // Bindings to f1186

  // f1182
  logic [0:0] f1182_wen;
  logic [31:0] f1182_wdata;
  logic [0:0] f1182_clk;
  logic [0:0] f1182_rst;
  logic [31:0] f1182_rdata;
  sr_buffer_32_1 f1182(.wen(f1182_wen), .wdata(f1182_wdata), .clk(f1182_clk), .rst(f1182_rst), .rdata(f1182_rdata));
  assign f1182_clk = clk;
  assign f1182_rst = rst;
  // Bindings to f1182

  // f1184
  logic [0:0] f1184_wen;
  logic [31:0] f1184_wdata;
  logic [0:0] f1184_clk;
  logic [0:0] f1184_rst;
  logic [31:0] f1184_rdata;
  sr_buffer_32_1 f1184(.wen(f1184_wen), .wdata(f1184_wdata), .clk(f1184_clk), .rst(f1184_rst), .rdata(f1184_rdata));
  assign f1184_clk = clk;
  assign f1184_rst = rst;
  // Bindings to f1184

  // f1178
  logic [0:0] f1178_wen;
  logic [31:0] f1178_wdata;
  logic [0:0] f1178_clk;
  logic [0:0] f1178_rst;
  logic [31:0] f1178_rdata;
  sr_buffer_32_1 f1178(.wen(f1178_wen), .wdata(f1178_wdata), .clk(f1178_clk), .rst(f1178_rst), .rdata(f1178_rdata));
  assign f1178_clk = clk;
  assign f1178_rst = rst;
  // Bindings to f1178

  // f1176
  logic [0:0] f1176_wen;
  logic [31:0] f1176_wdata;
  logic [0:0] f1176_clk;
  logic [0:0] f1176_rst;
  logic [31:0] f1176_rdata;
  sr_buffer_32_1 f1176(.wen(f1176_wen), .wdata(f1176_wdata), .clk(f1176_clk), .rst(f1176_rst), .rdata(f1176_rdata));
  assign f1176_clk = clk;
  assign f1176_rst = rst;
  // Bindings to f1176

  // f1174
  logic [0:0] f1174_wen;
  logic [31:0] f1174_wdata;
  logic [0:0] f1174_clk;
  logic [0:0] f1174_rst;
  logic [31:0] f1174_rdata;
  sr_buffer_32_1 f1174(.wen(f1174_wen), .wdata(f1174_wdata), .clk(f1174_clk), .rst(f1174_rst), .rdata(f1174_rdata));
  assign f1174_clk = clk;
  assign f1174_rst = rst;
  // Bindings to f1174

  // f1172
  logic [0:0] f1172_wen;
  logic [31:0] f1172_wdata;
  logic [0:0] f1172_clk;
  logic [0:0] f1172_rst;
  logic [31:0] f1172_rdata;
  sr_buffer_32_1 f1172(.wen(f1172_wen), .wdata(f1172_wdata), .clk(f1172_clk), .rst(f1172_rst), .rdata(f1172_rdata));
  assign f1172_clk = clk;
  assign f1172_rst = rst;
  // Bindings to f1172

  // f1170
  logic [0:0] f1170_wen;
  logic [31:0] f1170_wdata;
  logic [0:0] f1170_clk;
  logic [0:0] f1170_rst;
  logic [31:0] f1170_rdata;
  sr_buffer_32_1 f1170(.wen(f1170_wen), .wdata(f1170_wdata), .clk(f1170_clk), .rst(f1170_rst), .rdata(f1170_rdata));
  assign f1170_clk = clk;
  assign f1170_rst = rst;
  // Bindings to f1170

  // f1168
  logic [0:0] f1168_wen;
  logic [31:0] f1168_wdata;
  logic [0:0] f1168_clk;
  logic [0:0] f1168_rst;
  logic [31:0] f1168_rdata;
  sr_buffer_32_1 f1168(.wen(f1168_wen), .wdata(f1168_wdata), .clk(f1168_clk), .rst(f1168_rst), .rdata(f1168_rdata));
  assign f1168_clk = clk;
  assign f1168_rst = rst;
  // Bindings to f1168

  // f1166
  logic [0:0] f1166_wen;
  logic [31:0] f1166_wdata;
  logic [0:0] f1166_clk;
  logic [0:0] f1166_rst;
  logic [31:0] f1166_rdata;
  sr_buffer_32_1 f1166(.wen(f1166_wen), .wdata(f1166_wdata), .clk(f1166_clk), .rst(f1166_rst), .rdata(f1166_rdata));
  assign f1166_clk = clk;
  assign f1166_rst = rst;
  // Bindings to f1166

  // f1164
  logic [0:0] f1164_wen;
  logic [31:0] f1164_wdata;
  logic [0:0] f1164_clk;
  logic [0:0] f1164_rst;
  logic [31:0] f1164_rdata;
  sr_buffer_32_1 f1164(.wen(f1164_wen), .wdata(f1164_wdata), .clk(f1164_clk), .rst(f1164_rst), .rdata(f1164_rdata));
  assign f1164_clk = clk;
  assign f1164_rst = rst;
  // Bindings to f1164

  // f1162
  logic [0:0] f1162_wen;
  logic [31:0] f1162_wdata;
  logic [0:0] f1162_clk;
  logic [0:0] f1162_rst;
  logic [31:0] f1162_rdata;
  sr_buffer_32_1 f1162(.wen(f1162_wen), .wdata(f1162_wdata), .clk(f1162_clk), .rst(f1162_rst), .rdata(f1162_rdata));
  assign f1162_clk = clk;
  assign f1162_rst = rst;
  // Bindings to f1162

  // f1154
  logic [0:0] f1154_wen;
  logic [31:0] f1154_wdata;
  logic [0:0] f1154_clk;
  logic [0:0] f1154_rst;
  logic [31:0] f1154_rdata;
  sr_buffer_32_1 f1154(.wen(f1154_wen), .wdata(f1154_wdata), .clk(f1154_clk), .rst(f1154_rst), .rdata(f1154_rdata));
  assign f1154_clk = clk;
  assign f1154_rst = rst;
  // Bindings to f1154

  // f1160
  logic [0:0] f1160_wen;
  logic [31:0] f1160_wdata;
  logic [0:0] f1160_clk;
  logic [0:0] f1160_rst;
  logic [31:0] f1160_rdata;
  sr_buffer_32_1 f1160(.wen(f1160_wen), .wdata(f1160_wdata), .clk(f1160_clk), .rst(f1160_rst), .rdata(f1160_rdata));
  assign f1160_clk = clk;
  assign f1160_rst = rst;
  // Bindings to f1160

  // f1158
  logic [0:0] f1158_wen;
  logic [31:0] f1158_wdata;
  logic [0:0] f1158_clk;
  logic [0:0] f1158_rst;
  logic [31:0] f1158_rdata;
  sr_buffer_32_1 f1158(.wen(f1158_wen), .wdata(f1158_wdata), .clk(f1158_clk), .rst(f1158_rst), .rdata(f1158_rdata));
  assign f1158_clk = clk;
  assign f1158_rst = rst;
  // Bindings to f1158

  // f1156
  logic [0:0] f1156_wen;
  logic [31:0] f1156_wdata;
  logic [0:0] f1156_clk;
  logic [0:0] f1156_rst;
  logic [31:0] f1156_rdata;
  sr_buffer_32_1 f1156(.wen(f1156_wen), .wdata(f1156_wdata), .clk(f1156_clk), .rst(f1156_rst), .rdata(f1156_rdata));
  assign f1156_clk = clk;
  assign f1156_rst = rst;
  // Bindings to f1156

  // f1152
  logic [0:0] f1152_wen;
  logic [31:0] f1152_wdata;
  logic [0:0] f1152_clk;
  logic [0:0] f1152_rst;
  logic [31:0] f1152_rdata;
  sr_buffer_32_1 f1152(.wen(f1152_wen), .wdata(f1152_wdata), .clk(f1152_clk), .rst(f1152_rst), .rdata(f1152_rdata));
  assign f1152_clk = clk;
  assign f1152_rst = rst;
  // Bindings to f1152

  // f1150
  logic [0:0] f1150_wen;
  logic [31:0] f1150_wdata;
  logic [0:0] f1150_clk;
  logic [0:0] f1150_rst;
  logic [31:0] f1150_rdata;
  sr_buffer_32_1 f1150(.wen(f1150_wen), .wdata(f1150_wdata), .clk(f1150_clk), .rst(f1150_rst), .rdata(f1150_rdata));
  assign f1150_clk = clk;
  assign f1150_rst = rst;
  // Bindings to f1150

  // f1140
  logic [0:0] f1140_wen;
  logic [31:0] f1140_wdata;
  logic [0:0] f1140_clk;
  logic [0:0] f1140_rst;
  logic [31:0] f1140_rdata;
  sr_buffer_32_1 f1140(.wen(f1140_wen), .wdata(f1140_wdata), .clk(f1140_clk), .rst(f1140_rst), .rdata(f1140_rdata));
  assign f1140_clk = clk;
  assign f1140_rst = rst;
  // Bindings to f1140

  // f1148
  logic [0:0] f1148_wen;
  logic [31:0] f1148_wdata;
  logic [0:0] f1148_clk;
  logic [0:0] f1148_rst;
  logic [31:0] f1148_rdata;
  sr_buffer_32_1 f1148(.wen(f1148_wen), .wdata(f1148_wdata), .clk(f1148_clk), .rst(f1148_rst), .rdata(f1148_rdata));
  assign f1148_clk = clk;
  assign f1148_rst = rst;
  // Bindings to f1148

  // f1146
  logic [0:0] f1146_wen;
  logic [31:0] f1146_wdata;
  logic [0:0] f1146_clk;
  logic [0:0] f1146_rst;
  logic [31:0] f1146_rdata;
  sr_buffer_32_1 f1146(.wen(f1146_wen), .wdata(f1146_wdata), .clk(f1146_clk), .rst(f1146_rst), .rdata(f1146_rdata));
  assign f1146_clk = clk;
  assign f1146_rst = rst;
  // Bindings to f1146

  // f1142
  logic [0:0] f1142_wen;
  logic [31:0] f1142_wdata;
  logic [0:0] f1142_clk;
  logic [0:0] f1142_rst;
  logic [31:0] f1142_rdata;
  sr_buffer_32_1 f1142(.wen(f1142_wen), .wdata(f1142_wdata), .clk(f1142_clk), .rst(f1142_rst), .rdata(f1142_rdata));
  assign f1142_clk = clk;
  assign f1142_rst = rst;
  // Bindings to f1142

  // f1144
  logic [0:0] f1144_wen;
  logic [31:0] f1144_wdata;
  logic [0:0] f1144_clk;
  logic [0:0] f1144_rst;
  logic [31:0] f1144_rdata;
  sr_buffer_32_1 f1144(.wen(f1144_wen), .wdata(f1144_wdata), .clk(f1144_clk), .rst(f1144_rst), .rdata(f1144_rdata));
  assign f1144_clk = clk;
  assign f1144_rst = rst;
  // Bindings to f1144

  // f1136
  logic [0:0] f1136_wen;
  logic [31:0] f1136_wdata;
  logic [0:0] f1136_clk;
  logic [0:0] f1136_rst;
  logic [31:0] f1136_rdata;
  sr_buffer_32_1 f1136(.wen(f1136_wen), .wdata(f1136_wdata), .clk(f1136_clk), .rst(f1136_rst), .rdata(f1136_rdata));
  assign f1136_clk = clk;
  assign f1136_rst = rst;
  // Bindings to f1136

  // f1138
  logic [0:0] f1138_wen;
  logic [31:0] f1138_wdata;
  logic [0:0] f1138_clk;
  logic [0:0] f1138_rst;
  logic [31:0] f1138_rdata;
  sr_buffer_32_1 f1138(.wen(f1138_wen), .wdata(f1138_wdata), .clk(f1138_clk), .rst(f1138_rst), .rdata(f1138_rdata));
  assign f1138_clk = clk;
  assign f1138_rst = rst;
  // Bindings to f1138

  // f1120
  logic [0:0] f1120_wen;
  logic [31:0] f1120_wdata;
  logic [0:0] f1120_clk;
  logic [0:0] f1120_rst;
  logic [31:0] f1120_rdata;
  sr_buffer_32_1 f1120(.wen(f1120_wen), .wdata(f1120_wdata), .clk(f1120_clk), .rst(f1120_rst), .rdata(f1120_rdata));
  assign f1120_clk = clk;
  assign f1120_rst = rst;
  // Bindings to f1120

  // f1134
  logic [0:0] f1134_wen;
  logic [31:0] f1134_wdata;
  logic [0:0] f1134_clk;
  logic [0:0] f1134_rst;
  logic [31:0] f1134_rdata;
  sr_buffer_32_1 f1134(.wen(f1134_wen), .wdata(f1134_wdata), .clk(f1134_clk), .rst(f1134_rst), .rdata(f1134_rdata));
  assign f1134_clk = clk;
  assign f1134_rst = rst;
  // Bindings to f1134

  // f1132
  logic [0:0] f1132_wen;
  logic [31:0] f1132_wdata;
  logic [0:0] f1132_clk;
  logic [0:0] f1132_rst;
  logic [31:0] f1132_rdata;
  sr_buffer_32_1 f1132(.wen(f1132_wen), .wdata(f1132_wdata), .clk(f1132_clk), .rst(f1132_rst), .rdata(f1132_rdata));
  assign f1132_clk = clk;
  assign f1132_rst = rst;
  // Bindings to f1132

  // f1130
  logic [0:0] f1130_wen;
  logic [31:0] f1130_wdata;
  logic [0:0] f1130_clk;
  logic [0:0] f1130_rst;
  logic [31:0] f1130_rdata;
  sr_buffer_32_1 f1130(.wen(f1130_wen), .wdata(f1130_wdata), .clk(f1130_clk), .rst(f1130_rst), .rdata(f1130_rdata));
  assign f1130_clk = clk;
  assign f1130_rst = rst;
  // Bindings to f1130

  // f1128
  logic [0:0] f1128_wen;
  logic [31:0] f1128_wdata;
  logic [0:0] f1128_clk;
  logic [0:0] f1128_rst;
  logic [31:0] f1128_rdata;
  sr_buffer_32_1 f1128(.wen(f1128_wen), .wdata(f1128_wdata), .clk(f1128_clk), .rst(f1128_rst), .rdata(f1128_rdata));
  assign f1128_clk = clk;
  assign f1128_rst = rst;
  // Bindings to f1128

  // f1122
  logic [0:0] f1122_wen;
  logic [31:0] f1122_wdata;
  logic [0:0] f1122_clk;
  logic [0:0] f1122_rst;
  logic [31:0] f1122_rdata;
  sr_buffer_32_1 f1122(.wen(f1122_wen), .wdata(f1122_wdata), .clk(f1122_clk), .rst(f1122_rst), .rdata(f1122_rdata));
  assign f1122_clk = clk;
  assign f1122_rst = rst;
  // Bindings to f1122

  // f1126
  logic [0:0] f1126_wen;
  logic [31:0] f1126_wdata;
  logic [0:0] f1126_clk;
  logic [0:0] f1126_rst;
  logic [31:0] f1126_rdata;
  sr_buffer_32_1 f1126(.wen(f1126_wen), .wdata(f1126_wdata), .clk(f1126_clk), .rst(f1126_rst), .rdata(f1126_rdata));
  assign f1126_clk = clk;
  assign f1126_rst = rst;
  // Bindings to f1126

  // f1124
  logic [0:0] f1124_wen;
  logic [31:0] f1124_wdata;
  logic [0:0] f1124_clk;
  logic [0:0] f1124_rst;
  logic [31:0] f1124_rdata;
  sr_buffer_32_1 f1124(.wen(f1124_wen), .wdata(f1124_wdata), .clk(f1124_clk), .rst(f1124_rst), .rdata(f1124_rdata));
  assign f1124_clk = clk;
  assign f1124_rst = rst;
  // Bindings to f1124

  // f1118
  logic [0:0] f1118_wen;
  logic [31:0] f1118_wdata;
  logic [0:0] f1118_clk;
  logic [0:0] f1118_rst;
  logic [31:0] f1118_rdata;
  sr_buffer_32_1 f1118(.wen(f1118_wen), .wdata(f1118_wdata), .clk(f1118_clk), .rst(f1118_rst), .rdata(f1118_rdata));
  assign f1118_clk = clk;
  assign f1118_rst = rst;
  // Bindings to f1118

  // f1116
  logic [0:0] f1116_wen;
  logic [31:0] f1116_wdata;
  logic [0:0] f1116_clk;
  logic [0:0] f1116_rst;
  logic [31:0] f1116_rdata;
  sr_buffer_32_1 f1116(.wen(f1116_wen), .wdata(f1116_wdata), .clk(f1116_clk), .rst(f1116_rst), .rdata(f1116_rdata));
  assign f1116_clk = clk;
  assign f1116_rst = rst;
  // Bindings to f1116

  // f1114
  logic [0:0] f1114_wen;
  logic [31:0] f1114_wdata;
  logic [0:0] f1114_clk;
  logic [0:0] f1114_rst;
  logic [31:0] f1114_rdata;
  sr_buffer_32_1 f1114(.wen(f1114_wen), .wdata(f1114_wdata), .clk(f1114_clk), .rst(f1114_rst), .rdata(f1114_rdata));
  assign f1114_clk = clk;
  assign f1114_rst = rst;
  // Bindings to f1114

  // f1112
  logic [0:0] f1112_wen;
  logic [31:0] f1112_wdata;
  logic [0:0] f1112_clk;
  logic [0:0] f1112_rst;
  logic [31:0] f1112_rdata;
  sr_buffer_32_1 f1112(.wen(f1112_wen), .wdata(f1112_wdata), .clk(f1112_clk), .rst(f1112_rst), .rdata(f1112_rdata));
  assign f1112_clk = clk;
  assign f1112_rst = rst;
  // Bindings to f1112

  // f1110
  logic [0:0] f1110_wen;
  logic [31:0] f1110_wdata;
  logic [0:0] f1110_clk;
  logic [0:0] f1110_rst;
  logic [31:0] f1110_rdata;
  sr_buffer_32_1 f1110(.wen(f1110_wen), .wdata(f1110_wdata), .clk(f1110_clk), .rst(f1110_rst), .rdata(f1110_rdata));
  assign f1110_clk = clk;
  assign f1110_rst = rst;
  // Bindings to f1110

  // f1108
  logic [0:0] f1108_wen;
  logic [31:0] f1108_wdata;
  logic [0:0] f1108_clk;
  logic [0:0] f1108_rst;
  logic [31:0] f1108_rdata;
  sr_buffer_32_1 f1108(.wen(f1108_wen), .wdata(f1108_wdata), .clk(f1108_clk), .rst(f1108_rst), .rdata(f1108_rdata));
  assign f1108_clk = clk;
  assign f1108_rst = rst;
  // Bindings to f1108

  // f1106
  logic [0:0] f1106_wen;
  logic [31:0] f1106_wdata;
  logic [0:0] f1106_clk;
  logic [0:0] f1106_rst;
  logic [31:0] f1106_rdata;
  sr_buffer_32_1 f1106(.wen(f1106_wen), .wdata(f1106_wdata), .clk(f1106_clk), .rst(f1106_rst), .rdata(f1106_rdata));
  assign f1106_clk = clk;
  assign f1106_rst = rst;
  // Bindings to f1106

  // f1094
  logic [0:0] f1094_wen;
  logic [31:0] f1094_wdata;
  logic [0:0] f1094_clk;
  logic [0:0] f1094_rst;
  logic [31:0] f1094_rdata;
  sr_buffer_32_1 f1094(.wen(f1094_wen), .wdata(f1094_wdata), .clk(f1094_clk), .rst(f1094_rst), .rdata(f1094_rdata));
  assign f1094_clk = clk;
  assign f1094_rst = rst;
  // Bindings to f1094

  // f1104
  logic [0:0] f1104_wen;
  logic [31:0] f1104_wdata;
  logic [0:0] f1104_clk;
  logic [0:0] f1104_rst;
  logic [31:0] f1104_rdata;
  sr_buffer_32_1 f1104(.wen(f1104_wen), .wdata(f1104_wdata), .clk(f1104_clk), .rst(f1104_rst), .rdata(f1104_rdata));
  assign f1104_clk = clk;
  assign f1104_rst = rst;
  // Bindings to f1104

  // f1102
  logic [0:0] f1102_wen;
  logic [31:0] f1102_wdata;
  logic [0:0] f1102_clk;
  logic [0:0] f1102_rst;
  logic [31:0] f1102_rdata;
  sr_buffer_32_1 f1102(.wen(f1102_wen), .wdata(f1102_wdata), .clk(f1102_clk), .rst(f1102_rst), .rdata(f1102_rdata));
  assign f1102_clk = clk;
  assign f1102_rst = rst;
  // Bindings to f1102

  // f1100
  logic [0:0] f1100_wen;
  logic [31:0] f1100_wdata;
  logic [0:0] f1100_clk;
  logic [0:0] f1100_rst;
  logic [31:0] f1100_rdata;
  sr_buffer_32_1 f1100(.wen(f1100_wen), .wdata(f1100_wdata), .clk(f1100_clk), .rst(f1100_rst), .rdata(f1100_rdata));
  assign f1100_clk = clk;
  assign f1100_rst = rst;
  // Bindings to f1100

  // f1096
  logic [0:0] f1096_wen;
  logic [31:0] f1096_wdata;
  logic [0:0] f1096_clk;
  logic [0:0] f1096_rst;
  logic [31:0] f1096_rdata;
  sr_buffer_32_1 f1096(.wen(f1096_wen), .wdata(f1096_wdata), .clk(f1096_clk), .rst(f1096_rst), .rdata(f1096_rdata));
  assign f1096_clk = clk;
  assign f1096_rst = rst;
  // Bindings to f1096

  // f1098
  logic [0:0] f1098_wen;
  logic [31:0] f1098_wdata;
  logic [0:0] f1098_clk;
  logic [0:0] f1098_rst;
  logic [31:0] f1098_rdata;
  sr_buffer_32_1 f1098(.wen(f1098_wen), .wdata(f1098_wdata), .clk(f1098_clk), .rst(f1098_rst), .rdata(f1098_rdata));
  assign f1098_clk = clk;
  assign f1098_rst = rst;
  // Bindings to f1098

  // f1092
  logic [0:0] f1092_wen;
  logic [31:0] f1092_wdata;
  logic [0:0] f1092_clk;
  logic [0:0] f1092_rst;
  logic [31:0] f1092_rdata;
  sr_buffer_32_1 f1092(.wen(f1092_wen), .wdata(f1092_wdata), .clk(f1092_clk), .rst(f1092_rst), .rdata(f1092_rdata));
  assign f1092_clk = clk;
  assign f1092_rst = rst;
  // Bindings to f1092

  // f1090
  logic [0:0] f1090_wen;
  logic [31:0] f1090_wdata;
  logic [0:0] f1090_clk;
  logic [0:0] f1090_rst;
  logic [31:0] f1090_rdata;
  sr_buffer_32_1 f1090(.wen(f1090_wen), .wdata(f1090_wdata), .clk(f1090_clk), .rst(f1090_rst), .rdata(f1090_rdata));
  assign f1090_clk = clk;
  assign f1090_rst = rst;
  // Bindings to f1090

  // f1084
  logic [0:0] f1084_wen;
  logic [31:0] f1084_wdata;
  logic [0:0] f1084_clk;
  logic [0:0] f1084_rst;
  logic [31:0] f1084_rdata;
  sr_buffer_32_1 f1084(.wen(f1084_wen), .wdata(f1084_wdata), .clk(f1084_clk), .rst(f1084_rst), .rdata(f1084_rdata));
  assign f1084_clk = clk;
  assign f1084_rst = rst;
  // Bindings to f1084

  // f1088
  logic [0:0] f1088_wen;
  logic [31:0] f1088_wdata;
  logic [0:0] f1088_clk;
  logic [0:0] f1088_rst;
  logic [31:0] f1088_rdata;
  sr_buffer_32_1 f1088(.wen(f1088_wen), .wdata(f1088_wdata), .clk(f1088_clk), .rst(f1088_rst), .rdata(f1088_rdata));
  assign f1088_clk = clk;
  assign f1088_rst = rst;
  // Bindings to f1088

  // f1086
  logic [0:0] f1086_wen;
  logic [31:0] f1086_wdata;
  logic [0:0] f1086_clk;
  logic [0:0] f1086_rst;
  logic [31:0] f1086_rdata;
  sr_buffer_32_1 f1086(.wen(f1086_wen), .wdata(f1086_wdata), .clk(f1086_clk), .rst(f1086_rst), .rdata(f1086_rdata));
  assign f1086_clk = clk;
  assign f1086_rst = rst;
  // Bindings to f1086

  // f1080
  logic [0:0] f1080_wen;
  logic [31:0] f1080_wdata;
  logic [0:0] f1080_clk;
  logic [0:0] f1080_rst;
  logic [31:0] f1080_rdata;
  sr_buffer_32_1 f1080(.wen(f1080_wen), .wdata(f1080_wdata), .clk(f1080_clk), .rst(f1080_rst), .rdata(f1080_rdata));
  assign f1080_clk = clk;
  assign f1080_rst = rst;
  // Bindings to f1080

  // f1082
  logic [0:0] f1082_wen;
  logic [31:0] f1082_wdata;
  logic [0:0] f1082_clk;
  logic [0:0] f1082_rst;
  logic [31:0] f1082_rdata;
  sr_buffer_32_1 f1082(.wen(f1082_wen), .wdata(f1082_wdata), .clk(f1082_clk), .rst(f1082_rst), .rdata(f1082_rdata));
  assign f1082_clk = clk;
  assign f1082_rst = rst;
  // Bindings to f1082

  // f1078
  logic [0:0] f1078_wen;
  logic [31:0] f1078_wdata;
  logic [0:0] f1078_clk;
  logic [0:0] f1078_rst;
  logic [31:0] f1078_rdata;
  sr_buffer_32_1 f1078(.wen(f1078_wen), .wdata(f1078_wdata), .clk(f1078_clk), .rst(f1078_rst), .rdata(f1078_rdata));
  assign f1078_clk = clk;
  assign f1078_rst = rst;
  // Bindings to f1078

  // f1074
  logic [0:0] f1074_wen;
  logic [31:0] f1074_wdata;
  logic [0:0] f1074_clk;
  logic [0:0] f1074_rst;
  logic [31:0] f1074_rdata;
  sr_buffer_32_1 f1074(.wen(f1074_wen), .wdata(f1074_wdata), .clk(f1074_clk), .rst(f1074_rst), .rdata(f1074_rdata));
  assign f1074_clk = clk;
  assign f1074_rst = rst;
  // Bindings to f1074

  // f1076
  logic [0:0] f1076_wen;
  logic [31:0] f1076_wdata;
  logic [0:0] f1076_clk;
  logic [0:0] f1076_rst;
  logic [31:0] f1076_rdata;
  sr_buffer_32_1 f1076(.wen(f1076_wen), .wdata(f1076_wdata), .clk(f1076_clk), .rst(f1076_rst), .rdata(f1076_rdata));
  assign f1076_clk = clk;
  assign f1076_rst = rst;
  // Bindings to f1076

  // f1072
  logic [0:0] f1072_wen;
  logic [31:0] f1072_wdata;
  logic [0:0] f1072_clk;
  logic [0:0] f1072_rst;
  logic [31:0] f1072_rdata;
  sr_buffer_32_1 f1072(.wen(f1072_wen), .wdata(f1072_wdata), .clk(f1072_clk), .rst(f1072_rst), .rdata(f1072_rdata));
  assign f1072_clk = clk;
  assign f1072_rst = rst;
  // Bindings to f1072

  // f1060
  logic [0:0] f1060_wen;
  logic [31:0] f1060_wdata;
  logic [0:0] f1060_clk;
  logic [0:0] f1060_rst;
  logic [31:0] f1060_rdata;
  sr_buffer_32_1 f1060(.wen(f1060_wen), .wdata(f1060_wdata), .clk(f1060_clk), .rst(f1060_rst), .rdata(f1060_rdata));
  assign f1060_clk = clk;
  assign f1060_rst = rst;
  // Bindings to f1060

  // f1070
  logic [0:0] f1070_wen;
  logic [31:0] f1070_wdata;
  logic [0:0] f1070_clk;
  logic [0:0] f1070_rst;
  logic [31:0] f1070_rdata;
  sr_buffer_32_1 f1070(.wen(f1070_wen), .wdata(f1070_wdata), .clk(f1070_clk), .rst(f1070_rst), .rdata(f1070_rdata));
  assign f1070_clk = clk;
  assign f1070_rst = rst;
  // Bindings to f1070

  // f1068
  logic [0:0] f1068_wen;
  logic [31:0] f1068_wdata;
  logic [0:0] f1068_clk;
  logic [0:0] f1068_rst;
  logic [31:0] f1068_rdata;
  sr_buffer_32_1 f1068(.wen(f1068_wen), .wdata(f1068_wdata), .clk(f1068_clk), .rst(f1068_rst), .rdata(f1068_rdata));
  assign f1068_clk = clk;
  assign f1068_rst = rst;
  // Bindings to f1068

  // f1066
  logic [0:0] f1066_wen;
  logic [31:0] f1066_wdata;
  logic [0:0] f1066_clk;
  logic [0:0] f1066_rst;
  logic [31:0] f1066_rdata;
  sr_buffer_32_1 f1066(.wen(f1066_wen), .wdata(f1066_wdata), .clk(f1066_clk), .rst(f1066_rst), .rdata(f1066_rdata));
  assign f1066_clk = clk;
  assign f1066_rst = rst;
  // Bindings to f1066

  // f1062
  logic [0:0] f1062_wen;
  logic [31:0] f1062_wdata;
  logic [0:0] f1062_clk;
  logic [0:0] f1062_rst;
  logic [31:0] f1062_rdata;
  sr_buffer_32_1 f1062(.wen(f1062_wen), .wdata(f1062_wdata), .clk(f1062_clk), .rst(f1062_rst), .rdata(f1062_rdata));
  assign f1062_clk = clk;
  assign f1062_rst = rst;
  // Bindings to f1062

  // f1064
  logic [0:0] f1064_wen;
  logic [31:0] f1064_wdata;
  logic [0:0] f1064_clk;
  logic [0:0] f1064_rst;
  logic [31:0] f1064_rdata;
  sr_buffer_32_1 f1064(.wen(f1064_wen), .wdata(f1064_wdata), .clk(f1064_clk), .rst(f1064_rst), .rdata(f1064_rdata));
  assign f1064_clk = clk;
  assign f1064_rst = rst;
  // Bindings to f1064

  // f1058
  logic [0:0] f1058_wen;
  logic [31:0] f1058_wdata;
  logic [0:0] f1058_clk;
  logic [0:0] f1058_rst;
  logic [31:0] f1058_rdata;
  sr_buffer_32_1 f1058(.wen(f1058_wen), .wdata(f1058_wdata), .clk(f1058_clk), .rst(f1058_rst), .rdata(f1058_rdata));
  assign f1058_clk = clk;
  assign f1058_rst = rst;
  // Bindings to f1058

  // f1056
  logic [0:0] f1056_wen;
  logic [31:0] f1056_wdata;
  logic [0:0] f1056_clk;
  logic [0:0] f1056_rst;
  logic [31:0] f1056_rdata;
  sr_buffer_32_1 f1056(.wen(f1056_wen), .wdata(f1056_wdata), .clk(f1056_clk), .rst(f1056_rst), .rdata(f1056_rdata));
  assign f1056_clk = clk;
  assign f1056_rst = rst;
  // Bindings to f1056

  // f1054
  logic [0:0] f1054_wen;
  logic [31:0] f1054_wdata;
  logic [0:0] f1054_clk;
  logic [0:0] f1054_rst;
  logic [31:0] f1054_rdata;
  sr_buffer_32_1 f1054(.wen(f1054_wen), .wdata(f1054_wdata), .clk(f1054_clk), .rst(f1054_rst), .rdata(f1054_rdata));
  assign f1054_clk = clk;
  assign f1054_rst = rst;
  // Bindings to f1054

  // f1052
  logic [0:0] f1052_wen;
  logic [31:0] f1052_wdata;
  logic [0:0] f1052_clk;
  logic [0:0] f1052_rst;
  logic [31:0] f1052_rdata;
  sr_buffer_32_1 f1052(.wen(f1052_wen), .wdata(f1052_wdata), .clk(f1052_clk), .rst(f1052_rst), .rdata(f1052_rdata));
  assign f1052_clk = clk;
  assign f1052_rst = rst;
  // Bindings to f1052

  // f1048
  logic [0:0] f1048_wen;
  logic [31:0] f1048_wdata;
  logic [0:0] f1048_clk;
  logic [0:0] f1048_rst;
  logic [31:0] f1048_rdata;
  sr_buffer_32_1 f1048(.wen(f1048_wen), .wdata(f1048_wdata), .clk(f1048_clk), .rst(f1048_rst), .rdata(f1048_rdata));
  assign f1048_clk = clk;
  assign f1048_rst = rst;
  // Bindings to f1048

  // f1050
  logic [0:0] f1050_wen;
  logic [31:0] f1050_wdata;
  logic [0:0] f1050_clk;
  logic [0:0] f1050_rst;
  logic [31:0] f1050_rdata;
  sr_buffer_32_1 f1050(.wen(f1050_wen), .wdata(f1050_wdata), .clk(f1050_clk), .rst(f1050_rst), .rdata(f1050_rdata));
  assign f1050_clk = clk;
  assign f1050_rst = rst;
  // Bindings to f1050

  // f1046
  logic [0:0] f1046_wen;
  logic [31:0] f1046_wdata;
  logic [0:0] f1046_clk;
  logic [0:0] f1046_rst;
  logic [31:0] f1046_rdata;
  sr_buffer_32_1 f1046(.wen(f1046_wen), .wdata(f1046_wdata), .clk(f1046_clk), .rst(f1046_rst), .rdata(f1046_rdata));
  assign f1046_clk = clk;
  assign f1046_rst = rst;
  // Bindings to f1046

  // f1042
  logic [0:0] f1042_wen;
  logic [31:0] f1042_wdata;
  logic [0:0] f1042_clk;
  logic [0:0] f1042_rst;
  logic [31:0] f1042_rdata;
  sr_buffer_32_1 f1042(.wen(f1042_wen), .wdata(f1042_wdata), .clk(f1042_clk), .rst(f1042_rst), .rdata(f1042_rdata));
  assign f1042_clk = clk;
  assign f1042_rst = rst;
  // Bindings to f1042

  // f1044
  logic [0:0] f1044_wen;
  logic [31:0] f1044_wdata;
  logic [0:0] f1044_clk;
  logic [0:0] f1044_rst;
  logic [31:0] f1044_rdata;
  sr_buffer_32_1 f1044(.wen(f1044_wen), .wdata(f1044_wdata), .clk(f1044_clk), .rst(f1044_rst), .rdata(f1044_rdata));
  assign f1044_clk = clk;
  assign f1044_rst = rst;
  // Bindings to f1044

  // f1038
  logic [0:0] f1038_wen;
  logic [31:0] f1038_wdata;
  logic [0:0] f1038_clk;
  logic [0:0] f1038_rst;
  logic [31:0] f1038_rdata;
  sr_buffer_32_1 f1038(.wen(f1038_wen), .wdata(f1038_wdata), .clk(f1038_clk), .rst(f1038_rst), .rdata(f1038_rdata));
  assign f1038_clk = clk;
  assign f1038_rst = rst;
  // Bindings to f1038

  // f1040
  logic [0:0] f1040_wen;
  logic [31:0] f1040_wdata;
  logic [0:0] f1040_clk;
  logic [0:0] f1040_rst;
  logic [31:0] f1040_rdata;
  sr_buffer_32_1 f1040(.wen(f1040_wen), .wdata(f1040_wdata), .clk(f1040_clk), .rst(f1040_rst), .rdata(f1040_rdata));
  assign f1040_clk = clk;
  assign f1040_rst = rst;
  // Bindings to f1040

  // f1034
  logic [0:0] f1034_wen;
  logic [31:0] f1034_wdata;
  logic [0:0] f1034_clk;
  logic [0:0] f1034_rst;
  logic [31:0] f1034_rdata;
  sr_buffer_32_1 f1034(.wen(f1034_wen), .wdata(f1034_wdata), .clk(f1034_clk), .rst(f1034_rst), .rdata(f1034_rdata));
  assign f1034_clk = clk;
  assign f1034_rst = rst;
  // Bindings to f1034

  // f1036
  logic [0:0] f1036_wen;
  logic [31:0] f1036_wdata;
  logic [0:0] f1036_clk;
  logic [0:0] f1036_rst;
  logic [31:0] f1036_rdata;
  sr_buffer_32_1 f1036(.wen(f1036_wen), .wdata(f1036_wdata), .clk(f1036_clk), .rst(f1036_rst), .rdata(f1036_rdata));
  assign f1036_clk = clk;
  assign f1036_rst = rst;
  // Bindings to f1036

  // f1032
  logic [0:0] f1032_wen;
  logic [31:0] f1032_wdata;
  logic [0:0] f1032_clk;
  logic [0:0] f1032_rst;
  logic [31:0] f1032_rdata;
  sr_buffer_32_1 f1032(.wen(f1032_wen), .wdata(f1032_wdata), .clk(f1032_clk), .rst(f1032_rst), .rdata(f1032_rdata));
  assign f1032_clk = clk;
  assign f1032_rst = rst;
  // Bindings to f1032

  // f1030
  logic [0:0] f1030_wen;
  logic [31:0] f1030_wdata;
  logic [0:0] f1030_clk;
  logic [0:0] f1030_rst;
  logic [31:0] f1030_rdata;
  sr_buffer_32_1 f1030(.wen(f1030_wen), .wdata(f1030_wdata), .clk(f1030_clk), .rst(f1030_rst), .rdata(f1030_rdata));
  assign f1030_clk = clk;
  assign f1030_rst = rst;
  // Bindings to f1030

  // f1028
  logic [0:0] f1028_wen;
  logic [31:0] f1028_wdata;
  logic [0:0] f1028_clk;
  logic [0:0] f1028_rst;
  logic [31:0] f1028_rdata;
  sr_buffer_32_1 f1028(.wen(f1028_wen), .wdata(f1028_wdata), .clk(f1028_clk), .rst(f1028_rst), .rdata(f1028_rdata));
  assign f1028_clk = clk;
  assign f1028_rst = rst;
  // Bindings to f1028

  // f1026
  logic [0:0] f1026_wen;
  logic [31:0] f1026_wdata;
  logic [0:0] f1026_clk;
  logic [0:0] f1026_rst;
  logic [31:0] f1026_rdata;
  sr_buffer_32_1 f1026(.wen(f1026_wen), .wdata(f1026_wdata), .clk(f1026_clk), .rst(f1026_rst), .rdata(f1026_rdata));
  assign f1026_clk = clk;
  assign f1026_rst = rst;
  // Bindings to f1026

  // f1022
  logic [0:0] f1022_wen;
  logic [31:0] f1022_wdata;
  logic [0:0] f1022_clk;
  logic [0:0] f1022_rst;
  logic [31:0] f1022_rdata;
  sr_buffer_32_1 f1022(.wen(f1022_wen), .wdata(f1022_wdata), .clk(f1022_clk), .rst(f1022_rst), .rdata(f1022_rdata));
  assign f1022_clk = clk;
  assign f1022_rst = rst;
  // Bindings to f1022

  // f1024
  logic [0:0] f1024_wen;
  logic [31:0] f1024_wdata;
  logic [0:0] f1024_clk;
  logic [0:0] f1024_rst;
  logic [31:0] f1024_rdata;
  sr_buffer_32_1 f1024(.wen(f1024_wen), .wdata(f1024_wdata), .clk(f1024_clk), .rst(f1024_rst), .rdata(f1024_rdata));
  assign f1024_clk = clk;
  assign f1024_rst = rst;
  // Bindings to f1024

  // f1020
  logic [0:0] f1020_wen;
  logic [31:0] f1020_wdata;
  logic [0:0] f1020_clk;
  logic [0:0] f1020_rst;
  logic [31:0] f1020_rdata;
  sr_buffer_32_1 f1020(.wen(f1020_wen), .wdata(f1020_wdata), .clk(f1020_clk), .rst(f1020_rst), .rdata(f1020_rdata));
  assign f1020_clk = clk;
  assign f1020_rst = rst;
  // Bindings to f1020

  // f1018
  logic [0:0] f1018_wen;
  logic [31:0] f1018_wdata;
  logic [0:0] f1018_clk;
  logic [0:0] f1018_rst;
  logic [31:0] f1018_rdata;
  sr_buffer_32_1 f1018(.wen(f1018_wen), .wdata(f1018_wdata), .clk(f1018_clk), .rst(f1018_rst), .rdata(f1018_rdata));
  assign f1018_clk = clk;
  assign f1018_rst = rst;
  // Bindings to f1018

  // f1008
  logic [0:0] f1008_wen;
  logic [31:0] f1008_wdata;
  logic [0:0] f1008_clk;
  logic [0:0] f1008_rst;
  logic [31:0] f1008_rdata;
  sr_buffer_32_1 f1008(.wen(f1008_wen), .wdata(f1008_wdata), .clk(f1008_clk), .rst(f1008_rst), .rdata(f1008_rdata));
  assign f1008_clk = clk;
  assign f1008_rst = rst;
  // Bindings to f1008

  // f1016
  logic [0:0] f1016_wen;
  logic [31:0] f1016_wdata;
  logic [0:0] f1016_clk;
  logic [0:0] f1016_rst;
  logic [31:0] f1016_rdata;
  sr_buffer_32_1 f1016(.wen(f1016_wen), .wdata(f1016_wdata), .clk(f1016_clk), .rst(f1016_rst), .rdata(f1016_rdata));
  assign f1016_clk = clk;
  assign f1016_rst = rst;
  // Bindings to f1016

  // f1014
  logic [0:0] f1014_wen;
  logic [31:0] f1014_wdata;
  logic [0:0] f1014_clk;
  logic [0:0] f1014_rst;
  logic [31:0] f1014_rdata;
  sr_buffer_32_1 f1014(.wen(f1014_wen), .wdata(f1014_wdata), .clk(f1014_clk), .rst(f1014_rst), .rdata(f1014_rdata));
  assign f1014_clk = clk;
  assign f1014_rst = rst;
  // Bindings to f1014

  // f1010
  logic [0:0] f1010_wen;
  logic [31:0] f1010_wdata;
  logic [0:0] f1010_clk;
  logic [0:0] f1010_rst;
  logic [31:0] f1010_rdata;
  sr_buffer_32_1 f1010(.wen(f1010_wen), .wdata(f1010_wdata), .clk(f1010_clk), .rst(f1010_rst), .rdata(f1010_rdata));
  assign f1010_clk = clk;
  assign f1010_rst = rst;
  // Bindings to f1010

  // f1012
  logic [0:0] f1012_wen;
  logic [31:0] f1012_wdata;
  logic [0:0] f1012_clk;
  logic [0:0] f1012_rst;
  logic [31:0] f1012_rdata;
  sr_buffer_32_1 f1012(.wen(f1012_wen), .wdata(f1012_wdata), .clk(f1012_clk), .rst(f1012_rst), .rdata(f1012_rdata));
  assign f1012_clk = clk;
  assign f1012_rst = rst;
  // Bindings to f1012

  // f1004
  logic [0:0] f1004_wen;
  logic [31:0] f1004_wdata;
  logic [0:0] f1004_clk;
  logic [0:0] f1004_rst;
  logic [31:0] f1004_rdata;
  sr_buffer_32_1 f1004(.wen(f1004_wen), .wdata(f1004_wdata), .clk(f1004_clk), .rst(f1004_rst), .rdata(f1004_rdata));
  assign f1004_clk = clk;
  assign f1004_rst = rst;
  // Bindings to f1004

  // f1006
  logic [0:0] f1006_wen;
  logic [31:0] f1006_wdata;
  logic [0:0] f1006_clk;
  logic [0:0] f1006_rst;
  logic [31:0] f1006_rdata;
  sr_buffer_32_1 f1006(.wen(f1006_wen), .wdata(f1006_wdata), .clk(f1006_clk), .rst(f1006_rst), .rdata(f1006_rdata));
  assign f1006_clk = clk;
  assign f1006_rst = rst;
  // Bindings to f1006

  // f1002
  logic [0:0] f1002_wen;
  logic [31:0] f1002_wdata;
  logic [0:0] f1002_clk;
  logic [0:0] f1002_rst;
  logic [31:0] f1002_rdata;
  sr_buffer_32_1 f1002(.wen(f1002_wen), .wdata(f1002_wdata), .clk(f1002_clk), .rst(f1002_rst), .rdata(f1002_rdata));
  assign f1002_clk = clk;
  assign f1002_rst = rst;
  // Bindings to f1002

  // f1000
  logic [0:0] f1000_wen;
  logic [31:0] f1000_wdata;
  logic [0:0] f1000_clk;
  logic [0:0] f1000_rst;
  logic [31:0] f1000_rdata;
  sr_buffer_32_1 f1000(.wen(f1000_wen), .wdata(f1000_wdata), .clk(f1000_clk), .rst(f1000_rst), .rdata(f1000_rdata));
  assign f1000_clk = clk;
  assign f1000_rst = rst;
  // Bindings to f1000

  // f998
  logic [0:0] f998_wen;
  logic [31:0] f998_wdata;
  logic [0:0] f998_clk;
  logic [0:0] f998_rst;
  logic [31:0] f998_rdata;
  sr_buffer_32_1 f998(.wen(f998_wen), .wdata(f998_wdata), .clk(f998_clk), .rst(f998_rst), .rdata(f998_rdata));
  assign f998_clk = clk;
  assign f998_rst = rst;
  // Bindings to f998

  // f996
  logic [0:0] f996_wen;
  logic [31:0] f996_wdata;
  logic [0:0] f996_clk;
  logic [0:0] f996_rst;
  logic [31:0] f996_rdata;
  sr_buffer_32_1 f996(.wen(f996_wen), .wdata(f996_wdata), .clk(f996_clk), .rst(f996_rst), .rdata(f996_rdata));
  assign f996_clk = clk;
  assign f996_rst = rst;
  // Bindings to f996

  // f994
  logic [0:0] f994_wen;
  logic [31:0] f994_wdata;
  logic [0:0] f994_clk;
  logic [0:0] f994_rst;
  logic [31:0] f994_rdata;
  sr_buffer_32_1 f994(.wen(f994_wen), .wdata(f994_wdata), .clk(f994_clk), .rst(f994_rst), .rdata(f994_rdata));
  assign f994_clk = clk;
  assign f994_rst = rst;
  // Bindings to f994

  // f988
  logic [0:0] f988_wen;
  logic [31:0] f988_wdata;
  logic [0:0] f988_clk;
  logic [0:0] f988_rst;
  logic [31:0] f988_rdata;
  sr_buffer_32_1 f988(.wen(f988_wen), .wdata(f988_wdata), .clk(f988_clk), .rst(f988_rst), .rdata(f988_rdata));
  assign f988_clk = clk;
  assign f988_rst = rst;
  // Bindings to f988

  // f992
  logic [0:0] f992_wen;
  logic [31:0] f992_wdata;
  logic [0:0] f992_clk;
  logic [0:0] f992_rst;
  logic [31:0] f992_rdata;
  sr_buffer_32_1 f992(.wen(f992_wen), .wdata(f992_wdata), .clk(f992_clk), .rst(f992_rst), .rdata(f992_rdata));
  assign f992_clk = clk;
  assign f992_rst = rst;
  // Bindings to f992

  // f990
  logic [0:0] f990_wen;
  logic [31:0] f990_wdata;
  logic [0:0] f990_clk;
  logic [0:0] f990_rst;
  logic [31:0] f990_rdata;
  sr_buffer_32_1 f990(.wen(f990_wen), .wdata(f990_wdata), .clk(f990_clk), .rst(f990_rst), .rdata(f990_rdata));
  assign f990_clk = clk;
  assign f990_rst = rst;
  // Bindings to f990

  // f968
  logic [0:0] f968_wen;
  logic [31:0] f968_wdata;
  logic [0:0] f968_clk;
  logic [0:0] f968_rst;
  logic [31:0] f968_rdata;
  sr_buffer_32_1 f968(.wen(f968_wen), .wdata(f968_wdata), .clk(f968_clk), .rst(f968_rst), .rdata(f968_rdata));
  assign f968_clk = clk;
  assign f968_rst = rst;
  // Bindings to f968

  // f986
  logic [0:0] f986_wen;
  logic [31:0] f986_wdata;
  logic [0:0] f986_clk;
  logic [0:0] f986_rst;
  logic [31:0] f986_rdata;
  sr_buffer_32_1 f986(.wen(f986_wen), .wdata(f986_wdata), .clk(f986_clk), .rst(f986_rst), .rdata(f986_rdata));
  assign f986_clk = clk;
  assign f986_rst = rst;
  // Bindings to f986

  // f982
  logic [0:0] f982_wen;
  logic [31:0] f982_wdata;
  logic [0:0] f982_clk;
  logic [0:0] f982_rst;
  logic [31:0] f982_rdata;
  sr_buffer_32_1 f982(.wen(f982_wen), .wdata(f982_wdata), .clk(f982_clk), .rst(f982_rst), .rdata(f982_rdata));
  assign f982_clk = clk;
  assign f982_rst = rst;
  // Bindings to f982

  // f984
  logic [0:0] f984_wen;
  logic [31:0] f984_wdata;
  logic [0:0] f984_clk;
  logic [0:0] f984_rst;
  logic [31:0] f984_rdata;
  sr_buffer_32_1 f984(.wen(f984_wen), .wdata(f984_wdata), .clk(f984_clk), .rst(f984_rst), .rdata(f984_rdata));
  assign f984_clk = clk;
  assign f984_rst = rst;
  // Bindings to f984

  // f980
  logic [0:0] f980_wen;
  logic [31:0] f980_wdata;
  logic [0:0] f980_clk;
  logic [0:0] f980_rst;
  logic [31:0] f980_rdata;
  sr_buffer_32_1 f980(.wen(f980_wen), .wdata(f980_wdata), .clk(f980_clk), .rst(f980_rst), .rdata(f980_rdata));
  assign f980_clk = clk;
  assign f980_rst = rst;
  // Bindings to f980

  // f978
  logic [0:0] f978_wen;
  logic [31:0] f978_wdata;
  logic [0:0] f978_clk;
  logic [0:0] f978_rst;
  logic [31:0] f978_rdata;
  sr_buffer_32_1 f978(.wen(f978_wen), .wdata(f978_wdata), .clk(f978_clk), .rst(f978_rst), .rdata(f978_rdata));
  assign f978_clk = clk;
  assign f978_rst = rst;
  // Bindings to f978

  // f976
  logic [0:0] f976_wen;
  logic [31:0] f976_wdata;
  logic [0:0] f976_clk;
  logic [0:0] f976_rst;
  logic [31:0] f976_rdata;
  sr_buffer_32_1 f976(.wen(f976_wen), .wdata(f976_wdata), .clk(f976_clk), .rst(f976_rst), .rdata(f976_rdata));
  assign f976_clk = clk;
  assign f976_rst = rst;
  // Bindings to f976

  // f974
  logic [0:0] f974_wen;
  logic [31:0] f974_wdata;
  logic [0:0] f974_clk;
  logic [0:0] f974_rst;
  logic [31:0] f974_rdata;
  sr_buffer_32_1 f974(.wen(f974_wen), .wdata(f974_wdata), .clk(f974_clk), .rst(f974_rst), .rdata(f974_rdata));
  assign f974_clk = clk;
  assign f974_rst = rst;
  // Bindings to f974

  // f970
  logic [0:0] f970_wen;
  logic [31:0] f970_wdata;
  logic [0:0] f970_clk;
  logic [0:0] f970_rst;
  logic [31:0] f970_rdata;
  sr_buffer_32_1 f970(.wen(f970_wen), .wdata(f970_wdata), .clk(f970_clk), .rst(f970_rst), .rdata(f970_rdata));
  assign f970_clk = clk;
  assign f970_rst = rst;
  // Bindings to f970

  // f972
  logic [0:0] f972_wen;
  logic [31:0] f972_wdata;
  logic [0:0] f972_clk;
  logic [0:0] f972_rst;
  logic [31:0] f972_rdata;
  sr_buffer_32_1 f972(.wen(f972_wen), .wdata(f972_wdata), .clk(f972_clk), .rst(f972_rst), .rdata(f972_rdata));
  assign f972_clk = clk;
  assign f972_rst = rst;
  // Bindings to f972

  // f966
  logic [0:0] f966_wen;
  logic [31:0] f966_wdata;
  logic [0:0] f966_clk;
  logic [0:0] f966_rst;
  logic [31:0] f966_rdata;
  sr_buffer_32_1 f966(.wen(f966_wen), .wdata(f966_wdata), .clk(f966_clk), .rst(f966_rst), .rdata(f966_rdata));
  assign f966_clk = clk;
  assign f966_rst = rst;
  // Bindings to f966

  // f962
  logic [0:0] f962_wen;
  logic [31:0] f962_wdata;
  logic [0:0] f962_clk;
  logic [0:0] f962_rst;
  logic [31:0] f962_rdata;
  sr_buffer_32_1 f962(.wen(f962_wen), .wdata(f962_wdata), .clk(f962_clk), .rst(f962_rst), .rdata(f962_rdata));
  assign f962_clk = clk;
  assign f962_rst = rst;
  // Bindings to f962

  // f964
  logic [0:0] f964_wen;
  logic [31:0] f964_wdata;
  logic [0:0] f964_clk;
  logic [0:0] f964_rst;
  logic [31:0] f964_rdata;
  sr_buffer_32_1 f964(.wen(f964_wen), .wdata(f964_wdata), .clk(f964_clk), .rst(f964_rst), .rdata(f964_rdata));
  assign f964_clk = clk;
  assign f964_rst = rst;
  // Bindings to f964

  // f954
  logic [0:0] f954_wen;
  logic [31:0] f954_wdata;
  logic [0:0] f954_clk;
  logic [0:0] f954_rst;
  logic [31:0] f954_rdata;
  sr_buffer_32_1 f954(.wen(f954_wen), .wdata(f954_wdata), .clk(f954_clk), .rst(f954_rst), .rdata(f954_rdata));
  assign f954_clk = clk;
  assign f954_rst = rst;
  // Bindings to f954

  // f960
  logic [0:0] f960_wen;
  logic [31:0] f960_wdata;
  logic [0:0] f960_clk;
  logic [0:0] f960_rst;
  logic [31:0] f960_rdata;
  sr_buffer_32_1 f960(.wen(f960_wen), .wdata(f960_wdata), .clk(f960_clk), .rst(f960_rst), .rdata(f960_rdata));
  assign f960_clk = clk;
  assign f960_rst = rst;
  // Bindings to f960

  // f958
  logic [0:0] f958_wen;
  logic [31:0] f958_wdata;
  logic [0:0] f958_clk;
  logic [0:0] f958_rst;
  logic [31:0] f958_rdata;
  sr_buffer_32_1 f958(.wen(f958_wen), .wdata(f958_wdata), .clk(f958_clk), .rst(f958_rst), .rdata(f958_rdata));
  assign f958_clk = clk;
  assign f958_rst = rst;
  // Bindings to f958

  // f956
  logic [0:0] f956_wen;
  logic [31:0] f956_wdata;
  logic [0:0] f956_clk;
  logic [0:0] f956_rst;
  logic [31:0] f956_rdata;
  sr_buffer_32_1 f956(.wen(f956_wen), .wdata(f956_wdata), .clk(f956_clk), .rst(f956_rst), .rdata(f956_rdata));
  assign f956_clk = clk;
  assign f956_rst = rst;
  // Bindings to f956

  // f952
  logic [0:0] f952_wen;
  logic [31:0] f952_wdata;
  logic [0:0] f952_clk;
  logic [0:0] f952_rst;
  logic [31:0] f952_rdata;
  sr_buffer_32_1 f952(.wen(f952_wen), .wdata(f952_wdata), .clk(f952_clk), .rst(f952_rst), .rdata(f952_rdata));
  assign f952_clk = clk;
  assign f952_rst = rst;
  // Bindings to f952

  // f950
  logic [0:0] f950_wen;
  logic [31:0] f950_wdata;
  logic [0:0] f950_clk;
  logic [0:0] f950_rst;
  logic [31:0] f950_rdata;
  sr_buffer_32_1 f950(.wen(f950_wen), .wdata(f950_wdata), .clk(f950_clk), .rst(f950_rst), .rdata(f950_rdata));
  assign f950_clk = clk;
  assign f950_rst = rst;
  // Bindings to f950

  // f948
  logic [0:0] f948_wen;
  logic [31:0] f948_wdata;
  logic [0:0] f948_clk;
  logic [0:0] f948_rst;
  logic [31:0] f948_rdata;
  sr_buffer_32_1 f948(.wen(f948_wen), .wdata(f948_wdata), .clk(f948_clk), .rst(f948_rst), .rdata(f948_rdata));
  assign f948_clk = clk;
  assign f948_rst = rst;
  // Bindings to f948

  // f946
  logic [0:0] f946_wen;
  logic [31:0] f946_wdata;
  logic [0:0] f946_clk;
  logic [0:0] f946_rst;
  logic [31:0] f946_rdata;
  sr_buffer_32_1 f946(.wen(f946_wen), .wdata(f946_wdata), .clk(f946_clk), .rst(f946_rst), .rdata(f946_rdata));
  assign f946_clk = clk;
  assign f946_rst = rst;
  // Bindings to f946

  // f944
  logic [0:0] f944_wen;
  logic [31:0] f944_wdata;
  logic [0:0] f944_clk;
  logic [0:0] f944_rst;
  logic [31:0] f944_rdata;
  sr_buffer_32_1 f944(.wen(f944_wen), .wdata(f944_wdata), .clk(f944_clk), .rst(f944_rst), .rdata(f944_rdata));
  assign f944_clk = clk;
  assign f944_rst = rst;
  // Bindings to f944

  // f942
  logic [0:0] f942_wen;
  logic [31:0] f942_wdata;
  logic [0:0] f942_clk;
  logic [0:0] f942_rst;
  logic [31:0] f942_rdata;
  sr_buffer_32_1 f942(.wen(f942_wen), .wdata(f942_wdata), .clk(f942_clk), .rst(f942_rst), .rdata(f942_rdata));
  assign f942_clk = clk;
  assign f942_rst = rst;
  // Bindings to f942

  // f940
  logic [0:0] f940_wen;
  logic [31:0] f940_wdata;
  logic [0:0] f940_clk;
  logic [0:0] f940_rst;
  logic [31:0] f940_rdata;
  sr_buffer_32_1 f940(.wen(f940_wen), .wdata(f940_wdata), .clk(f940_clk), .rst(f940_rst), .rdata(f940_rdata));
  assign f940_clk = clk;
  assign f940_rst = rst;
  // Bindings to f940

  // f938
  logic [0:0] f938_wen;
  logic [31:0] f938_wdata;
  logic [0:0] f938_clk;
  logic [0:0] f938_rst;
  logic [31:0] f938_rdata;
  sr_buffer_32_1 f938(.wen(f938_wen), .wdata(f938_wdata), .clk(f938_clk), .rst(f938_rst), .rdata(f938_rdata));
  assign f938_clk = clk;
  assign f938_rst = rst;
  // Bindings to f938

  // f934
  logic [0:0] f934_wen;
  logic [31:0] f934_wdata;
  logic [0:0] f934_clk;
  logic [0:0] f934_rst;
  logic [31:0] f934_rdata;
  sr_buffer_32_1 f934(.wen(f934_wen), .wdata(f934_wdata), .clk(f934_clk), .rst(f934_rst), .rdata(f934_rdata));
  assign f934_clk = clk;
  assign f934_rst = rst;
  // Bindings to f934

  // f936
  logic [0:0] f936_wen;
  logic [31:0] f936_wdata;
  logic [0:0] f936_clk;
  logic [0:0] f936_rst;
  logic [31:0] f936_rdata;
  sr_buffer_32_1 f936(.wen(f936_wen), .wdata(f936_wdata), .clk(f936_clk), .rst(f936_rst), .rdata(f936_rdata));
  assign f936_clk = clk;
  assign f936_rst = rst;
  // Bindings to f936

  // f932
  logic [0:0] f932_wen;
  logic [31:0] f932_wdata;
  logic [0:0] f932_clk;
  logic [0:0] f932_rst;
  logic [31:0] f932_rdata;
  sr_buffer_32_1 f932(.wen(f932_wen), .wdata(f932_wdata), .clk(f932_clk), .rst(f932_rst), .rdata(f932_rdata));
  assign f932_clk = clk;
  assign f932_rst = rst;
  // Bindings to f932

  // f930
  logic [0:0] f930_wen;
  logic [31:0] f930_wdata;
  logic [0:0] f930_clk;
  logic [0:0] f930_rst;
  logic [31:0] f930_rdata;
  sr_buffer_32_1 f930(.wen(f930_wen), .wdata(f930_wdata), .clk(f930_clk), .rst(f930_rst), .rdata(f930_rdata));
  assign f930_clk = clk;
  assign f930_rst = rst;
  // Bindings to f930

  // f928
  logic [0:0] f928_wen;
  logic [31:0] f928_wdata;
  logic [0:0] f928_clk;
  logic [0:0] f928_rst;
  logic [31:0] f928_rdata;
  sr_buffer_32_1 f928(.wen(f928_wen), .wdata(f928_wdata), .clk(f928_clk), .rst(f928_rst), .rdata(f928_rdata));
  assign f928_clk = clk;
  assign f928_rst = rst;
  // Bindings to f928

  // f906
  logic [0:0] f906_wen;
  logic [31:0] f906_wdata;
  logic [0:0] f906_clk;
  logic [0:0] f906_rst;
  logic [31:0] f906_rdata;
  sr_buffer_32_1 f906(.wen(f906_wen), .wdata(f906_wdata), .clk(f906_clk), .rst(f906_rst), .rdata(f906_rdata));
  assign f906_clk = clk;
  assign f906_rst = rst;
  // Bindings to f906

  // f926
  logic [0:0] f926_wen;
  logic [31:0] f926_wdata;
  logic [0:0] f926_clk;
  logic [0:0] f926_rst;
  logic [31:0] f926_rdata;
  sr_buffer_32_1 f926(.wen(f926_wen), .wdata(f926_wdata), .clk(f926_clk), .rst(f926_rst), .rdata(f926_rdata));
  assign f926_clk = clk;
  assign f926_rst = rst;
  // Bindings to f926

  // f922
  logic [0:0] f922_wen;
  logic [31:0] f922_wdata;
  logic [0:0] f922_clk;
  logic [0:0] f922_rst;
  logic [31:0] f922_rdata;
  sr_buffer_32_1 f922(.wen(f922_wen), .wdata(f922_wdata), .clk(f922_clk), .rst(f922_rst), .rdata(f922_rdata));
  assign f922_clk = clk;
  assign f922_rst = rst;
  // Bindings to f922

  // f924
  logic [0:0] f924_wen;
  logic [31:0] f924_wdata;
  logic [0:0] f924_clk;
  logic [0:0] f924_rst;
  logic [31:0] f924_rdata;
  sr_buffer_32_1 f924(.wen(f924_wen), .wdata(f924_wdata), .clk(f924_clk), .rst(f924_rst), .rdata(f924_rdata));
  assign f924_clk = clk;
  assign f924_rst = rst;
  // Bindings to f924

  // f920
  logic [0:0] f920_wen;
  logic [31:0] f920_wdata;
  logic [0:0] f920_clk;
  logic [0:0] f920_rst;
  logic [31:0] f920_rdata;
  sr_buffer_32_1 f920(.wen(f920_wen), .wdata(f920_wdata), .clk(f920_clk), .rst(f920_rst), .rdata(f920_rdata));
  assign f920_clk = clk;
  assign f920_rst = rst;
  // Bindings to f920

  // f918
  logic [0:0] f918_wen;
  logic [31:0] f918_wdata;
  logic [0:0] f918_clk;
  logic [0:0] f918_rst;
  logic [31:0] f918_rdata;
  sr_buffer_32_1 f918(.wen(f918_wen), .wdata(f918_wdata), .clk(f918_clk), .rst(f918_rst), .rdata(f918_rdata));
  assign f918_clk = clk;
  assign f918_rst = rst;
  // Bindings to f918

  // f916
  logic [0:0] f916_wen;
  logic [31:0] f916_wdata;
  logic [0:0] f916_clk;
  logic [0:0] f916_rst;
  logic [31:0] f916_rdata;
  sr_buffer_32_1 f916(.wen(f916_wen), .wdata(f916_wdata), .clk(f916_clk), .rst(f916_rst), .rdata(f916_rdata));
  assign f916_clk = clk;
  assign f916_rst = rst;
  // Bindings to f916

  // f908
  logic [0:0] f908_wen;
  logic [31:0] f908_wdata;
  logic [0:0] f908_clk;
  logic [0:0] f908_rst;
  logic [31:0] f908_rdata;
  sr_buffer_32_1 f908(.wen(f908_wen), .wdata(f908_wdata), .clk(f908_clk), .rst(f908_rst), .rdata(f908_rdata));
  assign f908_clk = clk;
  assign f908_rst = rst;
  // Bindings to f908

  // f914
  logic [0:0] f914_wen;
  logic [31:0] f914_wdata;
  logic [0:0] f914_clk;
  logic [0:0] f914_rst;
  logic [31:0] f914_rdata;
  sr_buffer_32_1 f914(.wen(f914_wen), .wdata(f914_wdata), .clk(f914_clk), .rst(f914_rst), .rdata(f914_rdata));
  assign f914_clk = clk;
  assign f914_rst = rst;
  // Bindings to f914

  // f912
  logic [0:0] f912_wen;
  logic [31:0] f912_wdata;
  logic [0:0] f912_clk;
  logic [0:0] f912_rst;
  logic [31:0] f912_rdata;
  sr_buffer_32_1 f912(.wen(f912_wen), .wdata(f912_wdata), .clk(f912_clk), .rst(f912_rst), .rdata(f912_rdata));
  assign f912_clk = clk;
  assign f912_rst = rst;
  // Bindings to f912

  // f910
  logic [0:0] f910_wen;
  logic [31:0] f910_wdata;
  logic [0:0] f910_clk;
  logic [0:0] f910_rst;
  logic [31:0] f910_rdata;
  sr_buffer_32_1 f910(.wen(f910_wen), .wdata(f910_wdata), .clk(f910_clk), .rst(f910_rst), .rdata(f910_rdata));
  assign f910_clk = clk;
  assign f910_rst = rst;
  // Bindings to f910

  // f904
  logic [0:0] f904_wen;
  logic [31:0] f904_wdata;
  logic [0:0] f904_clk;
  logic [0:0] f904_rst;
  logic [31:0] f904_rdata;
  sr_buffer_32_1 f904(.wen(f904_wen), .wdata(f904_wdata), .clk(f904_clk), .rst(f904_rst), .rdata(f904_rdata));
  assign f904_clk = clk;
  assign f904_rst = rst;
  // Bindings to f904

  // f902
  logic [0:0] f902_wen;
  logic [31:0] f902_wdata;
  logic [0:0] f902_clk;
  logic [0:0] f902_rst;
  logic [31:0] f902_rdata;
  sr_buffer_32_1 f902(.wen(f902_wen), .wdata(f902_wdata), .clk(f902_clk), .rst(f902_rst), .rdata(f902_rdata));
  assign f902_clk = clk;
  assign f902_rst = rst;
  // Bindings to f902

  // f896
  logic [0:0] f896_wen;
  logic [31:0] f896_wdata;
  logic [0:0] f896_clk;
  logic [0:0] f896_rst;
  logic [31:0] f896_rdata;
  sr_buffer_32_1 f896(.wen(f896_wen), .wdata(f896_wdata), .clk(f896_clk), .rst(f896_rst), .rdata(f896_rdata));
  assign f896_clk = clk;
  assign f896_rst = rst;
  // Bindings to f896

  // f898
  logic [0:0] f898_wen;
  logic [31:0] f898_wdata;
  logic [0:0] f898_clk;
  logic [0:0] f898_rst;
  logic [31:0] f898_rdata;
  sr_buffer_32_1 f898(.wen(f898_wen), .wdata(f898_wdata), .clk(f898_clk), .rst(f898_rst), .rdata(f898_rdata));
  assign f898_clk = clk;
  assign f898_rst = rst;
  // Bindings to f898

  // f856
  logic [0:0] f856_wen;
  logic [31:0] f856_wdata;
  logic [0:0] f856_clk;
  logic [0:0] f856_rst;
  logic [31:0] f856_rdata;
  sr_buffer_32_1 f856(.wen(f856_wen), .wdata(f856_wdata), .clk(f856_clk), .rst(f856_rst), .rdata(f856_rdata));
  assign f856_clk = clk;
  assign f856_rst = rst;
  // Bindings to f856

  // f894
  logic [0:0] f894_wen;
  logic [31:0] f894_wdata;
  logic [0:0] f894_clk;
  logic [0:0] f894_rst;
  logic [31:0] f894_rdata;
  sr_buffer_32_1 f894(.wen(f894_wen), .wdata(f894_wdata), .clk(f894_clk), .rst(f894_rst), .rdata(f894_rdata));
  assign f894_clk = clk;
  assign f894_rst = rst;
  // Bindings to f894

  // f892
  logic [0:0] f892_wen;
  logic [31:0] f892_wdata;
  logic [0:0] f892_clk;
  logic [0:0] f892_rst;
  logic [31:0] f892_rdata;
  sr_buffer_32_1 f892(.wen(f892_wen), .wdata(f892_wdata), .clk(f892_clk), .rst(f892_rst), .rdata(f892_rdata));
  assign f892_clk = clk;
  assign f892_rst = rst;
  // Bindings to f892

  // f888
  logic [0:0] f888_wen;
  logic [31:0] f888_wdata;
  logic [0:0] f888_clk;
  logic [0:0] f888_rst;
  logic [31:0] f888_rdata;
  sr_buffer_32_1 f888(.wen(f888_wen), .wdata(f888_wdata), .clk(f888_clk), .rst(f888_rst), .rdata(f888_rdata));
  assign f888_clk = clk;
  assign f888_rst = rst;
  // Bindings to f888

  // f886
  logic [0:0] f886_wen;
  logic [31:0] f886_wdata;
  logic [0:0] f886_clk;
  logic [0:0] f886_rst;
  logic [31:0] f886_rdata;
  sr_buffer_32_1 f886(.wen(f886_wen), .wdata(f886_wdata), .clk(f886_clk), .rst(f886_rst), .rdata(f886_rdata));
  assign f886_clk = clk;
  assign f886_rst = rst;
  // Bindings to f886

  // f884
  logic [0:0] f884_wen;
  logic [31:0] f884_wdata;
  logic [0:0] f884_clk;
  logic [0:0] f884_rst;
  logic [31:0] f884_rdata;
  sr_buffer_32_1 f884(.wen(f884_wen), .wdata(f884_wdata), .clk(f884_clk), .rst(f884_rst), .rdata(f884_rdata));
  assign f884_clk = clk;
  assign f884_rst = rst;
  // Bindings to f884

  // f880
  logic [0:0] f880_wen;
  logic [31:0] f880_wdata;
  logic [0:0] f880_clk;
  logic [0:0] f880_rst;
  logic [31:0] f880_rdata;
  sr_buffer_32_1 f880(.wen(f880_wen), .wdata(f880_wdata), .clk(f880_clk), .rst(f880_rst), .rdata(f880_rdata));
  assign f880_clk = clk;
  assign f880_rst = rst;
  // Bindings to f880

  // f882
  logic [0:0] f882_wen;
  logic [31:0] f882_wdata;
  logic [0:0] f882_clk;
  logic [0:0] f882_rst;
  logic [31:0] f882_rdata;
  sr_buffer_32_1 f882(.wen(f882_wen), .wdata(f882_wdata), .clk(f882_clk), .rst(f882_rst), .rdata(f882_rdata));
  assign f882_clk = clk;
  assign f882_rst = rst;
  // Bindings to f882

  // f878
  logic [0:0] f878_wen;
  logic [31:0] f878_wdata;
  logic [0:0] f878_clk;
  logic [0:0] f878_rst;
  logic [31:0] f878_rdata;
  sr_buffer_32_1 f878(.wen(f878_wen), .wdata(f878_wdata), .clk(f878_clk), .rst(f878_rst), .rdata(f878_rdata));
  assign f878_clk = clk;
  assign f878_rst = rst;
  // Bindings to f878

  // f876
  logic [0:0] f876_wen;
  logic [31:0] f876_wdata;
  logic [0:0] f876_clk;
  logic [0:0] f876_rst;
  logic [31:0] f876_rdata;
  sr_buffer_32_1 f876(.wen(f876_wen), .wdata(f876_wdata), .clk(f876_clk), .rst(f876_rst), .rdata(f876_rdata));
  assign f876_clk = clk;
  assign f876_rst = rst;
  // Bindings to f876

  // f874
  logic [0:0] f874_wen;
  logic [31:0] f874_wdata;
  logic [0:0] f874_clk;
  logic [0:0] f874_rst;
  logic [31:0] f874_rdata;
  sr_buffer_32_1 f874(.wen(f874_wen), .wdata(f874_wdata), .clk(f874_clk), .rst(f874_rst), .rdata(f874_rdata));
  assign f874_clk = clk;
  assign f874_rst = rst;
  // Bindings to f874

  // f858
  logic [0:0] f858_wen;
  logic [31:0] f858_wdata;
  logic [0:0] f858_clk;
  logic [0:0] f858_rst;
  logic [31:0] f858_rdata;
  sr_buffer_32_1 f858(.wen(f858_wen), .wdata(f858_wdata), .clk(f858_clk), .rst(f858_rst), .rdata(f858_rdata));
  assign f858_clk = clk;
  assign f858_rst = rst;
  // Bindings to f858

  // f870
  logic [0:0] f870_wen;
  logic [31:0] f870_wdata;
  logic [0:0] f870_clk;
  logic [0:0] f870_rst;
  logic [31:0] f870_rdata;
  sr_buffer_32_1 f870(.wen(f870_wen), .wdata(f870_wdata), .clk(f870_clk), .rst(f870_rst), .rdata(f870_rdata));
  assign f870_clk = clk;
  assign f870_rst = rst;
  // Bindings to f870

  // f868
  logic [0:0] f868_wen;
  logic [31:0] f868_wdata;
  logic [0:0] f868_clk;
  logic [0:0] f868_rst;
  logic [31:0] f868_rdata;
  sr_buffer_32_1 f868(.wen(f868_wen), .wdata(f868_wdata), .clk(f868_clk), .rst(f868_rst), .rdata(f868_rdata));
  assign f868_clk = clk;
  assign f868_rst = rst;
  // Bindings to f868

  // f864
  logic [0:0] f864_wen;
  logic [31:0] f864_wdata;
  logic [0:0] f864_clk;
  logic [0:0] f864_rst;
  logic [31:0] f864_rdata;
  sr_buffer_32_1 f864(.wen(f864_wen), .wdata(f864_wdata), .clk(f864_clk), .rst(f864_rst), .rdata(f864_rdata));
  assign f864_clk = clk;
  assign f864_rst = rst;
  // Bindings to f864

  // f860
  logic [0:0] f860_wen;
  logic [31:0] f860_wdata;
  logic [0:0] f860_clk;
  logic [0:0] f860_rst;
  logic [31:0] f860_rdata;
  sr_buffer_32_1 f860(.wen(f860_wen), .wdata(f860_wdata), .clk(f860_clk), .rst(f860_rst), .rdata(f860_rdata));
  assign f860_clk = clk;
  assign f860_rst = rst;
  // Bindings to f860

  // f862
  logic [0:0] f862_wen;
  logic [31:0] f862_wdata;
  logic [0:0] f862_clk;
  logic [0:0] f862_rst;
  logic [31:0] f862_rdata;
  sr_buffer_32_1 f862(.wen(f862_wen), .wdata(f862_wdata), .clk(f862_clk), .rst(f862_rst), .rdata(f862_rdata));
  assign f862_clk = clk;
  assign f862_rst = rst;
  // Bindings to f862

  // f854
  logic [0:0] f854_wen;
  logic [31:0] f854_wdata;
  logic [0:0] f854_clk;
  logic [0:0] f854_rst;
  logic [31:0] f854_rdata;
  sr_buffer_32_1 f854(.wen(f854_wen), .wdata(f854_wdata), .clk(f854_clk), .rst(f854_rst), .rdata(f854_rdata));
  assign f854_clk = clk;
  assign f854_rst = rst;
  // Bindings to f854

  // f850
  logic [0:0] f850_wen;
  logic [31:0] f850_wdata;
  logic [0:0] f850_clk;
  logic [0:0] f850_rst;
  logic [31:0] f850_rdata;
  sr_buffer_32_1 f850(.wen(f850_wen), .wdata(f850_wdata), .clk(f850_clk), .rst(f850_rst), .rdata(f850_rdata));
  assign f850_clk = clk;
  assign f850_rst = rst;
  // Bindings to f850

  // f852
  logic [0:0] f852_wen;
  logic [31:0] f852_wdata;
  logic [0:0] f852_clk;
  logic [0:0] f852_rst;
  logic [31:0] f852_rdata;
  sr_buffer_32_1 f852(.wen(f852_wen), .wdata(f852_wdata), .clk(f852_clk), .rst(f852_rst), .rdata(f852_rdata));
  assign f852_clk = clk;
  assign f852_rst = rst;
  // Bindings to f852

  // f848
  logic [0:0] f848_wen;
  logic [31:0] f848_wdata;
  logic [0:0] f848_clk;
  logic [0:0] f848_rst;
  logic [31:0] f848_rdata;
  sr_buffer_32_1 f848(.wen(f848_wen), .wdata(f848_wdata), .clk(f848_clk), .rst(f848_rst), .rdata(f848_rdata));
  assign f848_clk = clk;
  assign f848_rst = rst;
  // Bindings to f848

  // f846
  logic [0:0] f846_wen;
  logic [31:0] f846_wdata;
  logic [0:0] f846_clk;
  logic [0:0] f846_rst;
  logic [31:0] f846_rdata;
  sr_buffer_32_1 f846(.wen(f846_wen), .wdata(f846_wdata), .clk(f846_clk), .rst(f846_rst), .rdata(f846_rdata));
  assign f846_clk = clk;
  assign f846_rst = rst;
  // Bindings to f846

  // f842
  logic [0:0] f842_wen;
  logic [31:0] f842_wdata;
  logic [0:0] f842_clk;
  logic [0:0] f842_rst;
  logic [31:0] f842_rdata;
  sr_buffer_32_1 f842(.wen(f842_wen), .wdata(f842_wdata), .clk(f842_clk), .rst(f842_rst), .rdata(f842_rdata));
  assign f842_clk = clk;
  assign f842_rst = rst;
  // Bindings to f842

  // f844
  logic [0:0] f844_wen;
  logic [31:0] f844_wdata;
  logic [0:0] f844_clk;
  logic [0:0] f844_rst;
  logic [31:0] f844_rdata;
  sr_buffer_32_1 f844(.wen(f844_wen), .wdata(f844_wdata), .clk(f844_clk), .rst(f844_rst), .rdata(f844_rdata));
  assign f844_clk = clk;
  assign f844_rst = rst;
  // Bindings to f844

  // f840
  logic [0:0] f840_wen;
  logic [31:0] f840_wdata;
  logic [0:0] f840_clk;
  logic [0:0] f840_rst;
  logic [31:0] f840_rdata;
  sr_buffer_32_1 f840(.wen(f840_wen), .wdata(f840_wdata), .clk(f840_clk), .rst(f840_rst), .rdata(f840_rdata));
  assign f840_clk = clk;
  assign f840_rst = rst;
  // Bindings to f840

  // f838
  logic [0:0] f838_wen;
  logic [31:0] f838_wdata;
  logic [0:0] f838_clk;
  logic [0:0] f838_rst;
  logic [31:0] f838_rdata;
  sr_buffer_32_1 f838(.wen(f838_wen), .wdata(f838_wdata), .clk(f838_clk), .rst(f838_rst), .rdata(f838_rdata));
  assign f838_clk = clk;
  assign f838_rst = rst;
  // Bindings to f838



endmodule


module bright_gauss_blur_2_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module bright_gauss_blur_2_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 633;
    end
  end

endmodule


module bright_gauss_blur_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1264;
    end
  end

endmodule


module bright_gauss_blur_2_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1263;
    end
  end

endmodule


module bright_gauss_blur_2_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 632;
    end
  end

endmodule


module bright_gauss_blur_2_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module bright_laplace_us_0_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (-1 + d1 == 0) ? ((4416 - floord(d0, 2))) : (d1 == 0) ? (3792) : ((-1 - d1) % 2 == 0 && -3 + d1 >= 0) ? ((4416 - floord(d0, 2))) : ((-d1) % 2 == 0 && -2 + d1 >= 0) ? (3792) : 0;
    end
  end

endmodule


module in_wire_bright_gauss_ds_1_update_0_write_wen(output [0:0] bright_gauss_ds_1_update_0_write_wen);

endmodule


module bright_gauss_blur_2_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (627 - d0 >= 0) ? (1262) : (-628 + d0 == 0) ? (1262) : 0;
    end
  end

endmodule


module bright_gauss_blur_2_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module bright_gauss_blur_2_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (627 - d0 >= 0) ? (631) : (-628 + d0 == 0) ? (631) : 0;
    end
  end

endmodule


module in_wire_bright_gauss_ds_1_update_0_write_wdata(output [31:0] bright_gauss_ds_1_update_0_write_wdata);

endmodule


module bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_312 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_312 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5



endmodule


module in_wire_bright_gauss_blur_2_update_0_read_dummy(output [287:0] bright_gauss_blur_2_update_0_read_dummy);

endmodule


module out_wire_bright_gauss_blur_2_update_0_read_rdata(input [287:0] bright_gauss_blur_2_update_0_read_rdata);

endmodule


module in_wire_bright_laplace_diff_1_update_0_read_dummy(output [31:0] bright_laplace_diff_1_update_0_read_dummy);

endmodule


module out_wire_bright_laplace_diff_1_update_0_read_rdata(input [31:0] bright_laplace_diff_1_update_0_read_rdata);

endmodule


module in_wire_bright_laplace_us_0_update_0_read_dummy(output [31:0] bright_laplace_us_0_update_0_read_dummy);

endmodule


module out_wire_bright_laplace_us_0_update_0_read_rdata(input [31:0] bright_laplace_us_0_update_0_read_rdata);

endmodule


module bright_gauss_blur_3_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (311 - d0 >= 0) ? (630) : (-312 + d0 == 0) ? (630) : 0;
    end
  end

endmodule


module sr_buffer_32_631(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 631;

  reg [31:0] data [630:0];

  reg [31:0] rdata_d;

  reg [9:0] waddr;

  wire [9:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module bright_gauss_blur_3_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 317;
    end
  end

endmodule


module bright_gauss_blur_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 632;
    end
  end

endmodule


module bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_631 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f314
  logic [0:0] f314_wen;
  logic [31:0] f314_wdata;
  logic [0:0] f314_clk;
  logic [0:0] f314_rst;
  logic [31:0] f314_rdata;
  sr_buffer_32_1 f314(.wen(f314_wen), .wdata(f314_wdata), .clk(f314_clk), .rst(f314_rst), .rdata(f314_rdata));
  assign f314_clk = clk;
  assign f314_rst = rst;
  // Bindings to f314

  // f316
  logic [0:0] f316_wen;
  logic [31:0] f316_wdata;
  logic [0:0] f316_clk;
  logic [0:0] f316_rst;
  logic [31:0] f316_rdata;
  sr_buffer_32_1 f316(.wen(f316_wen), .wdata(f316_wdata), .clk(f316_clk), .rst(f316_rst), .rdata(f316_rdata));
  assign f316_clk = clk;
  assign f316_rst = rst;
  // Bindings to f316

  // f318
  logic [0:0] f318_wen;
  logic [31:0] f318_wdata;
  logic [0:0] f318_clk;
  logic [0:0] f318_rst;
  logic [31:0] f318_rdata;
  sr_buffer_32_1 f318(.wen(f318_wen), .wdata(f318_wdata), .clk(f318_clk), .rst(f318_rst), .rdata(f318_rdata));
  assign f318_clk = clk;
  assign f318_rst = rst;
  // Bindings to f318

  // f320
  logic [0:0] f320_wen;
  logic [31:0] f320_wdata;
  logic [0:0] f320_clk;
  logic [0:0] f320_rst;
  logic [31:0] f320_rdata;
  sr_buffer_32_1 f320(.wen(f320_wen), .wdata(f320_wdata), .clk(f320_clk), .rst(f320_rst), .rdata(f320_rdata));
  assign f320_clk = clk;
  assign f320_rst = rst;
  // Bindings to f320

  // f322
  logic [0:0] f322_wen;
  logic [31:0] f322_wdata;
  logic [0:0] f322_clk;
  logic [0:0] f322_rst;
  logic [31:0] f322_rdata;
  sr_buffer_32_1 f322(.wen(f322_wen), .wdata(f322_wdata), .clk(f322_clk), .rst(f322_rst), .rdata(f322_rdata));
  assign f322_clk = clk;
  assign f322_rst = rst;
  // Bindings to f322

  // f324
  logic [0:0] f324_wen;
  logic [31:0] f324_wdata;
  logic [0:0] f324_clk;
  logic [0:0] f324_rst;
  logic [31:0] f324_rdata;
  sr_buffer_32_1 f324(.wen(f324_wen), .wdata(f324_wdata), .clk(f324_clk), .rst(f324_rst), .rdata(f324_rdata));
  assign f324_clk = clk;
  assign f324_rst = rst;
  // Bindings to f324

  // f326
  logic [0:0] f326_wen;
  logic [31:0] f326_wdata;
  logic [0:0] f326_clk;
  logic [0:0] f326_rst;
  logic [31:0] f326_rdata;
  sr_buffer_32_1 f326(.wen(f326_wen), .wdata(f326_wdata), .clk(f326_clk), .rst(f326_rst), .rdata(f326_rdata));
  assign f326_clk = clk;
  assign f326_rst = rst;
  // Bindings to f326

  // f328
  logic [0:0] f328_wen;
  logic [31:0] f328_wdata;
  logic [0:0] f328_clk;
  logic [0:0] f328_rst;
  logic [31:0] f328_rdata;
  sr_buffer_32_1 f328(.wen(f328_wen), .wdata(f328_wdata), .clk(f328_clk), .rst(f328_rst), .rdata(f328_rdata));
  assign f328_clk = clk;
  assign f328_rst = rst;
  // Bindings to f328

  // f330
  logic [0:0] f330_wen;
  logic [31:0] f330_wdata;
  logic [0:0] f330_clk;
  logic [0:0] f330_rst;
  logic [31:0] f330_rdata;
  sr_buffer_32_1 f330(.wen(f330_wen), .wdata(f330_wdata), .clk(f330_clk), .rst(f330_rst), .rdata(f330_rdata));
  assign f330_clk = clk;
  assign f330_rst = rst;
  // Bindings to f330

  // f332
  logic [0:0] f332_wen;
  logic [31:0] f332_wdata;
  logic [0:0] f332_clk;
  logic [0:0] f332_rst;
  logic [31:0] f332_rdata;
  sr_buffer_32_1 f332(.wen(f332_wen), .wdata(f332_wdata), .clk(f332_clk), .rst(f332_rst), .rdata(f332_rdata));
  assign f332_clk = clk;
  assign f332_rst = rst;
  // Bindings to f332

  // f334
  logic [0:0] f334_wen;
  logic [31:0] f334_wdata;
  logic [0:0] f334_clk;
  logic [0:0] f334_rst;
  logic [31:0] f334_rdata;
  sr_buffer_32_1 f334(.wen(f334_wen), .wdata(f334_wdata), .clk(f334_clk), .rst(f334_rst), .rdata(f334_rdata));
  assign f334_clk = clk;
  assign f334_rst = rst;
  // Bindings to f334

  // f336
  logic [0:0] f336_wen;
  logic [31:0] f336_wdata;
  logic [0:0] f336_clk;
  logic [0:0] f336_rst;
  logic [31:0] f336_rdata;
  sr_buffer_32_1 f336(.wen(f336_wen), .wdata(f336_wdata), .clk(f336_clk), .rst(f336_rst), .rdata(f336_rdata));
  assign f336_clk = clk;
  assign f336_rst = rst;
  // Bindings to f336

  // f338
  logic [0:0] f338_wen;
  logic [31:0] f338_wdata;
  logic [0:0] f338_clk;
  logic [0:0] f338_rst;
  logic [31:0] f338_rdata;
  sr_buffer_32_1 f338(.wen(f338_wen), .wdata(f338_wdata), .clk(f338_clk), .rst(f338_rst), .rdata(f338_rdata));
  assign f338_clk = clk;
  assign f338_rst = rst;
  // Bindings to f338

  // f340
  logic [0:0] f340_wen;
  logic [31:0] f340_wdata;
  logic [0:0] f340_clk;
  logic [0:0] f340_rst;
  logic [31:0] f340_rdata;
  sr_buffer_32_1 f340(.wen(f340_wen), .wdata(f340_wdata), .clk(f340_clk), .rst(f340_rst), .rdata(f340_rdata));
  assign f340_clk = clk;
  assign f340_rst = rst;
  // Bindings to f340

  // f342
  logic [0:0] f342_wen;
  logic [31:0] f342_wdata;
  logic [0:0] f342_clk;
  logic [0:0] f342_rst;
  logic [31:0] f342_rdata;
  sr_buffer_32_1 f342(.wen(f342_wen), .wdata(f342_wdata), .clk(f342_clk), .rst(f342_rst), .rdata(f342_rdata));
  assign f342_clk = clk;
  assign f342_rst = rst;
  // Bindings to f342

  // f344
  logic [0:0] f344_wen;
  logic [31:0] f344_wdata;
  logic [0:0] f344_clk;
  logic [0:0] f344_rst;
  logic [31:0] f344_rdata;
  sr_buffer_32_1 f344(.wen(f344_wen), .wdata(f344_wdata), .clk(f344_clk), .rst(f344_rst), .rdata(f344_rdata));
  assign f344_clk = clk;
  assign f344_rst = rst;
  // Bindings to f344

  // f346
  logic [0:0] f346_wen;
  logic [31:0] f346_wdata;
  logic [0:0] f346_clk;
  logic [0:0] f346_rst;
  logic [31:0] f346_rdata;
  sr_buffer_32_1 f346(.wen(f346_wen), .wdata(f346_wdata), .clk(f346_clk), .rst(f346_rst), .rdata(f346_rdata));
  assign f346_clk = clk;
  assign f346_rst = rst;
  // Bindings to f346

  // f348
  logic [0:0] f348_wen;
  logic [31:0] f348_wdata;
  logic [0:0] f348_clk;
  logic [0:0] f348_rst;
  logic [31:0] f348_rdata;
  sr_buffer_32_1 f348(.wen(f348_wen), .wdata(f348_wdata), .clk(f348_clk), .rst(f348_rst), .rdata(f348_rdata));
  assign f348_clk = clk;
  assign f348_rst = rst;
  // Bindings to f348

  // f350
  logic [0:0] f350_wen;
  logic [31:0] f350_wdata;
  logic [0:0] f350_clk;
  logic [0:0] f350_rst;
  logic [31:0] f350_rdata;
  sr_buffer_32_1 f350(.wen(f350_wen), .wdata(f350_wdata), .clk(f350_clk), .rst(f350_rst), .rdata(f350_rdata));
  assign f350_clk = clk;
  assign f350_rst = rst;
  // Bindings to f350

  // f352
  logic [0:0] f352_wen;
  logic [31:0] f352_wdata;
  logic [0:0] f352_clk;
  logic [0:0] f352_rst;
  logic [31:0] f352_rdata;
  sr_buffer_32_1 f352(.wen(f352_wen), .wdata(f352_wdata), .clk(f352_clk), .rst(f352_rst), .rdata(f352_rdata));
  assign f352_clk = clk;
  assign f352_rst = rst;
  // Bindings to f352

  // f354
  logic [0:0] f354_wen;
  logic [31:0] f354_wdata;
  logic [0:0] f354_clk;
  logic [0:0] f354_rst;
  logic [31:0] f354_rdata;
  sr_buffer_32_1 f354(.wen(f354_wen), .wdata(f354_wdata), .clk(f354_clk), .rst(f354_rst), .rdata(f354_rdata));
  assign f354_clk = clk;
  assign f354_rst = rst;
  // Bindings to f354

  // f356
  logic [0:0] f356_wen;
  logic [31:0] f356_wdata;
  logic [0:0] f356_clk;
  logic [0:0] f356_rst;
  logic [31:0] f356_rdata;
  sr_buffer_32_1 f356(.wen(f356_wen), .wdata(f356_wdata), .clk(f356_clk), .rst(f356_rst), .rdata(f356_rdata));
  assign f356_clk = clk;
  assign f356_rst = rst;
  // Bindings to f356

  // f358
  logic [0:0] f358_wen;
  logic [31:0] f358_wdata;
  logic [0:0] f358_clk;
  logic [0:0] f358_rst;
  logic [31:0] f358_rdata;
  sr_buffer_32_1 f358(.wen(f358_wen), .wdata(f358_wdata), .clk(f358_clk), .rst(f358_rst), .rdata(f358_rdata));
  assign f358_clk = clk;
  assign f358_rst = rst;
  // Bindings to f358

  // f360
  logic [0:0] f360_wen;
  logic [31:0] f360_wdata;
  logic [0:0] f360_clk;
  logic [0:0] f360_rst;
  logic [31:0] f360_rdata;
  sr_buffer_32_1 f360(.wen(f360_wen), .wdata(f360_wdata), .clk(f360_clk), .rst(f360_rst), .rdata(f360_rdata));
  assign f360_clk = clk;
  assign f360_rst = rst;
  // Bindings to f360

  // f362
  logic [0:0] f362_wen;
  logic [31:0] f362_wdata;
  logic [0:0] f362_clk;
  logic [0:0] f362_rst;
  logic [31:0] f362_rdata;
  sr_buffer_32_1 f362(.wen(f362_wen), .wdata(f362_wdata), .clk(f362_clk), .rst(f362_rst), .rdata(f362_rdata));
  assign f362_clk = clk;
  assign f362_rst = rst;
  // Bindings to f362

  // f364
  logic [0:0] f364_wen;
  logic [31:0] f364_wdata;
  logic [0:0] f364_clk;
  logic [0:0] f364_rst;
  logic [31:0] f364_rdata;
  sr_buffer_32_1 f364(.wen(f364_wen), .wdata(f364_wdata), .clk(f364_clk), .rst(f364_rst), .rdata(f364_rdata));
  assign f364_clk = clk;
  assign f364_rst = rst;
  // Bindings to f364

  // f366
  logic [0:0] f366_wen;
  logic [31:0] f366_wdata;
  logic [0:0] f366_clk;
  logic [0:0] f366_rst;
  logic [31:0] f366_rdata;
  sr_buffer_32_1 f366(.wen(f366_wen), .wdata(f366_wdata), .clk(f366_clk), .rst(f366_rst), .rdata(f366_rdata));
  assign f366_clk = clk;
  assign f366_rst = rst;
  // Bindings to f366

  // f368
  logic [0:0] f368_wen;
  logic [31:0] f368_wdata;
  logic [0:0] f368_clk;
  logic [0:0] f368_rst;
  logic [31:0] f368_rdata;
  sr_buffer_32_1 f368(.wen(f368_wen), .wdata(f368_wdata), .clk(f368_clk), .rst(f368_rst), .rdata(f368_rdata));
  assign f368_clk = clk;
  assign f368_rst = rst;
  // Bindings to f368

  // f370
  logic [0:0] f370_wen;
  logic [31:0] f370_wdata;
  logic [0:0] f370_clk;
  logic [0:0] f370_rst;
  logic [31:0] f370_rdata;
  sr_buffer_32_1 f370(.wen(f370_wen), .wdata(f370_wdata), .clk(f370_clk), .rst(f370_rst), .rdata(f370_rdata));
  assign f370_clk = clk;
  assign f370_rst = rst;
  // Bindings to f370

  // f372
  logic [0:0] f372_wen;
  logic [31:0] f372_wdata;
  logic [0:0] f372_clk;
  logic [0:0] f372_rst;
  logic [31:0] f372_rdata;
  sr_buffer_32_1 f372(.wen(f372_wen), .wdata(f372_wdata), .clk(f372_clk), .rst(f372_rst), .rdata(f372_rdata));
  assign f372_clk = clk;
  assign f372_rst = rst;
  // Bindings to f372

  // f374
  logic [0:0] f374_wen;
  logic [31:0] f374_wdata;
  logic [0:0] f374_clk;
  logic [0:0] f374_rst;
  logic [31:0] f374_rdata;
  sr_buffer_32_1 f374(.wen(f374_wen), .wdata(f374_wdata), .clk(f374_clk), .rst(f374_rst), .rdata(f374_rdata));
  assign f374_clk = clk;
  assign f374_rst = rst;
  // Bindings to f374

  // f376
  logic [0:0] f376_wen;
  logic [31:0] f376_wdata;
  logic [0:0] f376_clk;
  logic [0:0] f376_rst;
  logic [31:0] f376_rdata;
  sr_buffer_32_1 f376(.wen(f376_wen), .wdata(f376_wdata), .clk(f376_clk), .rst(f376_rst), .rdata(f376_rdata));
  assign f376_clk = clk;
  assign f376_rst = rst;
  // Bindings to f376

  // f378
  logic [0:0] f378_wen;
  logic [31:0] f378_wdata;
  logic [0:0] f378_clk;
  logic [0:0] f378_rst;
  logic [31:0] f378_rdata;
  sr_buffer_32_1 f378(.wen(f378_wen), .wdata(f378_wdata), .clk(f378_clk), .rst(f378_rst), .rdata(f378_rdata));
  assign f378_clk = clk;
  assign f378_rst = rst;
  // Bindings to f378

  // f380
  logic [0:0] f380_wen;
  logic [31:0] f380_wdata;
  logic [0:0] f380_clk;
  logic [0:0] f380_rst;
  logic [31:0] f380_rdata;
  sr_buffer_32_1 f380(.wen(f380_wen), .wdata(f380_wdata), .clk(f380_clk), .rst(f380_rst), .rdata(f380_rdata));
  assign f380_clk = clk;
  assign f380_rst = rst;
  // Bindings to f380

  // f382
  logic [0:0] f382_wen;
  logic [31:0] f382_wdata;
  logic [0:0] f382_clk;
  logic [0:0] f382_rst;
  logic [31:0] f382_rdata;
  sr_buffer_32_1 f382(.wen(f382_wen), .wdata(f382_wdata), .clk(f382_clk), .rst(f382_rst), .rdata(f382_rdata));
  assign f382_clk = clk;
  assign f382_rst = rst;
  // Bindings to f382

  // f384
  logic [0:0] f384_wen;
  logic [31:0] f384_wdata;
  logic [0:0] f384_clk;
  logic [0:0] f384_rst;
  logic [31:0] f384_rdata;
  sr_buffer_32_1 f384(.wen(f384_wen), .wdata(f384_wdata), .clk(f384_clk), .rst(f384_rst), .rdata(f384_rdata));
  assign f384_clk = clk;
  assign f384_rst = rst;
  // Bindings to f384

  // f386
  logic [0:0] f386_wen;
  logic [31:0] f386_wdata;
  logic [0:0] f386_clk;
  logic [0:0] f386_rst;
  logic [31:0] f386_rdata;
  sr_buffer_32_1 f386(.wen(f386_wen), .wdata(f386_wdata), .clk(f386_clk), .rst(f386_rst), .rdata(f386_rdata));
  assign f386_clk = clk;
  assign f386_rst = rst;
  // Bindings to f386

  // f388
  logic [0:0] f388_wen;
  logic [31:0] f388_wdata;
  logic [0:0] f388_clk;
  logic [0:0] f388_rst;
  logic [31:0] f388_rdata;
  sr_buffer_32_1 f388(.wen(f388_wen), .wdata(f388_wdata), .clk(f388_clk), .rst(f388_rst), .rdata(f388_rdata));
  assign f388_clk = clk;
  assign f388_rst = rst;
  // Bindings to f388

  // f390
  logic [0:0] f390_wen;
  logic [31:0] f390_wdata;
  logic [0:0] f390_clk;
  logic [0:0] f390_rst;
  logic [31:0] f390_rdata;
  sr_buffer_32_1 f390(.wen(f390_wen), .wdata(f390_wdata), .clk(f390_clk), .rst(f390_rst), .rdata(f390_rdata));
  assign f390_clk = clk;
  assign f390_rst = rst;
  // Bindings to f390

  // f392
  logic [0:0] f392_wen;
  logic [31:0] f392_wdata;
  logic [0:0] f392_clk;
  logic [0:0] f392_rst;
  logic [31:0] f392_rdata;
  sr_buffer_32_1 f392(.wen(f392_wen), .wdata(f392_wdata), .clk(f392_clk), .rst(f392_rst), .rdata(f392_rdata));
  assign f392_clk = clk;
  assign f392_rst = rst;
  // Bindings to f392

  // f394
  logic [0:0] f394_wen;
  logic [31:0] f394_wdata;
  logic [0:0] f394_clk;
  logic [0:0] f394_rst;
  logic [31:0] f394_rdata;
  sr_buffer_32_1 f394(.wen(f394_wen), .wdata(f394_wdata), .clk(f394_clk), .rst(f394_rst), .rdata(f394_rdata));
  assign f394_clk = clk;
  assign f394_rst = rst;
  // Bindings to f394

  // f396
  logic [0:0] f396_wen;
  logic [31:0] f396_wdata;
  logic [0:0] f396_clk;
  logic [0:0] f396_rst;
  logic [31:0] f396_rdata;
  sr_buffer_32_1 f396(.wen(f396_wen), .wdata(f396_wdata), .clk(f396_clk), .rst(f396_rst), .rdata(f396_rdata));
  assign f396_clk = clk;
  assign f396_rst = rst;
  // Bindings to f396

  // f398
  logic [0:0] f398_wen;
  logic [31:0] f398_wdata;
  logic [0:0] f398_clk;
  logic [0:0] f398_rst;
  logic [31:0] f398_rdata;
  sr_buffer_32_1 f398(.wen(f398_wen), .wdata(f398_wdata), .clk(f398_clk), .rst(f398_rst), .rdata(f398_rdata));
  assign f398_clk = clk;
  assign f398_rst = rst;
  // Bindings to f398

  // f400
  logic [0:0] f400_wen;
  logic [31:0] f400_wdata;
  logic [0:0] f400_clk;
  logic [0:0] f400_rst;
  logic [31:0] f400_rdata;
  sr_buffer_32_1 f400(.wen(f400_wen), .wdata(f400_wdata), .clk(f400_clk), .rst(f400_rst), .rdata(f400_rdata));
  assign f400_clk = clk;
  assign f400_rst = rst;
  // Bindings to f400

  // f402
  logic [0:0] f402_wen;
  logic [31:0] f402_wdata;
  logic [0:0] f402_clk;
  logic [0:0] f402_rst;
  logic [31:0] f402_rdata;
  sr_buffer_32_1 f402(.wen(f402_wen), .wdata(f402_wdata), .clk(f402_clk), .rst(f402_rst), .rdata(f402_rdata));
  assign f402_clk = clk;
  assign f402_rst = rst;
  // Bindings to f402

  // f404
  logic [0:0] f404_wen;
  logic [31:0] f404_wdata;
  logic [0:0] f404_clk;
  logic [0:0] f404_rst;
  logic [31:0] f404_rdata;
  sr_buffer_32_1 f404(.wen(f404_wen), .wdata(f404_wdata), .clk(f404_clk), .rst(f404_rst), .rdata(f404_rdata));
  assign f404_clk = clk;
  assign f404_rst = rst;
  // Bindings to f404

  // f406
  logic [0:0] f406_wen;
  logic [31:0] f406_wdata;
  logic [0:0] f406_clk;
  logic [0:0] f406_rst;
  logic [31:0] f406_rdata;
  sr_buffer_32_1 f406(.wen(f406_wen), .wdata(f406_wdata), .clk(f406_clk), .rst(f406_rst), .rdata(f406_rdata));
  assign f406_clk = clk;
  assign f406_rst = rst;
  // Bindings to f406

  // f408
  logic [0:0] f408_wen;
  logic [31:0] f408_wdata;
  logic [0:0] f408_clk;
  logic [0:0] f408_rst;
  logic [31:0] f408_rdata;
  sr_buffer_32_1 f408(.wen(f408_wen), .wdata(f408_wdata), .clk(f408_clk), .rst(f408_rst), .rdata(f408_rdata));
  assign f408_clk = clk;
  assign f408_rst = rst;
  // Bindings to f408

  // f410
  logic [0:0] f410_wen;
  logic [31:0] f410_wdata;
  logic [0:0] f410_clk;
  logic [0:0] f410_rst;
  logic [31:0] f410_rdata;
  sr_buffer_32_1 f410(.wen(f410_wen), .wdata(f410_wdata), .clk(f410_clk), .rst(f410_rst), .rdata(f410_rdata));
  assign f410_clk = clk;
  assign f410_rst = rst;
  // Bindings to f410

  // f412
  logic [0:0] f412_wen;
  logic [31:0] f412_wdata;
  logic [0:0] f412_clk;
  logic [0:0] f412_rst;
  logic [31:0] f412_rdata;
  sr_buffer_32_1 f412(.wen(f412_wen), .wdata(f412_wdata), .clk(f412_clk), .rst(f412_rst), .rdata(f412_rdata));
  assign f412_clk = clk;
  assign f412_rst = rst;
  // Bindings to f412

  // f414
  logic [0:0] f414_wen;
  logic [31:0] f414_wdata;
  logic [0:0] f414_clk;
  logic [0:0] f414_rst;
  logic [31:0] f414_rdata;
  sr_buffer_32_1 f414(.wen(f414_wen), .wdata(f414_wdata), .clk(f414_clk), .rst(f414_rst), .rdata(f414_rdata));
  assign f414_clk = clk;
  assign f414_rst = rst;
  // Bindings to f414

  // f416
  logic [0:0] f416_wen;
  logic [31:0] f416_wdata;
  logic [0:0] f416_clk;
  logic [0:0] f416_rst;
  logic [31:0] f416_rdata;
  sr_buffer_32_1 f416(.wen(f416_wen), .wdata(f416_wdata), .clk(f416_clk), .rst(f416_rst), .rdata(f416_rdata));
  assign f416_clk = clk;
  assign f416_rst = rst;
  // Bindings to f416

  // f418
  logic [0:0] f418_wen;
  logic [31:0] f418_wdata;
  logic [0:0] f418_clk;
  logic [0:0] f418_rst;
  logic [31:0] f418_rdata;
  sr_buffer_32_1 f418(.wen(f418_wen), .wdata(f418_wdata), .clk(f418_clk), .rst(f418_rst), .rdata(f418_rdata));
  assign f418_clk = clk;
  assign f418_rst = rst;
  // Bindings to f418

  // f420
  logic [0:0] f420_wen;
  logic [31:0] f420_wdata;
  logic [0:0] f420_clk;
  logic [0:0] f420_rst;
  logic [31:0] f420_rdata;
  sr_buffer_32_1 f420(.wen(f420_wen), .wdata(f420_wdata), .clk(f420_clk), .rst(f420_rst), .rdata(f420_rdata));
  assign f420_clk = clk;
  assign f420_rst = rst;
  // Bindings to f420

  // f422
  logic [0:0] f422_wen;
  logic [31:0] f422_wdata;
  logic [0:0] f422_clk;
  logic [0:0] f422_rst;
  logic [31:0] f422_rdata;
  sr_buffer_32_1 f422(.wen(f422_wen), .wdata(f422_wdata), .clk(f422_clk), .rst(f422_rst), .rdata(f422_rdata));
  assign f422_clk = clk;
  assign f422_rst = rst;
  // Bindings to f422

  // f424
  logic [0:0] f424_wen;
  logic [31:0] f424_wdata;
  logic [0:0] f424_clk;
  logic [0:0] f424_rst;
  logic [31:0] f424_rdata;
  sr_buffer_32_1 f424(.wen(f424_wen), .wdata(f424_wdata), .clk(f424_clk), .rst(f424_rst), .rdata(f424_rdata));
  assign f424_clk = clk;
  assign f424_rst = rst;
  // Bindings to f424

  // f426
  logic [0:0] f426_wen;
  logic [31:0] f426_wdata;
  logic [0:0] f426_clk;
  logic [0:0] f426_rst;
  logic [31:0] f426_rdata;
  sr_buffer_32_1 f426(.wen(f426_wen), .wdata(f426_wdata), .clk(f426_clk), .rst(f426_rst), .rdata(f426_rdata));
  assign f426_clk = clk;
  assign f426_rst = rst;
  // Bindings to f426

  // f428
  logic [0:0] f428_wen;
  logic [31:0] f428_wdata;
  logic [0:0] f428_clk;
  logic [0:0] f428_rst;
  logic [31:0] f428_rdata;
  sr_buffer_32_1 f428(.wen(f428_wen), .wdata(f428_wdata), .clk(f428_clk), .rst(f428_rst), .rdata(f428_rdata));
  assign f428_clk = clk;
  assign f428_rst = rst;
  // Bindings to f428

  // f430
  logic [0:0] f430_wen;
  logic [31:0] f430_wdata;
  logic [0:0] f430_clk;
  logic [0:0] f430_rst;
  logic [31:0] f430_rdata;
  sr_buffer_32_1 f430(.wen(f430_wen), .wdata(f430_wdata), .clk(f430_clk), .rst(f430_rst), .rdata(f430_rdata));
  assign f430_clk = clk;
  assign f430_rst = rst;
  // Bindings to f430

  // f432
  logic [0:0] f432_wen;
  logic [31:0] f432_wdata;
  logic [0:0] f432_clk;
  logic [0:0] f432_rst;
  logic [31:0] f432_rdata;
  sr_buffer_32_1 f432(.wen(f432_wen), .wdata(f432_wdata), .clk(f432_clk), .rst(f432_rst), .rdata(f432_rdata));
  assign f432_clk = clk;
  assign f432_rst = rst;
  // Bindings to f432

  // f434
  logic [0:0] f434_wen;
  logic [31:0] f434_wdata;
  logic [0:0] f434_clk;
  logic [0:0] f434_rst;
  logic [31:0] f434_rdata;
  sr_buffer_32_1 f434(.wen(f434_wen), .wdata(f434_wdata), .clk(f434_clk), .rst(f434_rst), .rdata(f434_rdata));
  assign f434_clk = clk;
  assign f434_rst = rst;
  // Bindings to f434

  // f436
  logic [0:0] f436_wen;
  logic [31:0] f436_wdata;
  logic [0:0] f436_clk;
  logic [0:0] f436_rst;
  logic [31:0] f436_rdata;
  sr_buffer_32_1 f436(.wen(f436_wen), .wdata(f436_wdata), .clk(f436_clk), .rst(f436_rst), .rdata(f436_rdata));
  assign f436_clk = clk;
  assign f436_rst = rst;
  // Bindings to f436

  // f438
  logic [0:0] f438_wen;
  logic [31:0] f438_wdata;
  logic [0:0] f438_clk;
  logic [0:0] f438_rst;
  logic [31:0] f438_rdata;
  sr_buffer_32_1 f438(.wen(f438_wen), .wdata(f438_wdata), .clk(f438_clk), .rst(f438_rst), .rdata(f438_rdata));
  assign f438_clk = clk;
  assign f438_rst = rst;
  // Bindings to f438

  // f440
  logic [0:0] f440_wen;
  logic [31:0] f440_wdata;
  logic [0:0] f440_clk;
  logic [0:0] f440_rst;
  logic [31:0] f440_rdata;
  sr_buffer_32_1 f440(.wen(f440_wen), .wdata(f440_wdata), .clk(f440_clk), .rst(f440_rst), .rdata(f440_rdata));
  assign f440_clk = clk;
  assign f440_rst = rst;
  // Bindings to f440

  // f442
  logic [0:0] f442_wen;
  logic [31:0] f442_wdata;
  logic [0:0] f442_clk;
  logic [0:0] f442_rst;
  logic [31:0] f442_rdata;
  sr_buffer_32_1 f442(.wen(f442_wen), .wdata(f442_wdata), .clk(f442_clk), .rst(f442_rst), .rdata(f442_rdata));
  assign f442_clk = clk;
  assign f442_rst = rst;
  // Bindings to f442

  // f444
  logic [0:0] f444_wen;
  logic [31:0] f444_wdata;
  logic [0:0] f444_clk;
  logic [0:0] f444_rst;
  logic [31:0] f444_rdata;
  sr_buffer_32_1 f444(.wen(f444_wen), .wdata(f444_wdata), .clk(f444_clk), .rst(f444_rst), .rdata(f444_rdata));
  assign f444_clk = clk;
  assign f444_rst = rst;
  // Bindings to f444

  // f446
  logic [0:0] f446_wen;
  logic [31:0] f446_wdata;
  logic [0:0] f446_clk;
  logic [0:0] f446_rst;
  logic [31:0] f446_rdata;
  sr_buffer_32_1 f446(.wen(f446_wen), .wdata(f446_wdata), .clk(f446_clk), .rst(f446_rst), .rdata(f446_rdata));
  assign f446_clk = clk;
  assign f446_rst = rst;
  // Bindings to f446

  // f448
  logic [0:0] f448_wen;
  logic [31:0] f448_wdata;
  logic [0:0] f448_clk;
  logic [0:0] f448_rst;
  logic [31:0] f448_rdata;
  sr_buffer_32_1 f448(.wen(f448_wen), .wdata(f448_wdata), .clk(f448_clk), .rst(f448_rst), .rdata(f448_rdata));
  assign f448_clk = clk;
  assign f448_rst = rst;
  // Bindings to f448

  // f450
  logic [0:0] f450_wen;
  logic [31:0] f450_wdata;
  logic [0:0] f450_clk;
  logic [0:0] f450_rst;
  logic [31:0] f450_rdata;
  sr_buffer_32_1 f450(.wen(f450_wen), .wdata(f450_wdata), .clk(f450_clk), .rst(f450_rst), .rdata(f450_rdata));
  assign f450_clk = clk;
  assign f450_rst = rst;
  // Bindings to f450

  // f452
  logic [0:0] f452_wen;
  logic [31:0] f452_wdata;
  logic [0:0] f452_clk;
  logic [0:0] f452_rst;
  logic [31:0] f452_rdata;
  sr_buffer_32_1 f452(.wen(f452_wen), .wdata(f452_wdata), .clk(f452_clk), .rst(f452_rst), .rdata(f452_rdata));
  assign f452_clk = clk;
  assign f452_rst = rst;
  // Bindings to f452

  // f454
  logic [0:0] f454_wen;
  logic [31:0] f454_wdata;
  logic [0:0] f454_clk;
  logic [0:0] f454_rst;
  logic [31:0] f454_rdata;
  sr_buffer_32_1 f454(.wen(f454_wen), .wdata(f454_wdata), .clk(f454_clk), .rst(f454_rst), .rdata(f454_rdata));
  assign f454_clk = clk;
  assign f454_rst = rst;
  // Bindings to f454

  // f456
  logic [0:0] f456_wen;
  logic [31:0] f456_wdata;
  logic [0:0] f456_clk;
  logic [0:0] f456_rst;
  logic [31:0] f456_rdata;
  sr_buffer_32_1 f456(.wen(f456_wen), .wdata(f456_wdata), .clk(f456_clk), .rst(f456_rst), .rdata(f456_rdata));
  assign f456_clk = clk;
  assign f456_rst = rst;
  // Bindings to f456

  // f458
  logic [0:0] f458_wen;
  logic [31:0] f458_wdata;
  logic [0:0] f458_clk;
  logic [0:0] f458_rst;
  logic [31:0] f458_rdata;
  sr_buffer_32_1 f458(.wen(f458_wen), .wdata(f458_wdata), .clk(f458_clk), .rst(f458_rst), .rdata(f458_rdata));
  assign f458_clk = clk;
  assign f458_rst = rst;
  // Bindings to f458

  // f460
  logic [0:0] f460_wen;
  logic [31:0] f460_wdata;
  logic [0:0] f460_clk;
  logic [0:0] f460_rst;
  logic [31:0] f460_rdata;
  sr_buffer_32_1 f460(.wen(f460_wen), .wdata(f460_wdata), .clk(f460_clk), .rst(f460_rst), .rdata(f460_rdata));
  assign f460_clk = clk;
  assign f460_rst = rst;
  // Bindings to f460

  // f462
  logic [0:0] f462_wen;
  logic [31:0] f462_wdata;
  logic [0:0] f462_clk;
  logic [0:0] f462_rst;
  logic [31:0] f462_rdata;
  sr_buffer_32_1 f462(.wen(f462_wen), .wdata(f462_wdata), .clk(f462_clk), .rst(f462_rst), .rdata(f462_rdata));
  assign f462_clk = clk;
  assign f462_rst = rst;
  // Bindings to f462

  // f464
  logic [0:0] f464_wen;
  logic [31:0] f464_wdata;
  logic [0:0] f464_clk;
  logic [0:0] f464_rst;
  logic [31:0] f464_rdata;
  sr_buffer_32_1 f464(.wen(f464_wen), .wdata(f464_wdata), .clk(f464_clk), .rst(f464_rst), .rdata(f464_rdata));
  assign f464_clk = clk;
  assign f464_rst = rst;
  // Bindings to f464

  // f466
  logic [0:0] f466_wen;
  logic [31:0] f466_wdata;
  logic [0:0] f466_clk;
  logic [0:0] f466_rst;
  logic [31:0] f466_rdata;
  sr_buffer_32_1 f466(.wen(f466_wen), .wdata(f466_wdata), .clk(f466_clk), .rst(f466_rst), .rdata(f466_rdata));
  assign f466_clk = clk;
  assign f466_rst = rst;
  // Bindings to f466

  // f468
  logic [0:0] f468_wen;
  logic [31:0] f468_wdata;
  logic [0:0] f468_clk;
  logic [0:0] f468_rst;
  logic [31:0] f468_rdata;
  sr_buffer_32_1 f468(.wen(f468_wen), .wdata(f468_wdata), .clk(f468_clk), .rst(f468_rst), .rdata(f468_rdata));
  assign f468_clk = clk;
  assign f468_rst = rst;
  // Bindings to f468

  // f470
  logic [0:0] f470_wen;
  logic [31:0] f470_wdata;
  logic [0:0] f470_clk;
  logic [0:0] f470_rst;
  logic [31:0] f470_rdata;
  sr_buffer_32_1 f470(.wen(f470_wen), .wdata(f470_wdata), .clk(f470_clk), .rst(f470_rst), .rdata(f470_rdata));
  assign f470_clk = clk;
  assign f470_rst = rst;
  // Bindings to f470

  // f472
  logic [0:0] f472_wen;
  logic [31:0] f472_wdata;
  logic [0:0] f472_clk;
  logic [0:0] f472_rst;
  logic [31:0] f472_rdata;
  sr_buffer_32_1 f472(.wen(f472_wen), .wdata(f472_wdata), .clk(f472_clk), .rst(f472_rst), .rdata(f472_rdata));
  assign f472_clk = clk;
  assign f472_rst = rst;
  // Bindings to f472

  // f474
  logic [0:0] f474_wen;
  logic [31:0] f474_wdata;
  logic [0:0] f474_clk;
  logic [0:0] f474_rst;
  logic [31:0] f474_rdata;
  sr_buffer_32_1 f474(.wen(f474_wen), .wdata(f474_wdata), .clk(f474_clk), .rst(f474_rst), .rdata(f474_rdata));
  assign f474_clk = clk;
  assign f474_rst = rst;
  // Bindings to f474

  // f476
  logic [0:0] f476_wen;
  logic [31:0] f476_wdata;
  logic [0:0] f476_clk;
  logic [0:0] f476_rst;
  logic [31:0] f476_rdata;
  sr_buffer_32_1 f476(.wen(f476_wen), .wdata(f476_wdata), .clk(f476_clk), .rst(f476_rst), .rdata(f476_rdata));
  assign f476_clk = clk;
  assign f476_rst = rst;
  // Bindings to f476

  // f478
  logic [0:0] f478_wen;
  logic [31:0] f478_wdata;
  logic [0:0] f478_clk;
  logic [0:0] f478_rst;
  logic [31:0] f478_rdata;
  sr_buffer_32_1 f478(.wen(f478_wen), .wdata(f478_wdata), .clk(f478_clk), .rst(f478_rst), .rdata(f478_rdata));
  assign f478_clk = clk;
  assign f478_rst = rst;
  // Bindings to f478

  // f480
  logic [0:0] f480_wen;
  logic [31:0] f480_wdata;
  logic [0:0] f480_clk;
  logic [0:0] f480_rst;
  logic [31:0] f480_rdata;
  sr_buffer_32_1 f480(.wen(f480_wen), .wdata(f480_wdata), .clk(f480_clk), .rst(f480_rst), .rdata(f480_rdata));
  assign f480_clk = clk;
  assign f480_rst = rst;
  // Bindings to f480

  // f482
  logic [0:0] f482_wen;
  logic [31:0] f482_wdata;
  logic [0:0] f482_clk;
  logic [0:0] f482_rst;
  logic [31:0] f482_rdata;
  sr_buffer_32_1 f482(.wen(f482_wen), .wdata(f482_wdata), .clk(f482_clk), .rst(f482_rst), .rdata(f482_rdata));
  assign f482_clk = clk;
  assign f482_rst = rst;
  // Bindings to f482

  // f484
  logic [0:0] f484_wen;
  logic [31:0] f484_wdata;
  logic [0:0] f484_clk;
  logic [0:0] f484_rst;
  logic [31:0] f484_rdata;
  sr_buffer_32_1 f484(.wen(f484_wen), .wdata(f484_wdata), .clk(f484_clk), .rst(f484_rst), .rdata(f484_rdata));
  assign f484_clk = clk;
  assign f484_rst = rst;
  // Bindings to f484

  // f486
  logic [0:0] f486_wen;
  logic [31:0] f486_wdata;
  logic [0:0] f486_clk;
  logic [0:0] f486_rst;
  logic [31:0] f486_rdata;
  sr_buffer_32_1 f486(.wen(f486_wen), .wdata(f486_wdata), .clk(f486_clk), .rst(f486_rst), .rdata(f486_rdata));
  assign f486_clk = clk;
  assign f486_rst = rst;
  // Bindings to f486

  // f488
  logic [0:0] f488_wen;
  logic [31:0] f488_wdata;
  logic [0:0] f488_clk;
  logic [0:0] f488_rst;
  logic [31:0] f488_rdata;
  sr_buffer_32_1 f488(.wen(f488_wen), .wdata(f488_wdata), .clk(f488_clk), .rst(f488_rst), .rdata(f488_rdata));
  assign f488_clk = clk;
  assign f488_rst = rst;
  // Bindings to f488

  // f490
  logic [0:0] f490_wen;
  logic [31:0] f490_wdata;
  logic [0:0] f490_clk;
  logic [0:0] f490_rst;
  logic [31:0] f490_rdata;
  sr_buffer_32_1 f490(.wen(f490_wen), .wdata(f490_wdata), .clk(f490_clk), .rst(f490_rst), .rdata(f490_rdata));
  assign f490_clk = clk;
  assign f490_rst = rst;
  // Bindings to f490

  // f492
  logic [0:0] f492_wen;
  logic [31:0] f492_wdata;
  logic [0:0] f492_clk;
  logic [0:0] f492_rst;
  logic [31:0] f492_rdata;
  sr_buffer_32_1 f492(.wen(f492_wen), .wdata(f492_wdata), .clk(f492_clk), .rst(f492_rst), .rdata(f492_rdata));
  assign f492_clk = clk;
  assign f492_rst = rst;
  // Bindings to f492

  // f494
  logic [0:0] f494_wen;
  logic [31:0] f494_wdata;
  logic [0:0] f494_clk;
  logic [0:0] f494_rst;
  logic [31:0] f494_rdata;
  sr_buffer_32_1 f494(.wen(f494_wen), .wdata(f494_wdata), .clk(f494_clk), .rst(f494_rst), .rdata(f494_rdata));
  assign f494_clk = clk;
  assign f494_rst = rst;
  // Bindings to f494

  // f496
  logic [0:0] f496_wen;
  logic [31:0] f496_wdata;
  logic [0:0] f496_clk;
  logic [0:0] f496_rst;
  logic [31:0] f496_rdata;
  sr_buffer_32_1 f496(.wen(f496_wen), .wdata(f496_wdata), .clk(f496_clk), .rst(f496_rst), .rdata(f496_rdata));
  assign f496_clk = clk;
  assign f496_rst = rst;
  // Bindings to f496

  // f498
  logic [0:0] f498_wen;
  logic [31:0] f498_wdata;
  logic [0:0] f498_clk;
  logic [0:0] f498_rst;
  logic [31:0] f498_rdata;
  sr_buffer_32_1 f498(.wen(f498_wen), .wdata(f498_wdata), .clk(f498_clk), .rst(f498_rst), .rdata(f498_rdata));
  assign f498_clk = clk;
  assign f498_rst = rst;
  // Bindings to f498

  // f500
  logic [0:0] f500_wen;
  logic [31:0] f500_wdata;
  logic [0:0] f500_clk;
  logic [0:0] f500_rst;
  logic [31:0] f500_rdata;
  sr_buffer_32_1 f500(.wen(f500_wen), .wdata(f500_wdata), .clk(f500_clk), .rst(f500_rst), .rdata(f500_rdata));
  assign f500_clk = clk;
  assign f500_rst = rst;
  // Bindings to f500

  // f502
  logic [0:0] f502_wen;
  logic [31:0] f502_wdata;
  logic [0:0] f502_clk;
  logic [0:0] f502_rst;
  logic [31:0] f502_rdata;
  sr_buffer_32_1 f502(.wen(f502_wen), .wdata(f502_wdata), .clk(f502_clk), .rst(f502_rst), .rdata(f502_rdata));
  assign f502_clk = clk;
  assign f502_rst = rst;
  // Bindings to f502

  // f504
  logic [0:0] f504_wen;
  logic [31:0] f504_wdata;
  logic [0:0] f504_clk;
  logic [0:0] f504_rst;
  logic [31:0] f504_rdata;
  sr_buffer_32_1 f504(.wen(f504_wen), .wdata(f504_wdata), .clk(f504_clk), .rst(f504_rst), .rdata(f504_rdata));
  assign f504_clk = clk;
  assign f504_rst = rst;
  // Bindings to f504

  // f506
  logic [0:0] f506_wen;
  logic [31:0] f506_wdata;
  logic [0:0] f506_clk;
  logic [0:0] f506_rst;
  logic [31:0] f506_rdata;
  sr_buffer_32_1 f506(.wen(f506_wen), .wdata(f506_wdata), .clk(f506_clk), .rst(f506_rst), .rdata(f506_rdata));
  assign f506_clk = clk;
  assign f506_rst = rst;
  // Bindings to f506

  // f508
  logic [0:0] f508_wen;
  logic [31:0] f508_wdata;
  logic [0:0] f508_clk;
  logic [0:0] f508_rst;
  logic [31:0] f508_rdata;
  sr_buffer_32_1 f508(.wen(f508_wen), .wdata(f508_wdata), .clk(f508_clk), .rst(f508_rst), .rdata(f508_rdata));
  assign f508_clk = clk;
  assign f508_rst = rst;
  // Bindings to f508

  // f510
  logic [0:0] f510_wen;
  logic [31:0] f510_wdata;
  logic [0:0] f510_clk;
  logic [0:0] f510_rst;
  logic [31:0] f510_rdata;
  sr_buffer_32_1 f510(.wen(f510_wen), .wdata(f510_wdata), .clk(f510_clk), .rst(f510_rst), .rdata(f510_rdata));
  assign f510_clk = clk;
  assign f510_rst = rst;
  // Bindings to f510

  // f512
  logic [0:0] f512_wen;
  logic [31:0] f512_wdata;
  logic [0:0] f512_clk;
  logic [0:0] f512_rst;
  logic [31:0] f512_rdata;
  sr_buffer_32_1 f512(.wen(f512_wen), .wdata(f512_wdata), .clk(f512_clk), .rst(f512_rst), .rdata(f512_rdata));
  assign f512_clk = clk;
  assign f512_rst = rst;
  // Bindings to f512

  // f514
  logic [0:0] f514_wen;
  logic [31:0] f514_wdata;
  logic [0:0] f514_clk;
  logic [0:0] f514_rst;
  logic [31:0] f514_rdata;
  sr_buffer_32_1 f514(.wen(f514_wen), .wdata(f514_wdata), .clk(f514_clk), .rst(f514_rst), .rdata(f514_rdata));
  assign f514_clk = clk;
  assign f514_rst = rst;
  // Bindings to f514

  // f516
  logic [0:0] f516_wen;
  logic [31:0] f516_wdata;
  logic [0:0] f516_clk;
  logic [0:0] f516_rst;
  logic [31:0] f516_rdata;
  sr_buffer_32_1 f516(.wen(f516_wen), .wdata(f516_wdata), .clk(f516_clk), .rst(f516_rst), .rdata(f516_rdata));
  assign f516_clk = clk;
  assign f516_rst = rst;
  // Bindings to f516

  // f518
  logic [0:0] f518_wen;
  logic [31:0] f518_wdata;
  logic [0:0] f518_clk;
  logic [0:0] f518_rst;
  logic [31:0] f518_rdata;
  sr_buffer_32_1 f518(.wen(f518_wen), .wdata(f518_wdata), .clk(f518_clk), .rst(f518_rst), .rdata(f518_rdata));
  assign f518_clk = clk;
  assign f518_rst = rst;
  // Bindings to f518

  // f520
  logic [0:0] f520_wen;
  logic [31:0] f520_wdata;
  logic [0:0] f520_clk;
  logic [0:0] f520_rst;
  logic [31:0] f520_rdata;
  sr_buffer_32_1 f520(.wen(f520_wen), .wdata(f520_wdata), .clk(f520_clk), .rst(f520_rst), .rdata(f520_rdata));
  assign f520_clk = clk;
  assign f520_rst = rst;
  // Bindings to f520

  // f522
  logic [0:0] f522_wen;
  logic [31:0] f522_wdata;
  logic [0:0] f522_clk;
  logic [0:0] f522_rst;
  logic [31:0] f522_rdata;
  sr_buffer_32_1 f522(.wen(f522_wen), .wdata(f522_wdata), .clk(f522_clk), .rst(f522_rst), .rdata(f522_rdata));
  assign f522_clk = clk;
  assign f522_rst = rst;
  // Bindings to f522

  // f524
  logic [0:0] f524_wen;
  logic [31:0] f524_wdata;
  logic [0:0] f524_clk;
  logic [0:0] f524_rst;
  logic [31:0] f524_rdata;
  sr_buffer_32_1 f524(.wen(f524_wen), .wdata(f524_wdata), .clk(f524_clk), .rst(f524_rst), .rdata(f524_rdata));
  assign f524_clk = clk;
  assign f524_rst = rst;
  // Bindings to f524

  // f526
  logic [0:0] f526_wen;
  logic [31:0] f526_wdata;
  logic [0:0] f526_clk;
  logic [0:0] f526_rst;
  logic [31:0] f526_rdata;
  sr_buffer_32_1 f526(.wen(f526_wen), .wdata(f526_wdata), .clk(f526_clk), .rst(f526_rst), .rdata(f526_rdata));
  assign f526_clk = clk;
  assign f526_rst = rst;
  // Bindings to f526

  // f528
  logic [0:0] f528_wen;
  logic [31:0] f528_wdata;
  logic [0:0] f528_clk;
  logic [0:0] f528_rst;
  logic [31:0] f528_rdata;
  sr_buffer_32_1 f528(.wen(f528_wen), .wdata(f528_wdata), .clk(f528_clk), .rst(f528_rst), .rdata(f528_rdata));
  assign f528_clk = clk;
  assign f528_rst = rst;
  // Bindings to f528

  // f530
  logic [0:0] f530_wen;
  logic [31:0] f530_wdata;
  logic [0:0] f530_clk;
  logic [0:0] f530_rst;
  logic [31:0] f530_rdata;
  sr_buffer_32_1 f530(.wen(f530_wen), .wdata(f530_wdata), .clk(f530_clk), .rst(f530_rst), .rdata(f530_rdata));
  assign f530_clk = clk;
  assign f530_rst = rst;
  // Bindings to f530

  // f532
  logic [0:0] f532_wen;
  logic [31:0] f532_wdata;
  logic [0:0] f532_clk;
  logic [0:0] f532_rst;
  logic [31:0] f532_rdata;
  sr_buffer_32_1 f532(.wen(f532_wen), .wdata(f532_wdata), .clk(f532_clk), .rst(f532_rst), .rdata(f532_rdata));
  assign f532_clk = clk;
  assign f532_rst = rst;
  // Bindings to f532

  // f534
  logic [0:0] f534_wen;
  logic [31:0] f534_wdata;
  logic [0:0] f534_clk;
  logic [0:0] f534_rst;
  logic [31:0] f534_rdata;
  sr_buffer_32_1 f534(.wen(f534_wen), .wdata(f534_wdata), .clk(f534_clk), .rst(f534_rst), .rdata(f534_rdata));
  assign f534_clk = clk;
  assign f534_rst = rst;
  // Bindings to f534

  // f536
  logic [0:0] f536_wen;
  logic [31:0] f536_wdata;
  logic [0:0] f536_clk;
  logic [0:0] f536_rst;
  logic [31:0] f536_rdata;
  sr_buffer_32_1 f536(.wen(f536_wen), .wdata(f536_wdata), .clk(f536_clk), .rst(f536_rst), .rdata(f536_rdata));
  assign f536_clk = clk;
  assign f536_rst = rst;
  // Bindings to f536

  // f538
  logic [0:0] f538_wen;
  logic [31:0] f538_wdata;
  logic [0:0] f538_clk;
  logic [0:0] f538_rst;
  logic [31:0] f538_rdata;
  sr_buffer_32_1 f538(.wen(f538_wen), .wdata(f538_wdata), .clk(f538_clk), .rst(f538_rst), .rdata(f538_rdata));
  assign f538_clk = clk;
  assign f538_rst = rst;
  // Bindings to f538

  // f540
  logic [0:0] f540_wen;
  logic [31:0] f540_wdata;
  logic [0:0] f540_clk;
  logic [0:0] f540_rst;
  logic [31:0] f540_rdata;
  sr_buffer_32_1 f540(.wen(f540_wen), .wdata(f540_wdata), .clk(f540_clk), .rst(f540_rst), .rdata(f540_rdata));
  assign f540_clk = clk;
  assign f540_rst = rst;
  // Bindings to f540

  // f542
  logic [0:0] f542_wen;
  logic [31:0] f542_wdata;
  logic [0:0] f542_clk;
  logic [0:0] f542_rst;
  logic [31:0] f542_rdata;
  sr_buffer_32_1 f542(.wen(f542_wen), .wdata(f542_wdata), .clk(f542_clk), .rst(f542_rst), .rdata(f542_rdata));
  assign f542_clk = clk;
  assign f542_rst = rst;
  // Bindings to f542

  // f544
  logic [0:0] f544_wen;
  logic [31:0] f544_wdata;
  logic [0:0] f544_clk;
  logic [0:0] f544_rst;
  logic [31:0] f544_rdata;
  sr_buffer_32_1 f544(.wen(f544_wen), .wdata(f544_wdata), .clk(f544_clk), .rst(f544_rst), .rdata(f544_rdata));
  assign f544_clk = clk;
  assign f544_rst = rst;
  // Bindings to f544

  // f546
  logic [0:0] f546_wen;
  logic [31:0] f546_wdata;
  logic [0:0] f546_clk;
  logic [0:0] f546_rst;
  logic [31:0] f546_rdata;
  sr_buffer_32_1 f546(.wen(f546_wen), .wdata(f546_wdata), .clk(f546_clk), .rst(f546_rst), .rdata(f546_rdata));
  assign f546_clk = clk;
  assign f546_rst = rst;
  // Bindings to f546

  // f548
  logic [0:0] f548_wen;
  logic [31:0] f548_wdata;
  logic [0:0] f548_clk;
  logic [0:0] f548_rst;
  logic [31:0] f548_rdata;
  sr_buffer_32_1 f548(.wen(f548_wen), .wdata(f548_wdata), .clk(f548_clk), .rst(f548_rst), .rdata(f548_rdata));
  assign f548_clk = clk;
  assign f548_rst = rst;
  // Bindings to f548

  // f550
  logic [0:0] f550_wen;
  logic [31:0] f550_wdata;
  logic [0:0] f550_clk;
  logic [0:0] f550_rst;
  logic [31:0] f550_rdata;
  sr_buffer_32_1 f550(.wen(f550_wen), .wdata(f550_wdata), .clk(f550_clk), .rst(f550_rst), .rdata(f550_rdata));
  assign f550_clk = clk;
  assign f550_rst = rst;
  // Bindings to f550

  // f552
  logic [0:0] f552_wen;
  logic [31:0] f552_wdata;
  logic [0:0] f552_clk;
  logic [0:0] f552_rst;
  logic [31:0] f552_rdata;
  sr_buffer_32_1 f552(.wen(f552_wen), .wdata(f552_wdata), .clk(f552_clk), .rst(f552_rst), .rdata(f552_rdata));
  assign f552_clk = clk;
  assign f552_rst = rst;
  // Bindings to f552

  // f554
  logic [0:0] f554_wen;
  logic [31:0] f554_wdata;
  logic [0:0] f554_clk;
  logic [0:0] f554_rst;
  logic [31:0] f554_rdata;
  sr_buffer_32_1 f554(.wen(f554_wen), .wdata(f554_wdata), .clk(f554_clk), .rst(f554_rst), .rdata(f554_rdata));
  assign f554_clk = clk;
  assign f554_rst = rst;
  // Bindings to f554

  // f556
  logic [0:0] f556_wen;
  logic [31:0] f556_wdata;
  logic [0:0] f556_clk;
  logic [0:0] f556_rst;
  logic [31:0] f556_rdata;
  sr_buffer_32_1 f556(.wen(f556_wen), .wdata(f556_wdata), .clk(f556_clk), .rst(f556_rst), .rdata(f556_rdata));
  assign f556_clk = clk;
  assign f556_rst = rst;
  // Bindings to f556

  // f558
  logic [0:0] f558_wen;
  logic [31:0] f558_wdata;
  logic [0:0] f558_clk;
  logic [0:0] f558_rst;
  logic [31:0] f558_rdata;
  sr_buffer_32_1 f558(.wen(f558_wen), .wdata(f558_wdata), .clk(f558_clk), .rst(f558_rst), .rdata(f558_rdata));
  assign f558_clk = clk;
  assign f558_rst = rst;
  // Bindings to f558

  // f560
  logic [0:0] f560_wen;
  logic [31:0] f560_wdata;
  logic [0:0] f560_clk;
  logic [0:0] f560_rst;
  logic [31:0] f560_rdata;
  sr_buffer_32_1 f560(.wen(f560_wen), .wdata(f560_wdata), .clk(f560_clk), .rst(f560_rst), .rdata(f560_rdata));
  assign f560_clk = clk;
  assign f560_rst = rst;
  // Bindings to f560

  // f562
  logic [0:0] f562_wen;
  logic [31:0] f562_wdata;
  logic [0:0] f562_clk;
  logic [0:0] f562_rst;
  logic [31:0] f562_rdata;
  sr_buffer_32_1 f562(.wen(f562_wen), .wdata(f562_wdata), .clk(f562_clk), .rst(f562_rst), .rdata(f562_rdata));
  assign f562_clk = clk;
  assign f562_rst = rst;
  // Bindings to f562

  // f564
  logic [0:0] f564_wen;
  logic [31:0] f564_wdata;
  logic [0:0] f564_clk;
  logic [0:0] f564_rst;
  logic [31:0] f564_rdata;
  sr_buffer_32_1 f564(.wen(f564_wen), .wdata(f564_wdata), .clk(f564_clk), .rst(f564_rst), .rdata(f564_rdata));
  assign f564_clk = clk;
  assign f564_rst = rst;
  // Bindings to f564

  // f566
  logic [0:0] f566_wen;
  logic [31:0] f566_wdata;
  logic [0:0] f566_clk;
  logic [0:0] f566_rst;
  logic [31:0] f566_rdata;
  sr_buffer_32_1 f566(.wen(f566_wen), .wdata(f566_wdata), .clk(f566_clk), .rst(f566_rst), .rdata(f566_rdata));
  assign f566_clk = clk;
  assign f566_rst = rst;
  // Bindings to f566

  // f568
  logic [0:0] f568_wen;
  logic [31:0] f568_wdata;
  logic [0:0] f568_clk;
  logic [0:0] f568_rst;
  logic [31:0] f568_rdata;
  sr_buffer_32_1 f568(.wen(f568_wen), .wdata(f568_wdata), .clk(f568_clk), .rst(f568_rst), .rdata(f568_rdata));
  assign f568_clk = clk;
  assign f568_rst = rst;
  // Bindings to f568

  // f570
  logic [0:0] f570_wen;
  logic [31:0] f570_wdata;
  logic [0:0] f570_clk;
  logic [0:0] f570_rst;
  logic [31:0] f570_rdata;
  sr_buffer_32_1 f570(.wen(f570_wen), .wdata(f570_wdata), .clk(f570_clk), .rst(f570_rst), .rdata(f570_rdata));
  assign f570_clk = clk;
  assign f570_rst = rst;
  // Bindings to f570

  // f572
  logic [0:0] f572_wen;
  logic [31:0] f572_wdata;
  logic [0:0] f572_clk;
  logic [0:0] f572_rst;
  logic [31:0] f572_rdata;
  sr_buffer_32_1 f572(.wen(f572_wen), .wdata(f572_wdata), .clk(f572_clk), .rst(f572_rst), .rdata(f572_rdata));
  assign f572_clk = clk;
  assign f572_rst = rst;
  // Bindings to f572

  // f574
  logic [0:0] f574_wen;
  logic [31:0] f574_wdata;
  logic [0:0] f574_clk;
  logic [0:0] f574_rst;
  logic [31:0] f574_rdata;
  sr_buffer_32_1 f574(.wen(f574_wen), .wdata(f574_wdata), .clk(f574_clk), .rst(f574_rst), .rdata(f574_rdata));
  assign f574_clk = clk;
  assign f574_rst = rst;
  // Bindings to f574

  // f576
  logic [0:0] f576_wen;
  logic [31:0] f576_wdata;
  logic [0:0] f576_clk;
  logic [0:0] f576_rst;
  logic [31:0] f576_rdata;
  sr_buffer_32_1 f576(.wen(f576_wen), .wdata(f576_wdata), .clk(f576_clk), .rst(f576_rst), .rdata(f576_rdata));
  assign f576_clk = clk;
  assign f576_rst = rst;
  // Bindings to f576

  // f578
  logic [0:0] f578_wen;
  logic [31:0] f578_wdata;
  logic [0:0] f578_clk;
  logic [0:0] f578_rst;
  logic [31:0] f578_rdata;
  sr_buffer_32_1 f578(.wen(f578_wen), .wdata(f578_wdata), .clk(f578_clk), .rst(f578_rst), .rdata(f578_rdata));
  assign f578_clk = clk;
  assign f578_rst = rst;
  // Bindings to f578

  // f580
  logic [0:0] f580_wen;
  logic [31:0] f580_wdata;
  logic [0:0] f580_clk;
  logic [0:0] f580_rst;
  logic [31:0] f580_rdata;
  sr_buffer_32_1 f580(.wen(f580_wen), .wdata(f580_wdata), .clk(f580_clk), .rst(f580_rst), .rdata(f580_rdata));
  assign f580_clk = clk;
  assign f580_rst = rst;
  // Bindings to f580

  // f582
  logic [0:0] f582_wen;
  logic [31:0] f582_wdata;
  logic [0:0] f582_clk;
  logic [0:0] f582_rst;
  logic [31:0] f582_rdata;
  sr_buffer_32_1 f582(.wen(f582_wen), .wdata(f582_wdata), .clk(f582_clk), .rst(f582_rst), .rdata(f582_rdata));
  assign f582_clk = clk;
  assign f582_rst = rst;
  // Bindings to f582

  // f584
  logic [0:0] f584_wen;
  logic [31:0] f584_wdata;
  logic [0:0] f584_clk;
  logic [0:0] f584_rst;
  logic [31:0] f584_rdata;
  sr_buffer_32_1 f584(.wen(f584_wen), .wdata(f584_wdata), .clk(f584_clk), .rst(f584_rst), .rdata(f584_rdata));
  assign f584_clk = clk;
  assign f584_rst = rst;
  // Bindings to f584

  // f586
  logic [0:0] f586_wen;
  logic [31:0] f586_wdata;
  logic [0:0] f586_clk;
  logic [0:0] f586_rst;
  logic [31:0] f586_rdata;
  sr_buffer_32_1 f586(.wen(f586_wen), .wdata(f586_wdata), .clk(f586_clk), .rst(f586_rst), .rdata(f586_rdata));
  assign f586_clk = clk;
  assign f586_rst = rst;
  // Bindings to f586

  // f588
  logic [0:0] f588_wen;
  logic [31:0] f588_wdata;
  logic [0:0] f588_clk;
  logic [0:0] f588_rst;
  logic [31:0] f588_rdata;
  sr_buffer_32_1 f588(.wen(f588_wen), .wdata(f588_wdata), .clk(f588_clk), .rst(f588_rst), .rdata(f588_rdata));
  assign f588_clk = clk;
  assign f588_rst = rst;
  // Bindings to f588

  // f590
  logic [0:0] f590_wen;
  logic [31:0] f590_wdata;
  logic [0:0] f590_clk;
  logic [0:0] f590_rst;
  logic [31:0] f590_rdata;
  sr_buffer_32_1 f590(.wen(f590_wen), .wdata(f590_wdata), .clk(f590_clk), .rst(f590_rst), .rdata(f590_rdata));
  assign f590_clk = clk;
  assign f590_rst = rst;
  // Bindings to f590

  // f592
  logic [0:0] f592_wen;
  logic [31:0] f592_wdata;
  logic [0:0] f592_clk;
  logic [0:0] f592_rst;
  logic [31:0] f592_rdata;
  sr_buffer_32_1 f592(.wen(f592_wen), .wdata(f592_wdata), .clk(f592_clk), .rst(f592_rst), .rdata(f592_rdata));
  assign f592_clk = clk;
  assign f592_rst = rst;
  // Bindings to f592

  // f594
  logic [0:0] f594_wen;
  logic [31:0] f594_wdata;
  logic [0:0] f594_clk;
  logic [0:0] f594_rst;
  logic [31:0] f594_rdata;
  sr_buffer_32_1 f594(.wen(f594_wen), .wdata(f594_wdata), .clk(f594_clk), .rst(f594_rst), .rdata(f594_rdata));
  assign f594_clk = clk;
  assign f594_rst = rst;
  // Bindings to f594

  // f596
  logic [0:0] f596_wen;
  logic [31:0] f596_wdata;
  logic [0:0] f596_clk;
  logic [0:0] f596_rst;
  logic [31:0] f596_rdata;
  sr_buffer_32_1 f596(.wen(f596_wen), .wdata(f596_wdata), .clk(f596_clk), .rst(f596_rst), .rdata(f596_rdata));
  assign f596_clk = clk;
  assign f596_rst = rst;
  // Bindings to f596

  // f598
  logic [0:0] f598_wen;
  logic [31:0] f598_wdata;
  logic [0:0] f598_clk;
  logic [0:0] f598_rst;
  logic [31:0] f598_rdata;
  sr_buffer_32_1 f598(.wen(f598_wen), .wdata(f598_wdata), .clk(f598_clk), .rst(f598_rst), .rdata(f598_rdata));
  assign f598_clk = clk;
  assign f598_rst = rst;
  // Bindings to f598

  // f600
  logic [0:0] f600_wen;
  logic [31:0] f600_wdata;
  logic [0:0] f600_clk;
  logic [0:0] f600_rst;
  logic [31:0] f600_rdata;
  sr_buffer_32_1 f600(.wen(f600_wen), .wdata(f600_wdata), .clk(f600_clk), .rst(f600_rst), .rdata(f600_rdata));
  assign f600_clk = clk;
  assign f600_rst = rst;
  // Bindings to f600

  // f602
  logic [0:0] f602_wen;
  logic [31:0] f602_wdata;
  logic [0:0] f602_clk;
  logic [0:0] f602_rst;
  logic [31:0] f602_rdata;
  sr_buffer_32_1 f602(.wen(f602_wen), .wdata(f602_wdata), .clk(f602_clk), .rst(f602_rst), .rdata(f602_rdata));
  assign f602_clk = clk;
  assign f602_rst = rst;
  // Bindings to f602

  // f604
  logic [0:0] f604_wen;
  logic [31:0] f604_wdata;
  logic [0:0] f604_clk;
  logic [0:0] f604_rst;
  logic [31:0] f604_rdata;
  sr_buffer_32_1 f604(.wen(f604_wen), .wdata(f604_wdata), .clk(f604_clk), .rst(f604_rst), .rdata(f604_rdata));
  assign f604_clk = clk;
  assign f604_rst = rst;
  // Bindings to f604

  // f606
  logic [0:0] f606_wen;
  logic [31:0] f606_wdata;
  logic [0:0] f606_clk;
  logic [0:0] f606_rst;
  logic [31:0] f606_rdata;
  sr_buffer_32_1 f606(.wen(f606_wen), .wdata(f606_wdata), .clk(f606_clk), .rst(f606_rst), .rdata(f606_rdata));
  assign f606_clk = clk;
  assign f606_rst = rst;
  // Bindings to f606

  // f608
  logic [0:0] f608_wen;
  logic [31:0] f608_wdata;
  logic [0:0] f608_clk;
  logic [0:0] f608_rst;
  logic [31:0] f608_rdata;
  sr_buffer_32_1 f608(.wen(f608_wen), .wdata(f608_wdata), .clk(f608_clk), .rst(f608_rst), .rdata(f608_rdata));
  assign f608_clk = clk;
  assign f608_rst = rst;
  // Bindings to f608

  // f610
  logic [0:0] f610_wen;
  logic [31:0] f610_wdata;
  logic [0:0] f610_clk;
  logic [0:0] f610_rst;
  logic [31:0] f610_rdata;
  sr_buffer_32_1 f610(.wen(f610_wen), .wdata(f610_wdata), .clk(f610_clk), .rst(f610_rst), .rdata(f610_rdata));
  assign f610_clk = clk;
  assign f610_rst = rst;
  // Bindings to f610

  // f612
  logic [0:0] f612_wen;
  logic [31:0] f612_wdata;
  logic [0:0] f612_clk;
  logic [0:0] f612_rst;
  logic [31:0] f612_rdata;
  sr_buffer_32_1 f612(.wen(f612_wen), .wdata(f612_wdata), .clk(f612_clk), .rst(f612_rst), .rdata(f612_rdata));
  assign f612_clk = clk;
  assign f612_rst = rst;
  // Bindings to f612

  // f614
  logic [0:0] f614_wen;
  logic [31:0] f614_wdata;
  logic [0:0] f614_clk;
  logic [0:0] f614_rst;
  logic [31:0] f614_rdata;
  sr_buffer_32_1 f614(.wen(f614_wen), .wdata(f614_wdata), .clk(f614_clk), .rst(f614_rst), .rdata(f614_rdata));
  assign f614_clk = clk;
  assign f614_rst = rst;
  // Bindings to f614

  // f616
  logic [0:0] f616_wen;
  logic [31:0] f616_wdata;
  logic [0:0] f616_clk;
  logic [0:0] f616_rst;
  logic [31:0] f616_rdata;
  sr_buffer_32_1 f616(.wen(f616_wen), .wdata(f616_wdata), .clk(f616_clk), .rst(f616_rst), .rdata(f616_rdata));
  assign f616_clk = clk;
  assign f616_rst = rst;
  // Bindings to f616

  // f618
  logic [0:0] f618_wen;
  logic [31:0] f618_wdata;
  logic [0:0] f618_clk;
  logic [0:0] f618_rst;
  logic [31:0] f618_rdata;
  sr_buffer_32_1 f618(.wen(f618_wen), .wdata(f618_wdata), .clk(f618_clk), .rst(f618_rst), .rdata(f618_rdata));
  assign f618_clk = clk;
  assign f618_rst = rst;
  // Bindings to f618

  // f620
  logic [0:0] f620_wen;
  logic [31:0] f620_wdata;
  logic [0:0] f620_clk;
  logic [0:0] f620_rst;
  logic [31:0] f620_rdata;
  sr_buffer_32_1 f620(.wen(f620_wen), .wdata(f620_wdata), .clk(f620_clk), .rst(f620_rst), .rdata(f620_rdata));
  assign f620_clk = clk;
  assign f620_rst = rst;
  // Bindings to f620

  // f622
  logic [0:0] f622_wen;
  logic [31:0] f622_wdata;
  logic [0:0] f622_clk;
  logic [0:0] f622_rst;
  logic [31:0] f622_rdata;
  sr_buffer_32_1 f622(.wen(f622_wen), .wdata(f622_wdata), .clk(f622_clk), .rst(f622_rst), .rdata(f622_rdata));
  assign f622_clk = clk;
  assign f622_rst = rst;
  // Bindings to f622

  // f624
  logic [0:0] f624_wen;
  logic [31:0] f624_wdata;
  logic [0:0] f624_clk;
  logic [0:0] f624_rst;
  logic [31:0] f624_rdata;
  sr_buffer_32_1 f624(.wen(f624_wen), .wdata(f624_wdata), .clk(f624_clk), .rst(f624_rst), .rdata(f624_rdata));
  assign f624_clk = clk;
  assign f624_rst = rst;
  // Bindings to f624

  // f626
  logic [0:0] f626_wen;
  logic [31:0] f626_wdata;
  logic [0:0] f626_clk;
  logic [0:0] f626_rst;
  logic [31:0] f626_rdata;
  sr_buffer_32_1 f626(.wen(f626_wen), .wdata(f626_wdata), .clk(f626_clk), .rst(f626_rst), .rdata(f626_rdata));
  assign f626_clk = clk;
  assign f626_rst = rst;
  // Bindings to f626



endmodule


module bright_gauss_blur_3_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module bright_gauss_blur_3_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 631;
    end
  end

endmodule


module bright_gauss_blur_3_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 316;
    end
  end

endmodule


module bright_gauss_blur_3_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module bright_gauss_blur_3_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_gauss_ds_2_update_0_write_wen(output [0:0] bright_gauss_ds_2_update_0_write_wen);

endmodule


module bright_laplace_us_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (-1 + d1 == 0) ? ((944 - floord(d0, 2))) : (d1 == 0) ? (632) : ((-1 - d1) % 2 == 0 && -3 + d1 >= 0) ? ((944 - floord(d0, 2))) : ((-d1) % 2 == 0 && -2 + d1 >= 0) ? (632) : 0;
    end
  end

endmodule


module bright_gauss_blur_3_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (311 - d0 >= 0) ? (315) : (-312 + d0 == 0) ? (315) : 0;
    end
  end

endmodule


module in_wire_bright_gauss_ds_2_update_0_write_wdata(output [31:0] bright_gauss_ds_2_update_0_write_wdata);

endmodule


module bright_gauss_ds_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [287:0] bright_gauss_blur_3_update_0_read_dummy, output [31:0] bright_laplace_us_1_update_0_read_rdata, input [31:0] bright_laplace_us_1_update_0_read_dummy, output [31:0] bright_laplace_diff_2_update_0_read_rdata, input [31:0] bright_laplace_diff_2_update_0_read_dummy, output [287:0] bright_gauss_blur_3_update_0_read_rdata, input [0:0] bright_gauss_ds_2_update_0_write_wen, input [31:0] bright_gauss_ds_2_update_0_write_wdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;
  logic [31:0] rd_6;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;
  reg [31:0] rd_6_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;
      rd_6_stage_1 <= rd_6;


    end

  end


  // Data processing units...
  // bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_clk;
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_rst;
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_start;
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_done;
  bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10 bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10(.clk(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_clk), .rst(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_rst), .start(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_start), .done(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_done));
  assign bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_clk = clk;
  assign bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_merged_banks_10

  // Bindings to bright_gauss_blur_3_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_gauss_blur_3_update_0_read_dummy;

  // selector_bright_gauss_blur_3_rd2_select
  logic [0:0] selector_bright_gauss_blur_3_rd2_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd2_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd2_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd2_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd2_select_out;
  bright_gauss_blur_3_rd2_select selector_bright_gauss_blur_3_rd2_select(.clk(selector_bright_gauss_blur_3_rd2_select_clk), .rst(selector_bright_gauss_blur_3_rd2_select_rst), .d0(selector_bright_gauss_blur_3_rd2_select_d0), .d1(selector_bright_gauss_blur_3_rd2_select_d1), .out(selector_bright_gauss_blur_3_rd2_select_out));
  assign selector_bright_gauss_blur_3_rd2_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd2_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd2_select

  // selector_bright_gauss_blur_3_rd0_select
  logic [0:0] selector_bright_gauss_blur_3_rd0_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd0_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd0_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd0_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd0_select_out;
  bright_gauss_blur_3_rd0_select selector_bright_gauss_blur_3_rd0_select(.clk(selector_bright_gauss_blur_3_rd0_select_clk), .rst(selector_bright_gauss_blur_3_rd0_select_rst), .d0(selector_bright_gauss_blur_3_rd0_select_d0), .d1(selector_bright_gauss_blur_3_rd0_select_d1), .out(selector_bright_gauss_blur_3_rd0_select_out));
  assign selector_bright_gauss_blur_3_rd0_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd0_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd0_select

  // selector_bright_gauss_blur_3_rd1_select
  logic [0:0] selector_bright_gauss_blur_3_rd1_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd1_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd1_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd1_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd1_select_out;
  bright_gauss_blur_3_rd1_select selector_bright_gauss_blur_3_rd1_select(.clk(selector_bright_gauss_blur_3_rd1_select_clk), .rst(selector_bright_gauss_blur_3_rd1_select_rst), .d0(selector_bright_gauss_blur_3_rd1_select_d0), .d1(selector_bright_gauss_blur_3_rd1_select_d1), .out(selector_bright_gauss_blur_3_rd1_select_out));
  assign selector_bright_gauss_blur_3_rd1_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd1_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd1_select

  // Bindings to bright_laplace_us_1_update_0_read_rdata
    // wr_7
  assign bright_laplace_us_1_update_0_read_rdata = rd_6;

  // Bindings to bright_laplace_us_1_update_0_read_dummy
    // rd_6
  assign rd_6 = bright_laplace_us_1_update_0_read_dummy;

  // Bindings to bright_laplace_diff_2_update_0_read_rdata
    // wr_5
  assign bright_laplace_diff_2_update_0_read_rdata = rd_4;

  // Bindings to bright_laplace_diff_2_update_0_read_dummy
    // rd_4
  assign rd_4 = bright_laplace_diff_2_update_0_read_dummy;

  // Bindings to bright_gauss_blur_3_update_0_read_rdata
    // wr_3
  assign bright_gauss_blur_3_update_0_read_rdata = rd_2;

  // selector_bright_laplace_us_1_rd0_select
  logic [0:0] selector_bright_laplace_us_1_rd0_select_clk;
  logic [0:0] selector_bright_laplace_us_1_rd0_select_rst;
  logic [31:0] selector_bright_laplace_us_1_rd0_select_d0;
  logic [31:0] selector_bright_laplace_us_1_rd0_select_d1;
  logic [31:0] selector_bright_laplace_us_1_rd0_select_out;
  bright_laplace_us_1_rd0_select selector_bright_laplace_us_1_rd0_select(.clk(selector_bright_laplace_us_1_rd0_select_clk), .rst(selector_bright_laplace_us_1_rd0_select_rst), .d0(selector_bright_laplace_us_1_rd0_select_d0), .d1(selector_bright_laplace_us_1_rd0_select_d1), .out(selector_bright_laplace_us_1_rd0_select_out));
  assign selector_bright_laplace_us_1_rd0_select_clk = clk;
  assign selector_bright_laplace_us_1_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_us_1_rd0_select

  // Bindings to bright_gauss_ds_2_update_0_write_wen
    // rd_0
  assign rd_0 = bright_gauss_ds_2_update_0_write_wen;

  // selector_bright_laplace_diff_2_rd0_select
  logic [0:0] selector_bright_laplace_diff_2_rd0_select_clk;
  logic [0:0] selector_bright_laplace_diff_2_rd0_select_rst;
  logic [31:0] selector_bright_laplace_diff_2_rd0_select_d0;
  logic [31:0] selector_bright_laplace_diff_2_rd0_select_d1;
  logic [31:0] selector_bright_laplace_diff_2_rd0_select_out;
  bright_laplace_diff_2_rd0_select selector_bright_laplace_diff_2_rd0_select(.clk(selector_bright_laplace_diff_2_rd0_select_clk), .rst(selector_bright_laplace_diff_2_rd0_select_rst), .d0(selector_bright_laplace_diff_2_rd0_select_d0), .d1(selector_bright_laplace_diff_2_rd0_select_d1), .out(selector_bright_laplace_diff_2_rd0_select_out));
  assign selector_bright_laplace_diff_2_rd0_select_clk = clk;
  assign selector_bright_laplace_diff_2_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_diff_2_rd0_select

  // selector_bright_gauss_blur_3_rd8_select
  logic [0:0] selector_bright_gauss_blur_3_rd8_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd8_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd8_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd8_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd8_select_out;
  bright_gauss_blur_3_rd8_select selector_bright_gauss_blur_3_rd8_select(.clk(selector_bright_gauss_blur_3_rd8_select_clk), .rst(selector_bright_gauss_blur_3_rd8_select_rst), .d0(selector_bright_gauss_blur_3_rd8_select_d0), .d1(selector_bright_gauss_blur_3_rd8_select_d1), .out(selector_bright_gauss_blur_3_rd8_select_out));
  assign selector_bright_gauss_blur_3_rd8_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd8_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd8_select

  // selector_bright_gauss_blur_3_rd7_select
  logic [0:0] selector_bright_gauss_blur_3_rd7_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd7_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd7_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd7_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd7_select_out;
  bright_gauss_blur_3_rd7_select selector_bright_gauss_blur_3_rd7_select(.clk(selector_bright_gauss_blur_3_rd7_select_clk), .rst(selector_bright_gauss_blur_3_rd7_select_rst), .d0(selector_bright_gauss_blur_3_rd7_select_d0), .d1(selector_bright_gauss_blur_3_rd7_select_d1), .out(selector_bright_gauss_blur_3_rd7_select_out));
  assign selector_bright_gauss_blur_3_rd7_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd7_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd7_select

  // selector_bright_gauss_blur_3_rd5_select
  logic [0:0] selector_bright_gauss_blur_3_rd5_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd5_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd5_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd5_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd5_select_out;
  bright_gauss_blur_3_rd5_select selector_bright_gauss_blur_3_rd5_select(.clk(selector_bright_gauss_blur_3_rd5_select_clk), .rst(selector_bright_gauss_blur_3_rd5_select_rst), .d0(selector_bright_gauss_blur_3_rd5_select_d0), .d1(selector_bright_gauss_blur_3_rd5_select_d1), .out(selector_bright_gauss_blur_3_rd5_select_out));
  assign selector_bright_gauss_blur_3_rd5_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd5_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd5_select

  // selector_bright_gauss_blur_3_rd6_select
  logic [0:0] selector_bright_gauss_blur_3_rd6_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd6_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd6_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd6_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd6_select_out;
  bright_gauss_blur_3_rd6_select selector_bright_gauss_blur_3_rd6_select(.clk(selector_bright_gauss_blur_3_rd6_select_clk), .rst(selector_bright_gauss_blur_3_rd6_select_rst), .d0(selector_bright_gauss_blur_3_rd6_select_d0), .d1(selector_bright_gauss_blur_3_rd6_select_d1), .out(selector_bright_gauss_blur_3_rd6_select_out));
  assign selector_bright_gauss_blur_3_rd6_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd6_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd6_select

  // selector_bright_gauss_blur_3_rd4_select
  logic [0:0] selector_bright_gauss_blur_3_rd4_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd4_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd4_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd4_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd4_select_out;
  bright_gauss_blur_3_rd4_select selector_bright_gauss_blur_3_rd4_select(.clk(selector_bright_gauss_blur_3_rd4_select_clk), .rst(selector_bright_gauss_blur_3_rd4_select_rst), .d0(selector_bright_gauss_blur_3_rd4_select_d0), .d1(selector_bright_gauss_blur_3_rd4_select_d1), .out(selector_bright_gauss_blur_3_rd4_select_out));
  assign selector_bright_gauss_blur_3_rd4_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd4_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd4_select

  // selector_bright_gauss_blur_3_rd3_select
  logic [0:0] selector_bright_gauss_blur_3_rd3_select_clk;
  logic [0:0] selector_bright_gauss_blur_3_rd3_select_rst;
  logic [31:0] selector_bright_gauss_blur_3_rd3_select_d0;
  logic [31:0] selector_bright_gauss_blur_3_rd3_select_d1;
  logic [31:0] selector_bright_gauss_blur_3_rd3_select_out;
  bright_gauss_blur_3_rd3_select selector_bright_gauss_blur_3_rd3_select(.clk(selector_bright_gauss_blur_3_rd3_select_clk), .rst(selector_bright_gauss_blur_3_rd3_select_rst), .d0(selector_bright_gauss_blur_3_rd3_select_d0), .d1(selector_bright_gauss_blur_3_rd3_select_d1), .out(selector_bright_gauss_blur_3_rd3_select_out));
  assign selector_bright_gauss_blur_3_rd3_select_clk = clk;
  assign selector_bright_gauss_blur_3_rd3_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_3_rd3_select

  // bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_clk;
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_rst;
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_start;
  logic [0:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_done;
  bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0 bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0(.clk(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_clk), .rst(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_rst), .start(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_start), .done(bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_done));
  assign bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_clk = clk;
  assign bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0_rst = rst;
  // Bindings to bright_gauss_ds_2_bright_gauss_ds_2_update_0_write0_to_bright_laplace_us_1_rd0

  // Bindings to bright_gauss_ds_2_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_gauss_ds_2_update_0_write_wdata;



endmodule


module in_wire_bright_gauss_blur_3_update_0_read_dummy(output [287:0] bright_gauss_blur_3_update_0_read_dummy);

endmodule


module out_wire_bright_gauss_blur_3_update_0_read_rdata(input [287:0] bright_gauss_blur_3_update_0_read_rdata);

endmodule


module in_wire_bright_laplace_diff_2_update_0_read_dummy(output [31:0] bright_laplace_diff_2_update_0_read_dummy);

endmodule


module out_wire_bright_laplace_diff_2_update_0_read_rdata(input [31:0] bright_laplace_diff_2_update_0_read_rdata);

endmodule


module in_wire_bright_laplace_us_1_update_0_read_dummy(output [31:0] bright_laplace_us_1_update_0_read_dummy);

endmodule


module out_wire_bright_laplace_us_1_update_0_read_rdata(input [31:0] bright_laplace_us_1_update_0_read_rdata);

endmodule


module bright_laplace_diff_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] fused_level_0_update_0_read_rdata, input [31:0] bright_laplace_diff_0_update_0_write_wdata, input [0:0] bright_laplace_diff_0_update_0_write_wen, input [31:0] fused_level_0_update_0_read_dummy);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to fused_level_0_update_0_read_rdata
    // wr_3
  assign fused_level_0_update_0_read_rdata = rd_2;

  // Bindings to bright_laplace_diff_0_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_laplace_diff_0_update_0_write_wdata;

  // Bindings to bright_laplace_diff_0_update_0_write_wen
    // rd_0
  assign rd_0 = bright_laplace_diff_0_update_0_write_wen;

  // bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1
  logic [0:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_done;
  bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1 bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1(.clk(bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_clk), .rst(bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_rst), .start(bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_start), .done(bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_done));
  assign bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_clk = clk;
  assign bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1

  // selector_fused_level_0_rd0_select
  logic [0:0] selector_fused_level_0_rd0_select_clk;
  logic [0:0] selector_fused_level_0_rd0_select_rst;
  logic [31:0] selector_fused_level_0_rd0_select_d0;
  logic [31:0] selector_fused_level_0_rd0_select_d1;
  logic [31:0] selector_fused_level_0_rd0_select_out;
  fused_level_0_rd0_select selector_fused_level_0_rd0_select(.clk(selector_fused_level_0_rd0_select_clk), .rst(selector_fused_level_0_rd0_select_rst), .d0(selector_fused_level_0_rd0_select_d0), .d1(selector_fused_level_0_rd0_select_d1), .out(selector_fused_level_0_rd0_select_out));
  assign selector_fused_level_0_rd0_select_clk = clk;
  assign selector_fused_level_0_rd0_select_rst = rst;
  // Bindings to selector_fused_level_0_rd0_select

  // Bindings to fused_level_0_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_0_update_0_read_dummy;



endmodule


module in_wire_bright_laplace_diff_1_update_0_write_wdata(output [31:0] bright_laplace_diff_1_update_0_write_wdata);

endmodule


module bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_laplace_diff_1_update_0_write_wen(output [0:0] bright_laplace_diff_1_update_0_write_wen);

endmodule


module in_wire_fused_level_1_update_0_read_dummy(output [31:0] fused_level_1_update_0_read_dummy);

endmodule


module out_wire_fused_level_1_update_0_read_rdata(input [31:0] fused_level_1_update_0_read_rdata);

endmodule


module bright_laplace_diff_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] bright_laplace_diff_1_update_0_write_wdata, output [31:0] fused_level_1_update_0_read_rdata, input [0:0] bright_laplace_diff_1_update_0_write_wen, input [31:0] fused_level_1_update_0_read_dummy);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1
  logic [0:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_done;
  bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1 bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1(.clk(bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_clk), .rst(bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_rst), .start(bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_start), .done(bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_done));
  assign bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_clk = clk;
  assign bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_laplace_diff_1_bright_laplace_diff_1_update_0_write0_merged_banks_1

  // Bindings to bright_laplace_diff_1_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_laplace_diff_1_update_0_write_wdata;

  // Bindings to fused_level_1_update_0_read_rdata
    // wr_3
  assign fused_level_1_update_0_read_rdata = rd_2;

  // Bindings to bright_laplace_diff_1_update_0_write_wen
    // rd_0
  assign rd_0 = bright_laplace_diff_1_update_0_write_wen;

  // selector_fused_level_1_rd0_select
  logic [0:0] selector_fused_level_1_rd0_select_clk;
  logic [0:0] selector_fused_level_1_rd0_select_rst;
  logic [31:0] selector_fused_level_1_rd0_select_d0;
  logic [31:0] selector_fused_level_1_rd0_select_d1;
  logic [31:0] selector_fused_level_1_rd0_select_out;
  fused_level_1_rd0_select selector_fused_level_1_rd0_select(.clk(selector_fused_level_1_rd0_select_clk), .rst(selector_fused_level_1_rd0_select_rst), .d0(selector_fused_level_1_rd0_select_d0), .d1(selector_fused_level_1_rd0_select_d1), .out(selector_fused_level_1_rd0_select_out));
  assign selector_fused_level_1_rd0_select_clk = clk;
  assign selector_fused_level_1_rd0_select_rst = rst;
  // Bindings to selector_fused_level_1_rd0_select

  // Bindings to fused_level_1_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_1_update_0_read_dummy;



endmodule


module in_wire_bright_laplace_diff_2_update_0_write_wen(output [0:0] bright_laplace_diff_2_update_0_write_wen);

endmodule


module in_wire_bright_laplace_diff_2_update_0_write_wdata(output [31:0] bright_laplace_diff_2_update_0_write_wdata);

endmodule


module bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_fused_level_2_update_0_read_dummy(output [31:0] fused_level_2_update_0_read_dummy);

endmodule


module out_wire_fused_level_2_update_0_read_rdata(input [31:0] fused_level_2_update_0_read_rdata);

endmodule


module in_wire_bright_laplace_us_0_update_0_write_wen(output [0:0] bright_laplace_us_0_update_0_write_wen);

endmodule


module bright_laplace_diff_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_laplace_diff_2_update_0_write_wen, input [31:0] fused_level_2_update_0_read_dummy, input [31:0] bright_laplace_diff_2_update_0_write_wdata, output [31:0] fused_level_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to bright_laplace_diff_2_update_0_write_wen
    // rd_0
  assign rd_0 = bright_laplace_diff_2_update_0_write_wen;

  // Bindings to fused_level_2_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_2_update_0_read_dummy;

  // selector_fused_level_2_rd0_select
  logic [0:0] selector_fused_level_2_rd0_select_clk;
  logic [0:0] selector_fused_level_2_rd0_select_rst;
  logic [31:0] selector_fused_level_2_rd0_select_d0;
  logic [31:0] selector_fused_level_2_rd0_select_d1;
  logic [31:0] selector_fused_level_2_rd0_select_out;
  fused_level_2_rd0_select selector_fused_level_2_rd0_select(.clk(selector_fused_level_2_rd0_select_clk), .rst(selector_fused_level_2_rd0_select_rst), .d0(selector_fused_level_2_rd0_select_d0), .d1(selector_fused_level_2_rd0_select_d1), .out(selector_fused_level_2_rd0_select_out));
  assign selector_fused_level_2_rd0_select_clk = clk;
  assign selector_fused_level_2_rd0_select_rst = rst;
  // Bindings to selector_fused_level_2_rd0_select

  // Bindings to bright_laplace_diff_2_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_laplace_diff_2_update_0_write_wdata;

  // bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1
  logic [0:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_done;
  bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1 bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1(.clk(bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_clk), .rst(bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_rst), .start(bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_start), .done(bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_done));
  assign bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_clk = clk;
  assign bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_laplace_diff_2_bright_laplace_diff_2_update_0_write0_merged_banks_1

  // Bindings to fused_level_2_update_0_read_rdata
    // wr_3
  assign fused_level_2_update_0_read_rdata = rd_2;



endmodule


module bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module bright_laplace_diff_0_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_laplace_us_0_update_0_write_wdata(output [31:0] bright_laplace_us_0_update_0_write_wdata);

endmodule


module in_wire_bright_laplace_us_1_update_0_write_wen(output [0:0] bright_laplace_us_1_update_0_write_wen);

endmodule


module bright_laplace_us_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_laplace_us_0_update_0_write_wen, input [31:0] bright_laplace_us_0_update_0_write_wdata, input [31:0] bright_laplace_diff_0_update_0_read_dummy, output [31:0] bright_laplace_diff_0_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to bright_laplace_us_0_update_0_write_wen
    // rd_0
  assign rd_0 = bright_laplace_us_0_update_0_write_wen;

  // bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1
  logic [0:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_done;
  bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1 bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1(.clk(bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_clk), .rst(bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_rst), .start(bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_start), .done(bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_done));
  assign bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_clk = clk;
  assign bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_laplace_us_0_bright_laplace_us_0_update_0_write0_merged_banks_1

  // selector_bright_laplace_diff_0_rd0_select
  logic [0:0] selector_bright_laplace_diff_0_rd0_select_clk;
  logic [0:0] selector_bright_laplace_diff_0_rd0_select_rst;
  logic [31:0] selector_bright_laplace_diff_0_rd0_select_d0;
  logic [31:0] selector_bright_laplace_diff_0_rd0_select_d1;
  logic [31:0] selector_bright_laplace_diff_0_rd0_select_out;
  bright_laplace_diff_0_rd0_select selector_bright_laplace_diff_0_rd0_select(.clk(selector_bright_laplace_diff_0_rd0_select_clk), .rst(selector_bright_laplace_diff_0_rd0_select_rst), .d0(selector_bright_laplace_diff_0_rd0_select_d0), .d1(selector_bright_laplace_diff_0_rd0_select_d1), .out(selector_bright_laplace_diff_0_rd0_select_out));
  assign selector_bright_laplace_diff_0_rd0_select_clk = clk;
  assign selector_bright_laplace_diff_0_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_diff_0_rd0_select

  // Bindings to bright_laplace_us_0_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_laplace_us_0_update_0_write_wdata;

  // Bindings to bright_laplace_diff_0_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_laplace_diff_0_update_0_read_dummy;

  // Bindings to bright_laplace_diff_0_update_0_read_rdata
    // wr_3
  assign bright_laplace_diff_0_update_0_read_rdata = rd_2;



endmodule


module in_wire_bright_laplace_us_1_update_0_write_wdata(output [31:0] bright_laplace_us_1_update_0_write_wdata);

endmodule


module bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module bright_laplace_diff_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_laplace_us_2_update_0_write_wen(output [0:0] bright_laplace_us_2_update_0_write_wen);

endmodule


module bright_laplace_diff_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module bright_laplace_us_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_laplace_us_1_update_0_write_wen, input [31:0] bright_laplace_us_1_update_0_write_wdata, input [31:0] bright_laplace_diff_1_update_0_read_dummy, output [31:0] bright_laplace_diff_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1
  logic [0:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_done;
  bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1 bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1(.clk(bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_clk), .rst(bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_rst), .start(bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_start), .done(bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_done));
  assign bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_clk = clk;
  assign bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_laplace_us_1_bright_laplace_us_1_update_0_write0_merged_banks_1

  // Bindings to bright_laplace_us_1_update_0_write_wen
    // rd_0
  assign rd_0 = bright_laplace_us_1_update_0_write_wen;

  // selector_bright_laplace_diff_1_rd0_select
  logic [0:0] selector_bright_laplace_diff_1_rd0_select_clk;
  logic [0:0] selector_bright_laplace_diff_1_rd0_select_rst;
  logic [31:0] selector_bright_laplace_diff_1_rd0_select_d0;
  logic [31:0] selector_bright_laplace_diff_1_rd0_select_d1;
  logic [31:0] selector_bright_laplace_diff_1_rd0_select_out;
  bright_laplace_diff_1_rd0_select selector_bright_laplace_diff_1_rd0_select(.clk(selector_bright_laplace_diff_1_rd0_select_clk), .rst(selector_bright_laplace_diff_1_rd0_select_rst), .d0(selector_bright_laplace_diff_1_rd0_select_d0), .d1(selector_bright_laplace_diff_1_rd0_select_d1), .out(selector_bright_laplace_diff_1_rd0_select_out));
  assign selector_bright_laplace_diff_1_rd0_select_clk = clk;
  assign selector_bright_laplace_diff_1_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_diff_1_rd0_select

  // Bindings to bright_laplace_us_1_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_laplace_us_1_update_0_write_wdata;

  // Bindings to bright_laplace_diff_1_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_laplace_diff_1_update_0_read_dummy;

  // Bindings to bright_laplace_diff_1_update_0_read_rdata
    // wr_3
  assign bright_laplace_diff_1_update_0_read_rdata = rd_2;



endmodule


module in_wire_bright_laplace_us_2_update_0_write_wdata(output [31:0] bright_laplace_us_2_update_0_write_wdata);

endmodule


module bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module bright_laplace_us_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_laplace_us_2_update_0_write_wen, input [31:0] bright_laplace_us_2_update_0_write_wdata, input [31:0] bright_laplace_diff_2_update_0_read_dummy, output [31:0] bright_laplace_diff_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1
  logic [0:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_done;
  bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1 bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1(.clk(bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_clk), .rst(bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_rst), .start(bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_start), .done(bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_done));
  assign bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_clk = clk;
  assign bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_laplace_us_2_bright_laplace_us_2_update_0_write0_merged_banks_1

  // Bindings to bright_laplace_us_2_update_0_write_wen
    // rd_0
  assign rd_0 = bright_laplace_us_2_update_0_write_wen;

  // Bindings to bright_laplace_us_2_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_laplace_us_2_update_0_write_wdata;

  // selector_bright_laplace_diff_2_rd0_select
  logic [0:0] selector_bright_laplace_diff_2_rd0_select_clk;
  logic [0:0] selector_bright_laplace_diff_2_rd0_select_rst;
  logic [31:0] selector_bright_laplace_diff_2_rd0_select_d0;
  logic [31:0] selector_bright_laplace_diff_2_rd0_select_d1;
  logic [31:0] selector_bright_laplace_diff_2_rd0_select_out;
  bright_laplace_diff_2_rd0_select selector_bright_laplace_diff_2_rd0_select(.clk(selector_bright_laplace_diff_2_rd0_select_clk), .rst(selector_bright_laplace_diff_2_rd0_select_rst), .d0(selector_bright_laplace_diff_2_rd0_select_d0), .d1(selector_bright_laplace_diff_2_rd0_select_d1), .out(selector_bright_laplace_diff_2_rd0_select_out));
  assign selector_bright_laplace_diff_2_rd0_select_clk = clk;
  assign selector_bright_laplace_diff_2_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_diff_2_rd0_select

  // Bindings to bright_laplace_diff_2_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_laplace_diff_2_update_0_read_dummy;

  // Bindings to bright_laplace_diff_2_update_0_read_rdata
    // wr_3
  assign bright_laplace_diff_2_update_0_read_rdata = rd_2;



endmodule


module bright_weights(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] weight_sums_update_0_read_dummy, input [0:0] bright_weights_update_0_write_wen, input [31:0] bright_weights_update_0_write_wdata, input [31:0] bright_weights_normed_update_0_read_dummy, output [31:0] bright_weights_normed_update_0_read_rdata, output [31:0] weight_sums_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // Bindings to weight_sums_update_0_read_dummy
    // rd_4
  assign rd_4 = weight_sums_update_0_read_dummy;

  // selector_weight_sums_rd0_select
  logic [0:0] selector_weight_sums_rd0_select_clk;
  logic [0:0] selector_weight_sums_rd0_select_rst;
  logic [31:0] selector_weight_sums_rd0_select_d0;
  logic [31:0] selector_weight_sums_rd0_select_d1;
  logic [31:0] selector_weight_sums_rd0_select_out;
  weight_sums_rd0_select selector_weight_sums_rd0_select(.clk(selector_weight_sums_rd0_select_clk), .rst(selector_weight_sums_rd0_select_rst), .d0(selector_weight_sums_rd0_select_d0), .d1(selector_weight_sums_rd0_select_d1), .out(selector_weight_sums_rd0_select_out));
  assign selector_weight_sums_rd0_select_clk = clk;
  assign selector_weight_sums_rd0_select_rst = rst;
  // Bindings to selector_weight_sums_rd0_select

  // Bindings to bright_weights_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_update_0_write_wen;

  // selector_bright_weights_normed_rd0_select
  logic [0:0] selector_bright_weights_normed_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_rd0_select_out;
  bright_weights_normed_rd0_select selector_bright_weights_normed_rd0_select(.clk(selector_bright_weights_normed_rd0_select_clk), .rst(selector_bright_weights_normed_rd0_select_rst), .d0(selector_bright_weights_normed_rd0_select_d0), .d1(selector_bright_weights_normed_rd0_select_d1), .out(selector_bright_weights_normed_rd0_select_out));
  assign selector_bright_weights_normed_rd0_select_clk = clk;
  assign selector_bright_weights_normed_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_rd0_select

  // Bindings to bright_weights_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_update_0_write_wdata;

  // Bindings to bright_weights_normed_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_update_0_read_dummy;

  // Bindings to bright_weights_normed_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_update_0_read_rdata = rd_2;

  // Bindings to weight_sums_update_0_read_rdata
    // wr_5
  assign weight_sums_update_0_read_rdata = rd_4;

  // bright_weights_bright_weights_update_0_write0_merged_banks_2
  logic [0:0] bright_weights_bright_weights_update_0_write0_merged_banks_2_clk;
  logic [0:0] bright_weights_bright_weights_update_0_write0_merged_banks_2_rst;
  logic [0:0] bright_weights_bright_weights_update_0_write0_merged_banks_2_start;
  logic [0:0] bright_weights_bright_weights_update_0_write0_merged_banks_2_done;
  bright_weights_bright_weights_update_0_write0_merged_banks_2 bright_weights_bright_weights_update_0_write0_merged_banks_2(.clk(bright_weights_bright_weights_update_0_write0_merged_banks_2_clk), .rst(bright_weights_bright_weights_update_0_write0_merged_banks_2_rst), .start(bright_weights_bright_weights_update_0_write0_merged_banks_2_start), .done(bright_weights_bright_weights_update_0_write0_merged_banks_2_done));
  assign bright_weights_bright_weights_update_0_write0_merged_banks_2_clk = clk;
  assign bright_weights_bright_weights_update_0_write0_merged_banks_2_rst = rst;
  // Bindings to bright_weights_bright_weights_update_0_write0_merged_banks_2



endmodule


module bright_weights_bright_weights_update_0_write0_merged_banks_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f17
  logic [0:0] f17_wen;
  logic [31:0] f17_wdata;
  logic [0:0] f17_clk;
  logic [0:0] f17_rst;
  logic [31:0] f17_rdata;
  sr_buffer_32_2527 f17(.wen(f17_wen), .wdata(f17_wdata), .clk(f17_clk), .rst(f17_rst), .rdata(f17_rdata));
  assign f17_clk = clk;
  assign f17_rst = rst;
  // Bindings to f17

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_628 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_628 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0



endmodule


module bright_weights_normed_gauss_blur_2_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (627 - d0 >= 0) ? (1262) : (-628 + d0 == 0) ? (1262) : 0;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_2_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 633;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1264;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_2_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_2_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1263;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_2_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 632;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_2_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module bright_weights_normed_gauss_blur_2_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_weights_normed_gauss_ds_1_update_0_write_wen(output [0:0] bright_weights_normed_gauss_ds_1_update_0_write_wen);

endmodule


module bright_weights_normed_gauss_blur_2_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (627 - d0 >= 0) ? (631) : (-628 + d0 == 0) ? (631) : 0;
    end
  end

endmodule


module in_wire_bright_weights_normed_gauss_ds_1_update_0_write_wdata(output [31:0] bright_weights_normed_gauss_ds_1_update_0_write_wdata);

endmodule


module in_wire_bright_weights_normed_gauss_blur_2_update_0_read_dummy(output [287:0] bright_weights_normed_gauss_blur_2_update_0_read_dummy);

endmodule


module out_wire_bright_weights_normed_gauss_blur_2_update_0_read_rdata(input [287:0] bright_weights_normed_gauss_blur_2_update_0_read_rdata);

endmodule


module bright_weights_normed_gauss_ds_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [287:0] bright_weights_normed_gauss_blur_2_update_0_read_dummy, input [31:0] bright_weights_normed_gauss_ds_1_update_0_write_wdata, input [0:0] bright_weights_normed_gauss_ds_1_update_0_write_wen, output [287:0] bright_weights_normed_gauss_blur_2_update_0_read_rdata, input [31:0] fused_level_1_update_0_read_dummy, output [31:0] fused_level_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10
  logic [0:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_clk;
  logic [0:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_rst;
  logic [0:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_start;
  logic [0:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_done;
  bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10 bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10(.clk(bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_clk), .rst(bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_rst), .start(bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_start), .done(bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_done));
  assign bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_clk = clk;
  assign bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10

  // Bindings to bright_weights_normed_gauss_blur_2_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_gauss_blur_2_update_0_read_dummy;

  // Bindings to bright_weights_normed_gauss_ds_1_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_normed_gauss_ds_1_update_0_write_wdata;

  // selector_bright_weights_normed_gauss_blur_2_rd8_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd8_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd8_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd8_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd8_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd8_select_out;
  bright_weights_normed_gauss_blur_2_rd8_select selector_bright_weights_normed_gauss_blur_2_rd8_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd8_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd8_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd8_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd8_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd8_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd8_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd8_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd8_select

  // Bindings to bright_weights_normed_gauss_ds_1_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_normed_gauss_ds_1_update_0_write_wen;

  // selector_bright_weights_normed_gauss_blur_2_rd7_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd7_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd7_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd7_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd7_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd7_select_out;
  bright_weights_normed_gauss_blur_2_rd7_select selector_bright_weights_normed_gauss_blur_2_rd7_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd7_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd7_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd7_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd7_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd7_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd7_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd7_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd7_select

  // selector_bright_weights_normed_gauss_blur_2_rd6_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd6_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd6_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd6_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd6_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd6_select_out;
  bright_weights_normed_gauss_blur_2_rd6_select selector_bright_weights_normed_gauss_blur_2_rd6_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd6_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd6_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd6_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd6_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd6_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd6_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd6_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd6_select

  // selector_bright_weights_normed_gauss_blur_2_rd5_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd5_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd5_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd5_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd5_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd5_select_out;
  bright_weights_normed_gauss_blur_2_rd5_select selector_bright_weights_normed_gauss_blur_2_rd5_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd5_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd5_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd5_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd5_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd5_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd5_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd5_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd5_select

  // selector_bright_weights_normed_gauss_blur_2_rd4_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd4_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd4_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd4_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd4_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd4_select_out;
  bright_weights_normed_gauss_blur_2_rd4_select selector_bright_weights_normed_gauss_blur_2_rd4_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd4_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd4_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd4_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd4_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd4_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd4_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd4_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd4_select

  // selector_bright_weights_normed_gauss_blur_2_rd3_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd3_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd3_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd3_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd3_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd3_select_out;
  bright_weights_normed_gauss_blur_2_rd3_select selector_bright_weights_normed_gauss_blur_2_rd3_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd3_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd3_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd3_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd3_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd3_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd3_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd3_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd3_select

  // selector_bright_weights_normed_gauss_blur_2_rd2_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd2_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd2_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd2_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd2_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd2_select_out;
  bright_weights_normed_gauss_blur_2_rd2_select selector_bright_weights_normed_gauss_blur_2_rd2_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd2_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd2_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd2_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd2_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd2_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd2_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd2_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd2_select

  // selector_bright_weights_normed_gauss_blur_2_rd0_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd0_select_out;
  bright_weights_normed_gauss_blur_2_rd0_select selector_bright_weights_normed_gauss_blur_2_rd0_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd0_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd0_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd0_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd0_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd0_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd0_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd0_select

  // selector_fused_level_1_rd0_select
  logic [0:0] selector_fused_level_1_rd0_select_clk;
  logic [0:0] selector_fused_level_1_rd0_select_rst;
  logic [31:0] selector_fused_level_1_rd0_select_d0;
  logic [31:0] selector_fused_level_1_rd0_select_d1;
  logic [31:0] selector_fused_level_1_rd0_select_out;
  fused_level_1_rd0_select selector_fused_level_1_rd0_select(.clk(selector_fused_level_1_rd0_select_clk), .rst(selector_fused_level_1_rd0_select_rst), .d0(selector_fused_level_1_rd0_select_d0), .d1(selector_fused_level_1_rd0_select_d1), .out(selector_fused_level_1_rd0_select_out));
  assign selector_fused_level_1_rd0_select_clk = clk;
  assign selector_fused_level_1_rd0_select_rst = rst;
  // Bindings to selector_fused_level_1_rd0_select

  // selector_bright_weights_normed_gauss_blur_2_rd1_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd1_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_2_rd1_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd1_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd1_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_2_rd1_select_out;
  bright_weights_normed_gauss_blur_2_rd1_select selector_bright_weights_normed_gauss_blur_2_rd1_select(.clk(selector_bright_weights_normed_gauss_blur_2_rd1_select_clk), .rst(selector_bright_weights_normed_gauss_blur_2_rd1_select_rst), .d0(selector_bright_weights_normed_gauss_blur_2_rd1_select_d0), .d1(selector_bright_weights_normed_gauss_blur_2_rd1_select_d1), .out(selector_bright_weights_normed_gauss_blur_2_rd1_select_out));
  assign selector_bright_weights_normed_gauss_blur_2_rd1_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_2_rd1_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_2_rd1_select

  // Bindings to bright_weights_normed_gauss_blur_2_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_gauss_blur_2_update_0_read_rdata = rd_2;

  // Bindings to fused_level_1_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_1_update_0_read_dummy;

  // Bindings to fused_level_1_update_0_read_rdata
    // wr_5
  assign fused_level_1_update_0_read_rdata = rd_4;



endmodule


module bright_weights_normed_gauss_ds_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [287:0] bright_weights_normed_gauss_blur_3_update_0_read_rdata, output [31:0] fused_level_2_update_0_read_rdata, input [31:0] fused_level_2_update_0_read_dummy, input [287:0] bright_weights_normed_gauss_blur_3_update_0_read_dummy, input [31:0] bright_weights_normed_gauss_ds_2_update_0_write_wdata, input [0:0] bright_weights_normed_gauss_ds_2_update_0_write_wen);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // Bindings to bright_weights_normed_gauss_blur_3_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_gauss_blur_3_update_0_read_rdata = rd_2;

  // selector_bright_weights_normed_gauss_blur_3_rd6_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd6_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd6_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd6_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd6_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd6_select_out;
  bright_weights_normed_gauss_blur_3_rd6_select selector_bright_weights_normed_gauss_blur_3_rd6_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd6_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd6_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd6_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd6_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd6_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd6_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd6_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd6_select

  // selector_bright_weights_normed_gauss_blur_3_rd0_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd0_select_out;
  bright_weights_normed_gauss_blur_3_rd0_select selector_bright_weights_normed_gauss_blur_3_rd0_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd0_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd0_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd0_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd0_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd0_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd0_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd0_select

  // Bindings to fused_level_2_update_0_read_rdata
    // wr_5
  assign fused_level_2_update_0_read_rdata = rd_4;

  // Bindings to fused_level_2_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_2_update_0_read_dummy;

  // Bindings to bright_weights_normed_gauss_blur_3_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_gauss_blur_3_update_0_read_dummy;

  // Bindings to bright_weights_normed_gauss_ds_2_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_normed_gauss_ds_2_update_0_write_wdata;

  // selector_bright_weights_normed_gauss_blur_3_rd8_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd8_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd8_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd8_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd8_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd8_select_out;
  bright_weights_normed_gauss_blur_3_rd8_select selector_bright_weights_normed_gauss_blur_3_rd8_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd8_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd8_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd8_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd8_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd8_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd8_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd8_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd8_select

  // selector_bright_weights_normed_gauss_blur_3_rd7_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd7_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd7_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd7_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd7_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd7_select_out;
  bright_weights_normed_gauss_blur_3_rd7_select selector_bright_weights_normed_gauss_blur_3_rd7_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd7_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd7_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd7_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd7_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd7_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd7_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd7_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd7_select

  // selector_bright_weights_normed_gauss_blur_3_rd5_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd5_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd5_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd5_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd5_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd5_select_out;
  bright_weights_normed_gauss_blur_3_rd5_select selector_bright_weights_normed_gauss_blur_3_rd5_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd5_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd5_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd5_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd5_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd5_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd5_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd5_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd5_select

  // selector_bright_weights_normed_gauss_blur_3_rd4_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd4_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd4_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd4_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd4_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd4_select_out;
  bright_weights_normed_gauss_blur_3_rd4_select selector_bright_weights_normed_gauss_blur_3_rd4_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd4_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd4_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd4_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd4_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd4_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd4_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd4_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd4_select

  // selector_bright_weights_normed_gauss_blur_3_rd3_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd3_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd3_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd3_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd3_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd3_select_out;
  bright_weights_normed_gauss_blur_3_rd3_select selector_bright_weights_normed_gauss_blur_3_rd3_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd3_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd3_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd3_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd3_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd3_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd3_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd3_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd3_select

  // selector_bright_weights_normed_gauss_blur_3_rd2_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd2_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd2_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd2_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd2_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd2_select_out;
  bright_weights_normed_gauss_blur_3_rd2_select selector_bright_weights_normed_gauss_blur_3_rd2_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd2_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd2_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd2_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd2_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd2_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd2_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd2_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd2_select

  // selector_bright_weights_normed_gauss_blur_3_rd1_select
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd1_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_blur_3_rd1_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd1_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd1_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_blur_3_rd1_select_out;
  bright_weights_normed_gauss_blur_3_rd1_select selector_bright_weights_normed_gauss_blur_3_rd1_select(.clk(selector_bright_weights_normed_gauss_blur_3_rd1_select_clk), .rst(selector_bright_weights_normed_gauss_blur_3_rd1_select_rst), .d0(selector_bright_weights_normed_gauss_blur_3_rd1_select_d0), .d1(selector_bright_weights_normed_gauss_blur_3_rd1_select_d1), .out(selector_bright_weights_normed_gauss_blur_3_rd1_select_out));
  assign selector_bright_weights_normed_gauss_blur_3_rd1_select_clk = clk;
  assign selector_bright_weights_normed_gauss_blur_3_rd1_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_blur_3_rd1_select

  // bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10
  logic [0:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_clk;
  logic [0:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_rst;
  logic [0:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_start;
  logic [0:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_done;
  bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10 bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10(.clk(bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_clk), .rst(bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_rst), .start(bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_start), .done(bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_done));
  assign bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_clk = clk;
  assign bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10

  // Bindings to bright_weights_normed_gauss_ds_2_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_normed_gauss_ds_2_update_0_write_wen;

  // selector_fused_level_2_rd0_select
  logic [0:0] selector_fused_level_2_rd0_select_clk;
  logic [0:0] selector_fused_level_2_rd0_select_rst;
  logic [31:0] selector_fused_level_2_rd0_select_d0;
  logic [31:0] selector_fused_level_2_rd0_select_d1;
  logic [31:0] selector_fused_level_2_rd0_select_out;
  fused_level_2_rd0_select selector_fused_level_2_rd0_select(.clk(selector_fused_level_2_rd0_select_clk), .rst(selector_fused_level_2_rd0_select_rst), .d0(selector_fused_level_2_rd0_select_d0), .d1(selector_fused_level_2_rd0_select_d1), .out(selector_fused_level_2_rd0_select_out));
  assign selector_fused_level_2_rd0_select_clk = clk;
  assign selector_fused_level_2_rd0_select_rst = rst;
  // Bindings to selector_fused_level_2_rd0_select



endmodule


module bright_weights_normed_gauss_ds_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_weights_normed_gauss_ds_3_update_0_write_wen, output [31:0] fused_level_3_update_0_read_rdata, input [31:0] bright_weights_normed_gauss_ds_3_update_0_write_wdata, input [31:0] fused_level_3_update_0_read_dummy);

  logic [31:0] rd_1;
  logic [0:0] rd_0;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_1_stage_1;
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_1_stage_1 <= rd_1;
      rd_0_stage_1 <= rd_0;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1
  logic [0:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_done;
  bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1 bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1(.clk(bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_clk), .rst(bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_rst), .start(bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_start), .done(bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_done));
  assign bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_clk = clk;
  assign bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1

  // Bindings to bright_weights_normed_gauss_ds_3_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_normed_gauss_ds_3_update_0_write_wen;

  // selector_fused_level_3_rd0_select
  logic [0:0] selector_fused_level_3_rd0_select_clk;
  logic [0:0] selector_fused_level_3_rd0_select_rst;
  logic [31:0] selector_fused_level_3_rd0_select_d0;
  logic [31:0] selector_fused_level_3_rd0_select_d1;
  logic [31:0] selector_fused_level_3_rd0_select_out;
  fused_level_3_rd0_select selector_fused_level_3_rd0_select(.clk(selector_fused_level_3_rd0_select_clk), .rst(selector_fused_level_3_rd0_select_rst), .d0(selector_fused_level_3_rd0_select_d0), .d1(selector_fused_level_3_rd0_select_d1), .out(selector_fused_level_3_rd0_select_out));
  assign selector_fused_level_3_rd0_select_clk = clk;
  assign selector_fused_level_3_rd0_select_rst = rst;
  // Bindings to selector_fused_level_3_rd0_select

  // Bindings to fused_level_3_update_0_read_rdata
    // wr_3
  assign fused_level_3_update_0_read_rdata = rd_2;

  // Bindings to bright_weights_normed_gauss_ds_3_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_normed_gauss_ds_3_update_0_write_wdata;

  // Bindings to fused_level_3_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_3_update_0_read_dummy;



endmodule


module dark_gauss_blur_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2528;
    end
  end

endmodule


module dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f388
  logic [0:0] f388_wen;
  logic [31:0] f388_wdata;
  logic [0:0] f388_clk;
  logic [0:0] f388_rst;
  logic [31:0] f388_rdata;
  sr_buffer_32_1 f388(.wen(f388_wen), .wdata(f388_wdata), .clk(f388_clk), .rst(f388_rst), .rdata(f388_rdata));
  assign f388_clk = clk;
  assign f388_rst = rst;
  // Bindings to f388

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f384
  logic [0:0] f384_wen;
  logic [31:0] f384_wdata;
  logic [0:0] f384_clk;
  logic [0:0] f384_rst;
  logic [31:0] f384_rdata;
  sr_buffer_32_1 f384(.wen(f384_wen), .wdata(f384_wdata), .clk(f384_clk), .rst(f384_rst), .rdata(f384_rdata));
  assign f384_clk = clk;
  assign f384_rst = rst;
  // Bindings to f384

  // f342
  logic [0:0] f342_wen;
  logic [31:0] f342_wdata;
  logic [0:0] f342_clk;
  logic [0:0] f342_rst;
  logic [31:0] f342_rdata;
  sr_buffer_32_1 f342(.wen(f342_wen), .wdata(f342_wdata), .clk(f342_clk), .rst(f342_rst), .rdata(f342_rdata));
  assign f342_clk = clk;
  assign f342_rst = rst;
  // Bindings to f342

  // f314
  logic [0:0] f314_wen;
  logic [31:0] f314_wdata;
  logic [0:0] f314_clk;
  logic [0:0] f314_rst;
  logic [31:0] f314_rdata;
  sr_buffer_32_1 f314(.wen(f314_wen), .wdata(f314_wdata), .clk(f314_clk), .rst(f314_rst), .rdata(f314_rdata));
  assign f314_clk = clk;
  assign f314_rst = rst;
  // Bindings to f314

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f386
  logic [0:0] f386_wen;
  logic [31:0] f386_wdata;
  logic [0:0] f386_clk;
  logic [0:0] f386_rst;
  logic [31:0] f386_rdata;
  sr_buffer_32_1 f386(.wen(f386_wen), .wdata(f386_wdata), .clk(f386_clk), .rst(f386_rst), .rdata(f386_rdata));
  assign f386_clk = clk;
  assign f386_rst = rst;
  // Bindings to f386

  // f382
  logic [0:0] f382_wen;
  logic [31:0] f382_wdata;
  logic [0:0] f382_clk;
  logic [0:0] f382_rst;
  logic [31:0] f382_rdata;
  sr_buffer_32_1 f382(.wen(f382_wen), .wdata(f382_wdata), .clk(f382_clk), .rst(f382_rst), .rdata(f382_rdata));
  assign f382_clk = clk;
  assign f382_rst = rst;
  // Bindings to f382

  // f380
  logic [0:0] f380_wen;
  logic [31:0] f380_wdata;
  logic [0:0] f380_clk;
  logic [0:0] f380_rst;
  logic [31:0] f380_rdata;
  sr_buffer_32_1 f380(.wen(f380_wen), .wdata(f380_wdata), .clk(f380_clk), .rst(f380_rst), .rdata(f380_rdata));
  assign f380_clk = clk;
  assign f380_rst = rst;
  // Bindings to f380

  // f378
  logic [0:0] f378_wen;
  logic [31:0] f378_wdata;
  logic [0:0] f378_clk;
  logic [0:0] f378_rst;
  logic [31:0] f378_rdata;
  sr_buffer_32_1 f378(.wen(f378_wen), .wdata(f378_wdata), .clk(f378_clk), .rst(f378_rst), .rdata(f378_rdata));
  assign f378_clk = clk;
  assign f378_rst = rst;
  // Bindings to f378

  // f376
  logic [0:0] f376_wen;
  logic [31:0] f376_wdata;
  logic [0:0] f376_clk;
  logic [0:0] f376_rst;
  logic [31:0] f376_rdata;
  sr_buffer_32_1 f376(.wen(f376_wen), .wdata(f376_wdata), .clk(f376_clk), .rst(f376_rst), .rdata(f376_rdata));
  assign f376_clk = clk;
  assign f376_rst = rst;
  // Bindings to f376

  // f374
  logic [0:0] f374_wen;
  logic [31:0] f374_wdata;
  logic [0:0] f374_clk;
  logic [0:0] f374_rst;
  logic [31:0] f374_rdata;
  sr_buffer_32_1 f374(.wen(f374_wen), .wdata(f374_wdata), .clk(f374_clk), .rst(f374_rst), .rdata(f374_rdata));
  assign f374_clk = clk;
  assign f374_rst = rst;
  // Bindings to f374

  // f372
  logic [0:0] f372_wen;
  logic [31:0] f372_wdata;
  logic [0:0] f372_clk;
  logic [0:0] f372_rst;
  logic [31:0] f372_rdata;
  sr_buffer_32_1 f372(.wen(f372_wen), .wdata(f372_wdata), .clk(f372_clk), .rst(f372_rst), .rdata(f372_rdata));
  assign f372_clk = clk;
  assign f372_rst = rst;
  // Bindings to f372

  // f368
  logic [0:0] f368_wen;
  logic [31:0] f368_wdata;
  logic [0:0] f368_clk;
  logic [0:0] f368_rst;
  logic [31:0] f368_rdata;
  sr_buffer_32_1 f368(.wen(f368_wen), .wdata(f368_wdata), .clk(f368_clk), .rst(f368_rst), .rdata(f368_rdata));
  assign f368_clk = clk;
  assign f368_rst = rst;
  // Bindings to f368

  // f370
  logic [0:0] f370_wen;
  logic [31:0] f370_wdata;
  logic [0:0] f370_clk;
  logic [0:0] f370_rst;
  logic [31:0] f370_rdata;
  sr_buffer_32_1 f370(.wen(f370_wen), .wdata(f370_wdata), .clk(f370_clk), .rst(f370_rst), .rdata(f370_rdata));
  assign f370_clk = clk;
  assign f370_rst = rst;
  // Bindings to f370

  // f340
  logic [0:0] f340_wen;
  logic [31:0] f340_wdata;
  logic [0:0] f340_clk;
  logic [0:0] f340_rst;
  logic [31:0] f340_rdata;
  sr_buffer_32_1 f340(.wen(f340_wen), .wdata(f340_wdata), .clk(f340_clk), .rst(f340_rst), .rdata(f340_rdata));
  assign f340_clk = clk;
  assign f340_rst = rst;
  // Bindings to f340

  // f366
  logic [0:0] f366_wen;
  logic [31:0] f366_wdata;
  logic [0:0] f366_clk;
  logic [0:0] f366_rst;
  logic [31:0] f366_rdata;
  sr_buffer_32_1 f366(.wen(f366_wen), .wdata(f366_wdata), .clk(f366_clk), .rst(f366_rst), .rdata(f366_rdata));
  assign f366_clk = clk;
  assign f366_rst = rst;
  // Bindings to f366

  // f358
  logic [0:0] f358_wen;
  logic [31:0] f358_wdata;
  logic [0:0] f358_clk;
  logic [0:0] f358_rst;
  logic [31:0] f358_rdata;
  sr_buffer_32_1 f358(.wen(f358_wen), .wdata(f358_wdata), .clk(f358_clk), .rst(f358_rst), .rdata(f358_rdata));
  assign f358_clk = clk;
  assign f358_rst = rst;
  // Bindings to f358

  // f364
  logic [0:0] f364_wen;
  logic [31:0] f364_wdata;
  logic [0:0] f364_clk;
  logic [0:0] f364_rst;
  logic [31:0] f364_rdata;
  sr_buffer_32_1 f364(.wen(f364_wen), .wdata(f364_wdata), .clk(f364_clk), .rst(f364_rst), .rdata(f364_rdata));
  assign f364_clk = clk;
  assign f364_rst = rst;
  // Bindings to f364

  // f362
  logic [0:0] f362_wen;
  logic [31:0] f362_wdata;
  logic [0:0] f362_clk;
  logic [0:0] f362_rst;
  logic [31:0] f362_rdata;
  sr_buffer_32_1 f362(.wen(f362_wen), .wdata(f362_wdata), .clk(f362_clk), .rst(f362_rst), .rdata(f362_rdata));
  assign f362_clk = clk;
  assign f362_rst = rst;
  // Bindings to f362

  // f360
  logic [0:0] f360_wen;
  logic [31:0] f360_wdata;
  logic [0:0] f360_clk;
  logic [0:0] f360_rst;
  logic [31:0] f360_rdata;
  sr_buffer_32_1 f360(.wen(f360_wen), .wdata(f360_wdata), .clk(f360_clk), .rst(f360_rst), .rdata(f360_rdata));
  assign f360_clk = clk;
  assign f360_rst = rst;
  // Bindings to f360

  // f356
  logic [0:0] f356_wen;
  logic [31:0] f356_wdata;
  logic [0:0] f356_clk;
  logic [0:0] f356_rst;
  logic [31:0] f356_rdata;
  sr_buffer_32_1 f356(.wen(f356_wen), .wdata(f356_wdata), .clk(f356_clk), .rst(f356_rst), .rdata(f356_rdata));
  assign f356_clk = clk;
  assign f356_rst = rst;
  // Bindings to f356

  // f354
  logic [0:0] f354_wen;
  logic [31:0] f354_wdata;
  logic [0:0] f354_clk;
  logic [0:0] f354_rst;
  logic [31:0] f354_rdata;
  sr_buffer_32_1 f354(.wen(f354_wen), .wdata(f354_wdata), .clk(f354_clk), .rst(f354_rst), .rdata(f354_rdata));
  assign f354_clk = clk;
  assign f354_rst = rst;
  // Bindings to f354

  // f352
  logic [0:0] f352_wen;
  logic [31:0] f352_wdata;
  logic [0:0] f352_clk;
  logic [0:0] f352_rst;
  logic [31:0] f352_rdata;
  sr_buffer_32_1 f352(.wen(f352_wen), .wdata(f352_wdata), .clk(f352_clk), .rst(f352_rst), .rdata(f352_rdata));
  assign f352_clk = clk;
  assign f352_rst = rst;
  // Bindings to f352

  // f348
  logic [0:0] f348_wen;
  logic [31:0] f348_wdata;
  logic [0:0] f348_clk;
  logic [0:0] f348_rst;
  logic [31:0] f348_rdata;
  sr_buffer_32_1 f348(.wen(f348_wen), .wdata(f348_wdata), .clk(f348_clk), .rst(f348_rst), .rdata(f348_rdata));
  assign f348_clk = clk;
  assign f348_rst = rst;
  // Bindings to f348

  // f350
  logic [0:0] f350_wen;
  logic [31:0] f350_wdata;
  logic [0:0] f350_clk;
  logic [0:0] f350_rst;
  logic [31:0] f350_rdata;
  sr_buffer_32_1 f350(.wen(f350_wen), .wdata(f350_wdata), .clk(f350_clk), .rst(f350_rst), .rdata(f350_rdata));
  assign f350_clk = clk;
  assign f350_rst = rst;
  // Bindings to f350

  // f346
  logic [0:0] f346_wen;
  logic [31:0] f346_wdata;
  logic [0:0] f346_clk;
  logic [0:0] f346_rst;
  logic [31:0] f346_rdata;
  sr_buffer_32_1 f346(.wen(f346_wen), .wdata(f346_wdata), .clk(f346_clk), .rst(f346_rst), .rdata(f346_rdata));
  assign f346_clk = clk;
  assign f346_rst = rst;
  // Bindings to f346

  // f344
  logic [0:0] f344_wen;
  logic [31:0] f344_wdata;
  logic [0:0] f344_clk;
  logic [0:0] f344_rst;
  logic [31:0] f344_rdata;
  sr_buffer_32_1 f344(.wen(f344_wen), .wdata(f344_wdata), .clk(f344_clk), .rst(f344_rst), .rdata(f344_rdata));
  assign f344_clk = clk;
  assign f344_rst = rst;
  // Bindings to f344

  // f338
  logic [0:0] f338_wen;
  logic [31:0] f338_wdata;
  logic [0:0] f338_clk;
  logic [0:0] f338_rst;
  logic [31:0] f338_rdata;
  sr_buffer_32_1 f338(.wen(f338_wen), .wdata(f338_wdata), .clk(f338_clk), .rst(f338_rst), .rdata(f338_rdata));
  assign f338_clk = clk;
  assign f338_rst = rst;
  // Bindings to f338

  // f336
  logic [0:0] f336_wen;
  logic [31:0] f336_wdata;
  logic [0:0] f336_clk;
  logic [0:0] f336_rst;
  logic [31:0] f336_rdata;
  sr_buffer_32_1 f336(.wen(f336_wen), .wdata(f336_wdata), .clk(f336_clk), .rst(f336_rst), .rdata(f336_rdata));
  assign f336_clk = clk;
  assign f336_rst = rst;
  // Bindings to f336

  // f334
  logic [0:0] f334_wen;
  logic [31:0] f334_wdata;
  logic [0:0] f334_clk;
  logic [0:0] f334_rst;
  logic [31:0] f334_rdata;
  sr_buffer_32_1 f334(.wen(f334_wen), .wdata(f334_wdata), .clk(f334_clk), .rst(f334_rst), .rdata(f334_rdata));
  assign f334_clk = clk;
  assign f334_rst = rst;
  // Bindings to f334

  // f330
  logic [0:0] f330_wen;
  logic [31:0] f330_wdata;
  logic [0:0] f330_clk;
  logic [0:0] f330_rst;
  logic [31:0] f330_rdata;
  sr_buffer_32_1 f330(.wen(f330_wen), .wdata(f330_wdata), .clk(f330_clk), .rst(f330_rst), .rdata(f330_rdata));
  assign f330_clk = clk;
  assign f330_rst = rst;
  // Bindings to f330

  // f332
  logic [0:0] f332_wen;
  logic [31:0] f332_wdata;
  logic [0:0] f332_clk;
  logic [0:0] f332_rst;
  logic [31:0] f332_rdata;
  sr_buffer_32_1 f332(.wen(f332_wen), .wdata(f332_wdata), .clk(f332_clk), .rst(f332_rst), .rdata(f332_rdata));
  assign f332_clk = clk;
  assign f332_rst = rst;
  // Bindings to f332

  // f328
  logic [0:0] f328_wen;
  logic [31:0] f328_wdata;
  logic [0:0] f328_clk;
  logic [0:0] f328_rst;
  logic [31:0] f328_rdata;
  sr_buffer_32_1 f328(.wen(f328_wen), .wdata(f328_wdata), .clk(f328_clk), .rst(f328_rst), .rdata(f328_rdata));
  assign f328_clk = clk;
  assign f328_rst = rst;
  // Bindings to f328

  // f324
  logic [0:0] f324_wen;
  logic [31:0] f324_wdata;
  logic [0:0] f324_clk;
  logic [0:0] f324_rst;
  logic [31:0] f324_rdata;
  sr_buffer_32_1 f324(.wen(f324_wen), .wdata(f324_wdata), .clk(f324_clk), .rst(f324_rst), .rdata(f324_rdata));
  assign f324_clk = clk;
  assign f324_rst = rst;
  // Bindings to f324

  // f326
  logic [0:0] f326_wen;
  logic [31:0] f326_wdata;
  logic [0:0] f326_clk;
  logic [0:0] f326_rst;
  logic [31:0] f326_rdata;
  sr_buffer_32_1 f326(.wen(f326_wen), .wdata(f326_wdata), .clk(f326_clk), .rst(f326_rst), .rdata(f326_rdata));
  assign f326_clk = clk;
  assign f326_rst = rst;
  // Bindings to f326

  // f322
  logic [0:0] f322_wen;
  logic [31:0] f322_wdata;
  logic [0:0] f322_clk;
  logic [0:0] f322_rst;
  logic [31:0] f322_rdata;
  sr_buffer_32_1 f322(.wen(f322_wen), .wdata(f322_wdata), .clk(f322_clk), .rst(f322_rst), .rdata(f322_rdata));
  assign f322_clk = clk;
  assign f322_rst = rst;
  // Bindings to f322

  // f320
  logic [0:0] f320_wen;
  logic [31:0] f320_wdata;
  logic [0:0] f320_clk;
  logic [0:0] f320_rst;
  logic [31:0] f320_rdata;
  sr_buffer_32_1 f320(.wen(f320_wen), .wdata(f320_wdata), .clk(f320_clk), .rst(f320_rst), .rdata(f320_rdata));
  assign f320_clk = clk;
  assign f320_rst = rst;
  // Bindings to f320

  // f316
  logic [0:0] f316_wen;
  logic [31:0] f316_wdata;
  logic [0:0] f316_clk;
  logic [0:0] f316_rst;
  logic [31:0] f316_rdata;
  sr_buffer_32_1 f316(.wen(f316_wen), .wdata(f316_wdata), .clk(f316_clk), .rst(f316_rst), .rdata(f316_rdata));
  assign f316_clk = clk;
  assign f316_rst = rst;
  // Bindings to f316

  // f318
  logic [0:0] f318_wen;
  logic [31:0] f318_wdata;
  logic [0:0] f318_clk;
  logic [0:0] f318_rst;
  logic [31:0] f318_rdata;
  sr_buffer_32_1 f318(.wen(f318_wen), .wdata(f318_wdata), .clk(f318_clk), .rst(f318_rst), .rdata(f318_rdata));
  assign f318_clk = clk;
  assign f318_rst = rst;
  // Bindings to f318

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_16431 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f390
  logic [0:0] f390_wen;
  logic [31:0] f390_wdata;
  logic [0:0] f390_clk;
  logic [0:0] f390_rst;
  logic [31:0] f390_rdata;
  sr_buffer_32_1 f390(.wen(f390_wen), .wdata(f390_wdata), .clk(f390_clk), .rst(f390_rst), .rdata(f390_rdata));
  assign f390_clk = clk;
  assign f390_rst = rst;
  // Bindings to f390

  // f392
  logic [0:0] f392_wen;
  logic [31:0] f392_wdata;
  logic [0:0] f392_clk;
  logic [0:0] f392_rst;
  logic [31:0] f392_rdata;
  sr_buffer_32_1 f392(.wen(f392_wen), .wdata(f392_wdata), .clk(f392_clk), .rst(f392_rst), .rdata(f392_rdata));
  assign f392_clk = clk;
  assign f392_rst = rst;
  // Bindings to f392

  // f394
  logic [0:0] f394_wen;
  logic [31:0] f394_wdata;
  logic [0:0] f394_clk;
  logic [0:0] f394_rst;
  logic [31:0] f394_rdata;
  sr_buffer_32_1 f394(.wen(f394_wen), .wdata(f394_wdata), .clk(f394_clk), .rst(f394_rst), .rdata(f394_rdata));
  assign f394_clk = clk;
  assign f394_rst = rst;
  // Bindings to f394

  // f396
  logic [0:0] f396_wen;
  logic [31:0] f396_wdata;
  logic [0:0] f396_clk;
  logic [0:0] f396_rst;
  logic [31:0] f396_rdata;
  sr_buffer_32_1 f396(.wen(f396_wen), .wdata(f396_wdata), .clk(f396_clk), .rst(f396_rst), .rdata(f396_rdata));
  assign f396_clk = clk;
  assign f396_rst = rst;
  // Bindings to f396

  // f398
  logic [0:0] f398_wen;
  logic [31:0] f398_wdata;
  logic [0:0] f398_clk;
  logic [0:0] f398_rst;
  logic [31:0] f398_rdata;
  sr_buffer_32_1 f398(.wen(f398_wen), .wdata(f398_wdata), .clk(f398_clk), .rst(f398_rst), .rdata(f398_rdata));
  assign f398_clk = clk;
  assign f398_rst = rst;
  // Bindings to f398

  // f400
  logic [0:0] f400_wen;
  logic [31:0] f400_wdata;
  logic [0:0] f400_clk;
  logic [0:0] f400_rst;
  logic [31:0] f400_rdata;
  sr_buffer_32_1 f400(.wen(f400_wen), .wdata(f400_wdata), .clk(f400_clk), .rst(f400_rst), .rdata(f400_rdata));
  assign f400_clk = clk;
  assign f400_rst = rst;
  // Bindings to f400

  // f402
  logic [0:0] f402_wen;
  logic [31:0] f402_wdata;
  logic [0:0] f402_clk;
  logic [0:0] f402_rst;
  logic [31:0] f402_rdata;
  sr_buffer_32_1 f402(.wen(f402_wen), .wdata(f402_wdata), .clk(f402_clk), .rst(f402_rst), .rdata(f402_rdata));
  assign f402_clk = clk;
  assign f402_rst = rst;
  // Bindings to f402

  // f404
  logic [0:0] f404_wen;
  logic [31:0] f404_wdata;
  logic [0:0] f404_clk;
  logic [0:0] f404_rst;
  logic [31:0] f404_rdata;
  sr_buffer_32_1 f404(.wen(f404_wen), .wdata(f404_wdata), .clk(f404_clk), .rst(f404_rst), .rdata(f404_rdata));
  assign f404_clk = clk;
  assign f404_rst = rst;
  // Bindings to f404

  // f406
  logic [0:0] f406_wen;
  logic [31:0] f406_wdata;
  logic [0:0] f406_clk;
  logic [0:0] f406_rst;
  logic [31:0] f406_rdata;
  sr_buffer_32_1 f406(.wen(f406_wen), .wdata(f406_wdata), .clk(f406_clk), .rst(f406_rst), .rdata(f406_rdata));
  assign f406_clk = clk;
  assign f406_rst = rst;
  // Bindings to f406

  // f408
  logic [0:0] f408_wen;
  logic [31:0] f408_wdata;
  logic [0:0] f408_clk;
  logic [0:0] f408_rst;
  logic [31:0] f408_rdata;
  sr_buffer_32_1 f408(.wen(f408_wen), .wdata(f408_wdata), .clk(f408_clk), .rst(f408_rst), .rdata(f408_rdata));
  assign f408_clk = clk;
  assign f408_rst = rst;
  // Bindings to f408

  // f410
  logic [0:0] f410_wen;
  logic [31:0] f410_wdata;
  logic [0:0] f410_clk;
  logic [0:0] f410_rst;
  logic [31:0] f410_rdata;
  sr_buffer_32_1 f410(.wen(f410_wen), .wdata(f410_wdata), .clk(f410_clk), .rst(f410_rst), .rdata(f410_rdata));
  assign f410_clk = clk;
  assign f410_rst = rst;
  // Bindings to f410

  // f412
  logic [0:0] f412_wen;
  logic [31:0] f412_wdata;
  logic [0:0] f412_clk;
  logic [0:0] f412_rst;
  logic [31:0] f412_rdata;
  sr_buffer_32_1 f412(.wen(f412_wen), .wdata(f412_wdata), .clk(f412_clk), .rst(f412_rst), .rdata(f412_rdata));
  assign f412_clk = clk;
  assign f412_rst = rst;
  // Bindings to f412

  // f414
  logic [0:0] f414_wen;
  logic [31:0] f414_wdata;
  logic [0:0] f414_clk;
  logic [0:0] f414_rst;
  logic [31:0] f414_rdata;
  sr_buffer_32_1 f414(.wen(f414_wen), .wdata(f414_wdata), .clk(f414_clk), .rst(f414_rst), .rdata(f414_rdata));
  assign f414_clk = clk;
  assign f414_rst = rst;
  // Bindings to f414

  // f416
  logic [0:0] f416_wen;
  logic [31:0] f416_wdata;
  logic [0:0] f416_clk;
  logic [0:0] f416_rst;
  logic [31:0] f416_rdata;
  sr_buffer_32_1 f416(.wen(f416_wen), .wdata(f416_wdata), .clk(f416_clk), .rst(f416_rst), .rdata(f416_rdata));
  assign f416_clk = clk;
  assign f416_rst = rst;
  // Bindings to f416

  // f418
  logic [0:0] f418_wen;
  logic [31:0] f418_wdata;
  logic [0:0] f418_clk;
  logic [0:0] f418_rst;
  logic [31:0] f418_rdata;
  sr_buffer_32_1 f418(.wen(f418_wen), .wdata(f418_wdata), .clk(f418_clk), .rst(f418_rst), .rdata(f418_rdata));
  assign f418_clk = clk;
  assign f418_rst = rst;
  // Bindings to f418

  // f420
  logic [0:0] f420_wen;
  logic [31:0] f420_wdata;
  logic [0:0] f420_clk;
  logic [0:0] f420_rst;
  logic [31:0] f420_rdata;
  sr_buffer_32_1 f420(.wen(f420_wen), .wdata(f420_wdata), .clk(f420_clk), .rst(f420_rst), .rdata(f420_rdata));
  assign f420_clk = clk;
  assign f420_rst = rst;
  // Bindings to f420

  // f422
  logic [0:0] f422_wen;
  logic [31:0] f422_wdata;
  logic [0:0] f422_clk;
  logic [0:0] f422_rst;
  logic [31:0] f422_rdata;
  sr_buffer_32_1 f422(.wen(f422_wen), .wdata(f422_wdata), .clk(f422_clk), .rst(f422_rst), .rdata(f422_rdata));
  assign f422_clk = clk;
  assign f422_rst = rst;
  // Bindings to f422

  // f424
  logic [0:0] f424_wen;
  logic [31:0] f424_wdata;
  logic [0:0] f424_clk;
  logic [0:0] f424_rst;
  logic [31:0] f424_rdata;
  sr_buffer_32_1 f424(.wen(f424_wen), .wdata(f424_wdata), .clk(f424_clk), .rst(f424_rst), .rdata(f424_rdata));
  assign f424_clk = clk;
  assign f424_rst = rst;
  // Bindings to f424

  // f426
  logic [0:0] f426_wen;
  logic [31:0] f426_wdata;
  logic [0:0] f426_clk;
  logic [0:0] f426_rst;
  logic [31:0] f426_rdata;
  sr_buffer_32_1 f426(.wen(f426_wen), .wdata(f426_wdata), .clk(f426_clk), .rst(f426_rst), .rdata(f426_rdata));
  assign f426_clk = clk;
  assign f426_rst = rst;
  // Bindings to f426

  // f428
  logic [0:0] f428_wen;
  logic [31:0] f428_wdata;
  logic [0:0] f428_clk;
  logic [0:0] f428_rst;
  logic [31:0] f428_rdata;
  sr_buffer_32_1 f428(.wen(f428_wen), .wdata(f428_wdata), .clk(f428_clk), .rst(f428_rst), .rdata(f428_rdata));
  assign f428_clk = clk;
  assign f428_rst = rst;
  // Bindings to f428

  // f430
  logic [0:0] f430_wen;
  logic [31:0] f430_wdata;
  logic [0:0] f430_clk;
  logic [0:0] f430_rst;
  logic [31:0] f430_rdata;
  sr_buffer_32_1 f430(.wen(f430_wen), .wdata(f430_wdata), .clk(f430_clk), .rst(f430_rst), .rdata(f430_rdata));
  assign f430_clk = clk;
  assign f430_rst = rst;
  // Bindings to f430

  // f432
  logic [0:0] f432_wen;
  logic [31:0] f432_wdata;
  logic [0:0] f432_clk;
  logic [0:0] f432_rst;
  logic [31:0] f432_rdata;
  sr_buffer_32_1 f432(.wen(f432_wen), .wdata(f432_wdata), .clk(f432_clk), .rst(f432_rst), .rdata(f432_rdata));
  assign f432_clk = clk;
  assign f432_rst = rst;
  // Bindings to f432

  // f434
  logic [0:0] f434_wen;
  logic [31:0] f434_wdata;
  logic [0:0] f434_clk;
  logic [0:0] f434_rst;
  logic [31:0] f434_rdata;
  sr_buffer_32_1 f434(.wen(f434_wen), .wdata(f434_wdata), .clk(f434_clk), .rst(f434_rst), .rdata(f434_rdata));
  assign f434_clk = clk;
  assign f434_rst = rst;
  // Bindings to f434

  // f436
  logic [0:0] f436_wen;
  logic [31:0] f436_wdata;
  logic [0:0] f436_clk;
  logic [0:0] f436_rst;
  logic [31:0] f436_rdata;
  sr_buffer_32_1 f436(.wen(f436_wen), .wdata(f436_wdata), .clk(f436_clk), .rst(f436_rst), .rdata(f436_rdata));
  assign f436_clk = clk;
  assign f436_rst = rst;
  // Bindings to f436

  // f438
  logic [0:0] f438_wen;
  logic [31:0] f438_wdata;
  logic [0:0] f438_clk;
  logic [0:0] f438_rst;
  logic [31:0] f438_rdata;
  sr_buffer_32_1 f438(.wen(f438_wen), .wdata(f438_wdata), .clk(f438_clk), .rst(f438_rst), .rdata(f438_rdata));
  assign f438_clk = clk;
  assign f438_rst = rst;
  // Bindings to f438

  // f440
  logic [0:0] f440_wen;
  logic [31:0] f440_wdata;
  logic [0:0] f440_clk;
  logic [0:0] f440_rst;
  logic [31:0] f440_rdata;
  sr_buffer_32_1 f440(.wen(f440_wen), .wdata(f440_wdata), .clk(f440_clk), .rst(f440_rst), .rdata(f440_rdata));
  assign f440_clk = clk;
  assign f440_rst = rst;
  // Bindings to f440

  // f442
  logic [0:0] f442_wen;
  logic [31:0] f442_wdata;
  logic [0:0] f442_clk;
  logic [0:0] f442_rst;
  logic [31:0] f442_rdata;
  sr_buffer_32_1 f442(.wen(f442_wen), .wdata(f442_wdata), .clk(f442_clk), .rst(f442_rst), .rdata(f442_rdata));
  assign f442_clk = clk;
  assign f442_rst = rst;
  // Bindings to f442

  // f444
  logic [0:0] f444_wen;
  logic [31:0] f444_wdata;
  logic [0:0] f444_clk;
  logic [0:0] f444_rst;
  logic [31:0] f444_rdata;
  sr_buffer_32_1 f444(.wen(f444_wen), .wdata(f444_wdata), .clk(f444_clk), .rst(f444_rst), .rdata(f444_rdata));
  assign f444_clk = clk;
  assign f444_rst = rst;
  // Bindings to f444

  // f446
  logic [0:0] f446_wen;
  logic [31:0] f446_wdata;
  logic [0:0] f446_clk;
  logic [0:0] f446_rst;
  logic [31:0] f446_rdata;
  sr_buffer_32_1 f446(.wen(f446_wen), .wdata(f446_wdata), .clk(f446_clk), .rst(f446_rst), .rdata(f446_rdata));
  assign f446_clk = clk;
  assign f446_rst = rst;
  // Bindings to f446

  // f448
  logic [0:0] f448_wen;
  logic [31:0] f448_wdata;
  logic [0:0] f448_clk;
  logic [0:0] f448_rst;
  logic [31:0] f448_rdata;
  sr_buffer_32_1 f448(.wen(f448_wen), .wdata(f448_wdata), .clk(f448_clk), .rst(f448_rst), .rdata(f448_rdata));
  assign f448_clk = clk;
  assign f448_rst = rst;
  // Bindings to f448

  // f450
  logic [0:0] f450_wen;
  logic [31:0] f450_wdata;
  logic [0:0] f450_clk;
  logic [0:0] f450_rst;
  logic [31:0] f450_rdata;
  sr_buffer_32_1 f450(.wen(f450_wen), .wdata(f450_wdata), .clk(f450_clk), .rst(f450_rst), .rdata(f450_rdata));
  assign f450_clk = clk;
  assign f450_rst = rst;
  // Bindings to f450

  // f452
  logic [0:0] f452_wen;
  logic [31:0] f452_wdata;
  logic [0:0] f452_clk;
  logic [0:0] f452_rst;
  logic [31:0] f452_rdata;
  sr_buffer_32_1 f452(.wen(f452_wen), .wdata(f452_wdata), .clk(f452_clk), .rst(f452_rst), .rdata(f452_rdata));
  assign f452_clk = clk;
  assign f452_rst = rst;
  // Bindings to f452

  // f454
  logic [0:0] f454_wen;
  logic [31:0] f454_wdata;
  logic [0:0] f454_clk;
  logic [0:0] f454_rst;
  logic [31:0] f454_rdata;
  sr_buffer_32_1 f454(.wen(f454_wen), .wdata(f454_wdata), .clk(f454_clk), .rst(f454_rst), .rdata(f454_rdata));
  assign f454_clk = clk;
  assign f454_rst = rst;
  // Bindings to f454

  // f456
  logic [0:0] f456_wen;
  logic [31:0] f456_wdata;
  logic [0:0] f456_clk;
  logic [0:0] f456_rst;
  logic [31:0] f456_rdata;
  sr_buffer_32_1 f456(.wen(f456_wen), .wdata(f456_wdata), .clk(f456_clk), .rst(f456_rst), .rdata(f456_rdata));
  assign f456_clk = clk;
  assign f456_rst = rst;
  // Bindings to f456

  // f458
  logic [0:0] f458_wen;
  logic [31:0] f458_wdata;
  logic [0:0] f458_clk;
  logic [0:0] f458_rst;
  logic [31:0] f458_rdata;
  sr_buffer_32_1 f458(.wen(f458_wen), .wdata(f458_wdata), .clk(f458_clk), .rst(f458_rst), .rdata(f458_rdata));
  assign f458_clk = clk;
  assign f458_rst = rst;
  // Bindings to f458

  // f460
  logic [0:0] f460_wen;
  logic [31:0] f460_wdata;
  logic [0:0] f460_clk;
  logic [0:0] f460_rst;
  logic [31:0] f460_rdata;
  sr_buffer_32_1 f460(.wen(f460_wen), .wdata(f460_wdata), .clk(f460_clk), .rst(f460_rst), .rdata(f460_rdata));
  assign f460_clk = clk;
  assign f460_rst = rst;
  // Bindings to f460

  // f462
  logic [0:0] f462_wen;
  logic [31:0] f462_wdata;
  logic [0:0] f462_clk;
  logic [0:0] f462_rst;
  logic [31:0] f462_rdata;
  sr_buffer_32_1 f462(.wen(f462_wen), .wdata(f462_wdata), .clk(f462_clk), .rst(f462_rst), .rdata(f462_rdata));
  assign f462_clk = clk;
  assign f462_rst = rst;
  // Bindings to f462

  // f464
  logic [0:0] f464_wen;
  logic [31:0] f464_wdata;
  logic [0:0] f464_clk;
  logic [0:0] f464_rst;
  logic [31:0] f464_rdata;
  sr_buffer_32_1 f464(.wen(f464_wen), .wdata(f464_wdata), .clk(f464_clk), .rst(f464_rst), .rdata(f464_rdata));
  assign f464_clk = clk;
  assign f464_rst = rst;
  // Bindings to f464

  // f466
  logic [0:0] f466_wen;
  logic [31:0] f466_wdata;
  logic [0:0] f466_clk;
  logic [0:0] f466_rst;
  logic [31:0] f466_rdata;
  sr_buffer_32_1 f466(.wen(f466_wen), .wdata(f466_wdata), .clk(f466_clk), .rst(f466_rst), .rdata(f466_rdata));
  assign f466_clk = clk;
  assign f466_rst = rst;
  // Bindings to f466

  // f468
  logic [0:0] f468_wen;
  logic [31:0] f468_wdata;
  logic [0:0] f468_clk;
  logic [0:0] f468_rst;
  logic [31:0] f468_rdata;
  sr_buffer_32_1 f468(.wen(f468_wen), .wdata(f468_wdata), .clk(f468_clk), .rst(f468_rst), .rdata(f468_rdata));
  assign f468_clk = clk;
  assign f468_rst = rst;
  // Bindings to f468

  // f470
  logic [0:0] f470_wen;
  logic [31:0] f470_wdata;
  logic [0:0] f470_clk;
  logic [0:0] f470_rst;
  logic [31:0] f470_rdata;
  sr_buffer_32_1 f470(.wen(f470_wen), .wdata(f470_wdata), .clk(f470_clk), .rst(f470_rst), .rdata(f470_rdata));
  assign f470_clk = clk;
  assign f470_rst = rst;
  // Bindings to f470

  // f472
  logic [0:0] f472_wen;
  logic [31:0] f472_wdata;
  logic [0:0] f472_clk;
  logic [0:0] f472_rst;
  logic [31:0] f472_rdata;
  sr_buffer_32_1 f472(.wen(f472_wen), .wdata(f472_wdata), .clk(f472_clk), .rst(f472_rst), .rdata(f472_rdata));
  assign f472_clk = clk;
  assign f472_rst = rst;
  // Bindings to f472

  // f474
  logic [0:0] f474_wen;
  logic [31:0] f474_wdata;
  logic [0:0] f474_clk;
  logic [0:0] f474_rst;
  logic [31:0] f474_rdata;
  sr_buffer_32_1 f474(.wen(f474_wen), .wdata(f474_wdata), .clk(f474_clk), .rst(f474_rst), .rdata(f474_rdata));
  assign f474_clk = clk;
  assign f474_rst = rst;
  // Bindings to f474

  // f476
  logic [0:0] f476_wen;
  logic [31:0] f476_wdata;
  logic [0:0] f476_clk;
  logic [0:0] f476_rst;
  logic [31:0] f476_rdata;
  sr_buffer_32_1 f476(.wen(f476_wen), .wdata(f476_wdata), .clk(f476_clk), .rst(f476_rst), .rdata(f476_rdata));
  assign f476_clk = clk;
  assign f476_rst = rst;
  // Bindings to f476

  // f478
  logic [0:0] f478_wen;
  logic [31:0] f478_wdata;
  logic [0:0] f478_clk;
  logic [0:0] f478_rst;
  logic [31:0] f478_rdata;
  sr_buffer_32_1 f478(.wen(f478_wen), .wdata(f478_wdata), .clk(f478_clk), .rst(f478_rst), .rdata(f478_rdata));
  assign f478_clk = clk;
  assign f478_rst = rst;
  // Bindings to f478

  // f480
  logic [0:0] f480_wen;
  logic [31:0] f480_wdata;
  logic [0:0] f480_clk;
  logic [0:0] f480_rst;
  logic [31:0] f480_rdata;
  sr_buffer_32_1 f480(.wen(f480_wen), .wdata(f480_wdata), .clk(f480_clk), .rst(f480_rst), .rdata(f480_rdata));
  assign f480_clk = clk;
  assign f480_rst = rst;
  // Bindings to f480

  // f482
  logic [0:0] f482_wen;
  logic [31:0] f482_wdata;
  logic [0:0] f482_clk;
  logic [0:0] f482_rst;
  logic [31:0] f482_rdata;
  sr_buffer_32_1 f482(.wen(f482_wen), .wdata(f482_wdata), .clk(f482_clk), .rst(f482_rst), .rdata(f482_rdata));
  assign f482_clk = clk;
  assign f482_rst = rst;
  // Bindings to f482

  // f484
  logic [0:0] f484_wen;
  logic [31:0] f484_wdata;
  logic [0:0] f484_clk;
  logic [0:0] f484_rst;
  logic [31:0] f484_rdata;
  sr_buffer_32_1 f484(.wen(f484_wen), .wdata(f484_wdata), .clk(f484_clk), .rst(f484_rst), .rdata(f484_rdata));
  assign f484_clk = clk;
  assign f484_rst = rst;
  // Bindings to f484

  // f486
  logic [0:0] f486_wen;
  logic [31:0] f486_wdata;
  logic [0:0] f486_clk;
  logic [0:0] f486_rst;
  logic [31:0] f486_rdata;
  sr_buffer_32_1 f486(.wen(f486_wen), .wdata(f486_wdata), .clk(f486_clk), .rst(f486_rst), .rdata(f486_rdata));
  assign f486_clk = clk;
  assign f486_rst = rst;
  // Bindings to f486

  // f488
  logic [0:0] f488_wen;
  logic [31:0] f488_wdata;
  logic [0:0] f488_clk;
  logic [0:0] f488_rst;
  logic [31:0] f488_rdata;
  sr_buffer_32_1 f488(.wen(f488_wen), .wdata(f488_wdata), .clk(f488_clk), .rst(f488_rst), .rdata(f488_rdata));
  assign f488_clk = clk;
  assign f488_rst = rst;
  // Bindings to f488

  // f490
  logic [0:0] f490_wen;
  logic [31:0] f490_wdata;
  logic [0:0] f490_clk;
  logic [0:0] f490_rst;
  logic [31:0] f490_rdata;
  sr_buffer_32_1 f490(.wen(f490_wen), .wdata(f490_wdata), .clk(f490_clk), .rst(f490_rst), .rdata(f490_rdata));
  assign f490_clk = clk;
  assign f490_rst = rst;
  // Bindings to f490

  // f492
  logic [0:0] f492_wen;
  logic [31:0] f492_wdata;
  logic [0:0] f492_clk;
  logic [0:0] f492_rst;
  logic [31:0] f492_rdata;
  sr_buffer_32_1 f492(.wen(f492_wen), .wdata(f492_wdata), .clk(f492_clk), .rst(f492_rst), .rdata(f492_rdata));
  assign f492_clk = clk;
  assign f492_rst = rst;
  // Bindings to f492

  // f494
  logic [0:0] f494_wen;
  logic [31:0] f494_wdata;
  logic [0:0] f494_clk;
  logic [0:0] f494_rst;
  logic [31:0] f494_rdata;
  sr_buffer_32_1 f494(.wen(f494_wen), .wdata(f494_wdata), .clk(f494_clk), .rst(f494_rst), .rdata(f494_rdata));
  assign f494_clk = clk;
  assign f494_rst = rst;
  // Bindings to f494

  // f496
  logic [0:0] f496_wen;
  logic [31:0] f496_wdata;
  logic [0:0] f496_clk;
  logic [0:0] f496_rst;
  logic [31:0] f496_rdata;
  sr_buffer_32_1 f496(.wen(f496_wen), .wdata(f496_wdata), .clk(f496_clk), .rst(f496_rst), .rdata(f496_rdata));
  assign f496_clk = clk;
  assign f496_rst = rst;
  // Bindings to f496

  // f498
  logic [0:0] f498_wen;
  logic [31:0] f498_wdata;
  logic [0:0] f498_clk;
  logic [0:0] f498_rst;
  logic [31:0] f498_rdata;
  sr_buffer_32_1 f498(.wen(f498_wen), .wdata(f498_wdata), .clk(f498_clk), .rst(f498_rst), .rdata(f498_rdata));
  assign f498_clk = clk;
  assign f498_rst = rst;
  // Bindings to f498

  // f500
  logic [0:0] f500_wen;
  logic [31:0] f500_wdata;
  logic [0:0] f500_clk;
  logic [0:0] f500_rst;
  logic [31:0] f500_rdata;
  sr_buffer_32_1 f500(.wen(f500_wen), .wdata(f500_wdata), .clk(f500_clk), .rst(f500_rst), .rdata(f500_rdata));
  assign f500_clk = clk;
  assign f500_rst = rst;
  // Bindings to f500

  // f502
  logic [0:0] f502_wen;
  logic [31:0] f502_wdata;
  logic [0:0] f502_clk;
  logic [0:0] f502_rst;
  logic [31:0] f502_rdata;
  sr_buffer_32_1 f502(.wen(f502_wen), .wdata(f502_wdata), .clk(f502_clk), .rst(f502_rst), .rdata(f502_rdata));
  assign f502_clk = clk;
  assign f502_rst = rst;
  // Bindings to f502

  // f504
  logic [0:0] f504_wen;
  logic [31:0] f504_wdata;
  logic [0:0] f504_clk;
  logic [0:0] f504_rst;
  logic [31:0] f504_rdata;
  sr_buffer_32_1 f504(.wen(f504_wen), .wdata(f504_wdata), .clk(f504_clk), .rst(f504_rst), .rdata(f504_rdata));
  assign f504_clk = clk;
  assign f504_rst = rst;
  // Bindings to f504

  // f506
  logic [0:0] f506_wen;
  logic [31:0] f506_wdata;
  logic [0:0] f506_clk;
  logic [0:0] f506_rst;
  logic [31:0] f506_rdata;
  sr_buffer_32_1 f506(.wen(f506_wen), .wdata(f506_wdata), .clk(f506_clk), .rst(f506_rst), .rdata(f506_rdata));
  assign f506_clk = clk;
  assign f506_rst = rst;
  // Bindings to f506

  // f508
  logic [0:0] f508_wen;
  logic [31:0] f508_wdata;
  logic [0:0] f508_clk;
  logic [0:0] f508_rst;
  logic [31:0] f508_rdata;
  sr_buffer_32_1 f508(.wen(f508_wen), .wdata(f508_wdata), .clk(f508_clk), .rst(f508_rst), .rdata(f508_rdata));
  assign f508_clk = clk;
  assign f508_rst = rst;
  // Bindings to f508

  // f510
  logic [0:0] f510_wen;
  logic [31:0] f510_wdata;
  logic [0:0] f510_clk;
  logic [0:0] f510_rst;
  logic [31:0] f510_rdata;
  sr_buffer_32_1 f510(.wen(f510_wen), .wdata(f510_wdata), .clk(f510_clk), .rst(f510_rst), .rdata(f510_rdata));
  assign f510_clk = clk;
  assign f510_rst = rst;
  // Bindings to f510

  // f512
  logic [0:0] f512_wen;
  logic [31:0] f512_wdata;
  logic [0:0] f512_clk;
  logic [0:0] f512_rst;
  logic [31:0] f512_rdata;
  sr_buffer_32_1 f512(.wen(f512_wen), .wdata(f512_wdata), .clk(f512_clk), .rst(f512_rst), .rdata(f512_rdata));
  assign f512_clk = clk;
  assign f512_rst = rst;
  // Bindings to f512

  // f514
  logic [0:0] f514_wen;
  logic [31:0] f514_wdata;
  logic [0:0] f514_clk;
  logic [0:0] f514_rst;
  logic [31:0] f514_rdata;
  sr_buffer_32_1 f514(.wen(f514_wen), .wdata(f514_wdata), .clk(f514_clk), .rst(f514_rst), .rdata(f514_rdata));
  assign f514_clk = clk;
  assign f514_rst = rst;
  // Bindings to f514

  // f516
  logic [0:0] f516_wen;
  logic [31:0] f516_wdata;
  logic [0:0] f516_clk;
  logic [0:0] f516_rst;
  logic [31:0] f516_rdata;
  sr_buffer_32_1 f516(.wen(f516_wen), .wdata(f516_wdata), .clk(f516_clk), .rst(f516_rst), .rdata(f516_rdata));
  assign f516_clk = clk;
  assign f516_rst = rst;
  // Bindings to f516

  // f518
  logic [0:0] f518_wen;
  logic [31:0] f518_wdata;
  logic [0:0] f518_clk;
  logic [0:0] f518_rst;
  logic [31:0] f518_rdata;
  sr_buffer_32_1 f518(.wen(f518_wen), .wdata(f518_wdata), .clk(f518_clk), .rst(f518_rst), .rdata(f518_rdata));
  assign f518_clk = clk;
  assign f518_rst = rst;
  // Bindings to f518

  // f520
  logic [0:0] f520_wen;
  logic [31:0] f520_wdata;
  logic [0:0] f520_clk;
  logic [0:0] f520_rst;
  logic [31:0] f520_rdata;
  sr_buffer_32_1 f520(.wen(f520_wen), .wdata(f520_wdata), .clk(f520_clk), .rst(f520_rst), .rdata(f520_rdata));
  assign f520_clk = clk;
  assign f520_rst = rst;
  // Bindings to f520

  // f522
  logic [0:0] f522_wen;
  logic [31:0] f522_wdata;
  logic [0:0] f522_clk;
  logic [0:0] f522_rst;
  logic [31:0] f522_rdata;
  sr_buffer_32_1 f522(.wen(f522_wen), .wdata(f522_wdata), .clk(f522_clk), .rst(f522_rst), .rdata(f522_rdata));
  assign f522_clk = clk;
  assign f522_rst = rst;
  // Bindings to f522

  // f524
  logic [0:0] f524_wen;
  logic [31:0] f524_wdata;
  logic [0:0] f524_clk;
  logic [0:0] f524_rst;
  logic [31:0] f524_rdata;
  sr_buffer_32_1 f524(.wen(f524_wen), .wdata(f524_wdata), .clk(f524_clk), .rst(f524_rst), .rdata(f524_rdata));
  assign f524_clk = clk;
  assign f524_rst = rst;
  // Bindings to f524

  // f526
  logic [0:0] f526_wen;
  logic [31:0] f526_wdata;
  logic [0:0] f526_clk;
  logic [0:0] f526_rst;
  logic [31:0] f526_rdata;
  sr_buffer_32_1 f526(.wen(f526_wen), .wdata(f526_wdata), .clk(f526_clk), .rst(f526_rst), .rdata(f526_rdata));
  assign f526_clk = clk;
  assign f526_rst = rst;
  // Bindings to f526

  // f528
  logic [0:0] f528_wen;
  logic [31:0] f528_wdata;
  logic [0:0] f528_clk;
  logic [0:0] f528_rst;
  logic [31:0] f528_rdata;
  sr_buffer_32_1 f528(.wen(f528_wen), .wdata(f528_wdata), .clk(f528_clk), .rst(f528_rst), .rdata(f528_rdata));
  assign f528_clk = clk;
  assign f528_rst = rst;
  // Bindings to f528

  // f530
  logic [0:0] f530_wen;
  logic [31:0] f530_wdata;
  logic [0:0] f530_clk;
  logic [0:0] f530_rst;
  logic [31:0] f530_rdata;
  sr_buffer_32_1 f530(.wen(f530_wen), .wdata(f530_wdata), .clk(f530_clk), .rst(f530_rst), .rdata(f530_rdata));
  assign f530_clk = clk;
  assign f530_rst = rst;
  // Bindings to f530

  // f532
  logic [0:0] f532_wen;
  logic [31:0] f532_wdata;
  logic [0:0] f532_clk;
  logic [0:0] f532_rst;
  logic [31:0] f532_rdata;
  sr_buffer_32_1 f532(.wen(f532_wen), .wdata(f532_wdata), .clk(f532_clk), .rst(f532_rst), .rdata(f532_rdata));
  assign f532_clk = clk;
  assign f532_rst = rst;
  // Bindings to f532

  // f534
  logic [0:0] f534_wen;
  logic [31:0] f534_wdata;
  logic [0:0] f534_clk;
  logic [0:0] f534_rst;
  logic [31:0] f534_rdata;
  sr_buffer_32_1 f534(.wen(f534_wen), .wdata(f534_wdata), .clk(f534_clk), .rst(f534_rst), .rdata(f534_rdata));
  assign f534_clk = clk;
  assign f534_rst = rst;
  // Bindings to f534

  // f536
  logic [0:0] f536_wen;
  logic [31:0] f536_wdata;
  logic [0:0] f536_clk;
  logic [0:0] f536_rst;
  logic [31:0] f536_rdata;
  sr_buffer_32_1 f536(.wen(f536_wen), .wdata(f536_wdata), .clk(f536_clk), .rst(f536_rst), .rdata(f536_rdata));
  assign f536_clk = clk;
  assign f536_rst = rst;
  // Bindings to f536

  // f538
  logic [0:0] f538_wen;
  logic [31:0] f538_wdata;
  logic [0:0] f538_clk;
  logic [0:0] f538_rst;
  logic [31:0] f538_rdata;
  sr_buffer_32_1 f538(.wen(f538_wen), .wdata(f538_wdata), .clk(f538_clk), .rst(f538_rst), .rdata(f538_rdata));
  assign f538_clk = clk;
  assign f538_rst = rst;
  // Bindings to f538

  // f540
  logic [0:0] f540_wen;
  logic [31:0] f540_wdata;
  logic [0:0] f540_clk;
  logic [0:0] f540_rst;
  logic [31:0] f540_rdata;
  sr_buffer_32_1 f540(.wen(f540_wen), .wdata(f540_wdata), .clk(f540_clk), .rst(f540_rst), .rdata(f540_rdata));
  assign f540_clk = clk;
  assign f540_rst = rst;
  // Bindings to f540

  // f542
  logic [0:0] f542_wen;
  logic [31:0] f542_wdata;
  logic [0:0] f542_clk;
  logic [0:0] f542_rst;
  logic [31:0] f542_rdata;
  sr_buffer_32_1 f542(.wen(f542_wen), .wdata(f542_wdata), .clk(f542_clk), .rst(f542_rst), .rdata(f542_rdata));
  assign f542_clk = clk;
  assign f542_rst = rst;
  // Bindings to f542

  // f544
  logic [0:0] f544_wen;
  logic [31:0] f544_wdata;
  logic [0:0] f544_clk;
  logic [0:0] f544_rst;
  logic [31:0] f544_rdata;
  sr_buffer_32_1 f544(.wen(f544_wen), .wdata(f544_wdata), .clk(f544_clk), .rst(f544_rst), .rdata(f544_rdata));
  assign f544_clk = clk;
  assign f544_rst = rst;
  // Bindings to f544

  // f546
  logic [0:0] f546_wen;
  logic [31:0] f546_wdata;
  logic [0:0] f546_clk;
  logic [0:0] f546_rst;
  logic [31:0] f546_rdata;
  sr_buffer_32_1 f546(.wen(f546_wen), .wdata(f546_wdata), .clk(f546_clk), .rst(f546_rst), .rdata(f546_rdata));
  assign f546_clk = clk;
  assign f546_rst = rst;
  // Bindings to f546

  // f548
  logic [0:0] f548_wen;
  logic [31:0] f548_wdata;
  logic [0:0] f548_clk;
  logic [0:0] f548_rst;
  logic [31:0] f548_rdata;
  sr_buffer_32_1 f548(.wen(f548_wen), .wdata(f548_wdata), .clk(f548_clk), .rst(f548_rst), .rdata(f548_rdata));
  assign f548_clk = clk;
  assign f548_rst = rst;
  // Bindings to f548

  // f550
  logic [0:0] f550_wen;
  logic [31:0] f550_wdata;
  logic [0:0] f550_clk;
  logic [0:0] f550_rst;
  logic [31:0] f550_rdata;
  sr_buffer_32_1 f550(.wen(f550_wen), .wdata(f550_wdata), .clk(f550_clk), .rst(f550_rst), .rdata(f550_rdata));
  assign f550_clk = clk;
  assign f550_rst = rst;
  // Bindings to f550

  // f552
  logic [0:0] f552_wen;
  logic [31:0] f552_wdata;
  logic [0:0] f552_clk;
  logic [0:0] f552_rst;
  logic [31:0] f552_rdata;
  sr_buffer_32_1 f552(.wen(f552_wen), .wdata(f552_wdata), .clk(f552_clk), .rst(f552_rst), .rdata(f552_rdata));
  assign f552_clk = clk;
  assign f552_rst = rst;
  // Bindings to f552

  // f554
  logic [0:0] f554_wen;
  logic [31:0] f554_wdata;
  logic [0:0] f554_clk;
  logic [0:0] f554_rst;
  logic [31:0] f554_rdata;
  sr_buffer_32_1 f554(.wen(f554_wen), .wdata(f554_wdata), .clk(f554_clk), .rst(f554_rst), .rdata(f554_rdata));
  assign f554_clk = clk;
  assign f554_rst = rst;
  // Bindings to f554

  // f556
  logic [0:0] f556_wen;
  logic [31:0] f556_wdata;
  logic [0:0] f556_clk;
  logic [0:0] f556_rst;
  logic [31:0] f556_rdata;
  sr_buffer_32_1 f556(.wen(f556_wen), .wdata(f556_wdata), .clk(f556_clk), .rst(f556_rst), .rdata(f556_rdata));
  assign f556_clk = clk;
  assign f556_rst = rst;
  // Bindings to f556

  // f558
  logic [0:0] f558_wen;
  logic [31:0] f558_wdata;
  logic [0:0] f558_clk;
  logic [0:0] f558_rst;
  logic [31:0] f558_rdata;
  sr_buffer_32_1 f558(.wen(f558_wen), .wdata(f558_wdata), .clk(f558_clk), .rst(f558_rst), .rdata(f558_rdata));
  assign f558_clk = clk;
  assign f558_rst = rst;
  // Bindings to f558

  // f560
  logic [0:0] f560_wen;
  logic [31:0] f560_wdata;
  logic [0:0] f560_clk;
  logic [0:0] f560_rst;
  logic [31:0] f560_rdata;
  sr_buffer_32_1 f560(.wen(f560_wen), .wdata(f560_wdata), .clk(f560_clk), .rst(f560_rst), .rdata(f560_rdata));
  assign f560_clk = clk;
  assign f560_rst = rst;
  // Bindings to f560

  // f562
  logic [0:0] f562_wen;
  logic [31:0] f562_wdata;
  logic [0:0] f562_clk;
  logic [0:0] f562_rst;
  logic [31:0] f562_rdata;
  sr_buffer_32_1 f562(.wen(f562_wen), .wdata(f562_wdata), .clk(f562_clk), .rst(f562_rst), .rdata(f562_rdata));
  assign f562_clk = clk;
  assign f562_rst = rst;
  // Bindings to f562

  // f564
  logic [0:0] f564_wen;
  logic [31:0] f564_wdata;
  logic [0:0] f564_clk;
  logic [0:0] f564_rst;
  logic [31:0] f564_rdata;
  sr_buffer_32_1 f564(.wen(f564_wen), .wdata(f564_wdata), .clk(f564_clk), .rst(f564_rst), .rdata(f564_rdata));
  assign f564_clk = clk;
  assign f564_rst = rst;
  // Bindings to f564

  // f566
  logic [0:0] f566_wen;
  logic [31:0] f566_wdata;
  logic [0:0] f566_clk;
  logic [0:0] f566_rst;
  logic [31:0] f566_rdata;
  sr_buffer_32_1 f566(.wen(f566_wen), .wdata(f566_wdata), .clk(f566_clk), .rst(f566_rst), .rdata(f566_rdata));
  assign f566_clk = clk;
  assign f566_rst = rst;
  // Bindings to f566

  // f568
  logic [0:0] f568_wen;
  logic [31:0] f568_wdata;
  logic [0:0] f568_clk;
  logic [0:0] f568_rst;
  logic [31:0] f568_rdata;
  sr_buffer_32_1 f568(.wen(f568_wen), .wdata(f568_wdata), .clk(f568_clk), .rst(f568_rst), .rdata(f568_rdata));
  assign f568_clk = clk;
  assign f568_rst = rst;
  // Bindings to f568

  // f570
  logic [0:0] f570_wen;
  logic [31:0] f570_wdata;
  logic [0:0] f570_clk;
  logic [0:0] f570_rst;
  logic [31:0] f570_rdata;
  sr_buffer_32_1 f570(.wen(f570_wen), .wdata(f570_wdata), .clk(f570_clk), .rst(f570_rst), .rdata(f570_rdata));
  assign f570_clk = clk;
  assign f570_rst = rst;
  // Bindings to f570

  // f572
  logic [0:0] f572_wen;
  logic [31:0] f572_wdata;
  logic [0:0] f572_clk;
  logic [0:0] f572_rst;
  logic [31:0] f572_rdata;
  sr_buffer_32_1 f572(.wen(f572_wen), .wdata(f572_wdata), .clk(f572_clk), .rst(f572_rst), .rdata(f572_rdata));
  assign f572_clk = clk;
  assign f572_rst = rst;
  // Bindings to f572

  // f574
  logic [0:0] f574_wen;
  logic [31:0] f574_wdata;
  logic [0:0] f574_clk;
  logic [0:0] f574_rst;
  logic [31:0] f574_rdata;
  sr_buffer_32_1 f574(.wen(f574_wen), .wdata(f574_wdata), .clk(f574_clk), .rst(f574_rst), .rdata(f574_rdata));
  assign f574_clk = clk;
  assign f574_rst = rst;
  // Bindings to f574

  // f576
  logic [0:0] f576_wen;
  logic [31:0] f576_wdata;
  logic [0:0] f576_clk;
  logic [0:0] f576_rst;
  logic [31:0] f576_rdata;
  sr_buffer_32_1 f576(.wen(f576_wen), .wdata(f576_wdata), .clk(f576_clk), .rst(f576_rst), .rdata(f576_rdata));
  assign f576_clk = clk;
  assign f576_rst = rst;
  // Bindings to f576

  // f578
  logic [0:0] f578_wen;
  logic [31:0] f578_wdata;
  logic [0:0] f578_clk;
  logic [0:0] f578_rst;
  logic [31:0] f578_rdata;
  sr_buffer_32_1 f578(.wen(f578_wen), .wdata(f578_wdata), .clk(f578_clk), .rst(f578_rst), .rdata(f578_rdata));
  assign f578_clk = clk;
  assign f578_rst = rst;
  // Bindings to f578

  // f580
  logic [0:0] f580_wen;
  logic [31:0] f580_wdata;
  logic [0:0] f580_clk;
  logic [0:0] f580_rst;
  logic [31:0] f580_rdata;
  sr_buffer_32_1 f580(.wen(f580_wen), .wdata(f580_wdata), .clk(f580_clk), .rst(f580_rst), .rdata(f580_rdata));
  assign f580_clk = clk;
  assign f580_rst = rst;
  // Bindings to f580

  // f582
  logic [0:0] f582_wen;
  logic [31:0] f582_wdata;
  logic [0:0] f582_clk;
  logic [0:0] f582_rst;
  logic [31:0] f582_rdata;
  sr_buffer_32_1 f582(.wen(f582_wen), .wdata(f582_wdata), .clk(f582_clk), .rst(f582_rst), .rdata(f582_rdata));
  assign f582_clk = clk;
  assign f582_rst = rst;
  // Bindings to f582

  // f584
  logic [0:0] f584_wen;
  logic [31:0] f584_wdata;
  logic [0:0] f584_clk;
  logic [0:0] f584_rst;
  logic [31:0] f584_rdata;
  sr_buffer_32_1 f584(.wen(f584_wen), .wdata(f584_wdata), .clk(f584_clk), .rst(f584_rst), .rdata(f584_rdata));
  assign f584_clk = clk;
  assign f584_rst = rst;
  // Bindings to f584

  // f586
  logic [0:0] f586_wen;
  logic [31:0] f586_wdata;
  logic [0:0] f586_clk;
  logic [0:0] f586_rst;
  logic [31:0] f586_rdata;
  sr_buffer_32_1 f586(.wen(f586_wen), .wdata(f586_wdata), .clk(f586_clk), .rst(f586_rst), .rdata(f586_rdata));
  assign f586_clk = clk;
  assign f586_rst = rst;
  // Bindings to f586

  // f588
  logic [0:0] f588_wen;
  logic [31:0] f588_wdata;
  logic [0:0] f588_clk;
  logic [0:0] f588_rst;
  logic [31:0] f588_rdata;
  sr_buffer_32_1 f588(.wen(f588_wen), .wdata(f588_wdata), .clk(f588_clk), .rst(f588_rst), .rdata(f588_rdata));
  assign f588_clk = clk;
  assign f588_rst = rst;
  // Bindings to f588

  // f590
  logic [0:0] f590_wen;
  logic [31:0] f590_wdata;
  logic [0:0] f590_clk;
  logic [0:0] f590_rst;
  logic [31:0] f590_rdata;
  sr_buffer_32_1 f590(.wen(f590_wen), .wdata(f590_wdata), .clk(f590_clk), .rst(f590_rst), .rdata(f590_rdata));
  assign f590_clk = clk;
  assign f590_rst = rst;
  // Bindings to f590

  // f592
  logic [0:0] f592_wen;
  logic [31:0] f592_wdata;
  logic [0:0] f592_clk;
  logic [0:0] f592_rst;
  logic [31:0] f592_rdata;
  sr_buffer_32_1 f592(.wen(f592_wen), .wdata(f592_wdata), .clk(f592_clk), .rst(f592_rst), .rdata(f592_rdata));
  assign f592_clk = clk;
  assign f592_rst = rst;
  // Bindings to f592

  // f594
  logic [0:0] f594_wen;
  logic [31:0] f594_wdata;
  logic [0:0] f594_clk;
  logic [0:0] f594_rst;
  logic [31:0] f594_rdata;
  sr_buffer_32_1 f594(.wen(f594_wen), .wdata(f594_wdata), .clk(f594_clk), .rst(f594_rst), .rdata(f594_rdata));
  assign f594_clk = clk;
  assign f594_rst = rst;
  // Bindings to f594

  // f596
  logic [0:0] f596_wen;
  logic [31:0] f596_wdata;
  logic [0:0] f596_clk;
  logic [0:0] f596_rst;
  logic [31:0] f596_rdata;
  sr_buffer_32_1 f596(.wen(f596_wen), .wdata(f596_wdata), .clk(f596_clk), .rst(f596_rst), .rdata(f596_rdata));
  assign f596_clk = clk;
  assign f596_rst = rst;
  // Bindings to f596

  // f598
  logic [0:0] f598_wen;
  logic [31:0] f598_wdata;
  logic [0:0] f598_clk;
  logic [0:0] f598_rst;
  logic [31:0] f598_rdata;
  sr_buffer_32_1 f598(.wen(f598_wen), .wdata(f598_wdata), .clk(f598_clk), .rst(f598_rst), .rdata(f598_rdata));
  assign f598_clk = clk;
  assign f598_rst = rst;
  // Bindings to f598

  // f600
  logic [0:0] f600_wen;
  logic [31:0] f600_wdata;
  logic [0:0] f600_clk;
  logic [0:0] f600_rst;
  logic [31:0] f600_rdata;
  sr_buffer_32_1 f600(.wen(f600_wen), .wdata(f600_wdata), .clk(f600_clk), .rst(f600_rst), .rdata(f600_rdata));
  assign f600_clk = clk;
  assign f600_rst = rst;
  // Bindings to f600

  // f602
  logic [0:0] f602_wen;
  logic [31:0] f602_wdata;
  logic [0:0] f602_clk;
  logic [0:0] f602_rst;
  logic [31:0] f602_rdata;
  sr_buffer_32_1 f602(.wen(f602_wen), .wdata(f602_wdata), .clk(f602_clk), .rst(f602_rst), .rdata(f602_rdata));
  assign f602_clk = clk;
  assign f602_rst = rst;
  // Bindings to f602

  // f604
  logic [0:0] f604_wen;
  logic [31:0] f604_wdata;
  logic [0:0] f604_clk;
  logic [0:0] f604_rst;
  logic [31:0] f604_rdata;
  sr_buffer_32_1 f604(.wen(f604_wen), .wdata(f604_wdata), .clk(f604_clk), .rst(f604_rst), .rdata(f604_rdata));
  assign f604_clk = clk;
  assign f604_rst = rst;
  // Bindings to f604

  // f606
  logic [0:0] f606_wen;
  logic [31:0] f606_wdata;
  logic [0:0] f606_clk;
  logic [0:0] f606_rst;
  logic [31:0] f606_rdata;
  sr_buffer_32_1 f606(.wen(f606_wen), .wdata(f606_wdata), .clk(f606_clk), .rst(f606_rst), .rdata(f606_rdata));
  assign f606_clk = clk;
  assign f606_rst = rst;
  // Bindings to f606

  // f608
  logic [0:0] f608_wen;
  logic [31:0] f608_wdata;
  logic [0:0] f608_clk;
  logic [0:0] f608_rst;
  logic [31:0] f608_rdata;
  sr_buffer_32_1 f608(.wen(f608_wen), .wdata(f608_wdata), .clk(f608_clk), .rst(f608_rst), .rdata(f608_rdata));
  assign f608_clk = clk;
  assign f608_rst = rst;
  // Bindings to f608

  // f610
  logic [0:0] f610_wen;
  logic [31:0] f610_wdata;
  logic [0:0] f610_clk;
  logic [0:0] f610_rst;
  logic [31:0] f610_rdata;
  sr_buffer_32_1 f610(.wen(f610_wen), .wdata(f610_wdata), .clk(f610_clk), .rst(f610_rst), .rdata(f610_rdata));
  assign f610_clk = clk;
  assign f610_rst = rst;
  // Bindings to f610

  // f612
  logic [0:0] f612_wen;
  logic [31:0] f612_wdata;
  logic [0:0] f612_clk;
  logic [0:0] f612_rst;
  logic [31:0] f612_rdata;
  sr_buffer_32_1 f612(.wen(f612_wen), .wdata(f612_wdata), .clk(f612_clk), .rst(f612_rst), .rdata(f612_rdata));
  assign f612_clk = clk;
  assign f612_rst = rst;
  // Bindings to f612

  // f614
  logic [0:0] f614_wen;
  logic [31:0] f614_wdata;
  logic [0:0] f614_clk;
  logic [0:0] f614_rst;
  logic [31:0] f614_rdata;
  sr_buffer_32_1 f614(.wen(f614_wen), .wdata(f614_wdata), .clk(f614_clk), .rst(f614_rst), .rdata(f614_rdata));
  assign f614_clk = clk;
  assign f614_rst = rst;
  // Bindings to f614

  // f616
  logic [0:0] f616_wen;
  logic [31:0] f616_wdata;
  logic [0:0] f616_clk;
  logic [0:0] f616_rst;
  logic [31:0] f616_rdata;
  sr_buffer_32_1 f616(.wen(f616_wen), .wdata(f616_wdata), .clk(f616_clk), .rst(f616_rst), .rdata(f616_rdata));
  assign f616_clk = clk;
  assign f616_rst = rst;
  // Bindings to f616

  // f618
  logic [0:0] f618_wen;
  logic [31:0] f618_wdata;
  logic [0:0] f618_clk;
  logic [0:0] f618_rst;
  logic [31:0] f618_rdata;
  sr_buffer_32_1 f618(.wen(f618_wen), .wdata(f618_wdata), .clk(f618_clk), .rst(f618_rst), .rdata(f618_rdata));
  assign f618_clk = clk;
  assign f618_rst = rst;
  // Bindings to f618

  // f620
  logic [0:0] f620_wen;
  logic [31:0] f620_wdata;
  logic [0:0] f620_clk;
  logic [0:0] f620_rst;
  logic [31:0] f620_rdata;
  sr_buffer_32_1 f620(.wen(f620_wen), .wdata(f620_wdata), .clk(f620_clk), .rst(f620_rst), .rdata(f620_rdata));
  assign f620_clk = clk;
  assign f620_rst = rst;
  // Bindings to f620

  // f622
  logic [0:0] f622_wen;
  logic [31:0] f622_wdata;
  logic [0:0] f622_clk;
  logic [0:0] f622_rst;
  logic [31:0] f622_rdata;
  sr_buffer_32_1 f622(.wen(f622_wen), .wdata(f622_wdata), .clk(f622_clk), .rst(f622_rst), .rdata(f622_rdata));
  assign f622_clk = clk;
  assign f622_rst = rst;
  // Bindings to f622

  // f624
  logic [0:0] f624_wen;
  logic [31:0] f624_wdata;
  logic [0:0] f624_clk;
  logic [0:0] f624_rst;
  logic [31:0] f624_rdata;
  sr_buffer_32_1 f624(.wen(f624_wen), .wdata(f624_wdata), .clk(f624_clk), .rst(f624_rst), .rdata(f624_rdata));
  assign f624_clk = clk;
  assign f624_rst = rst;
  // Bindings to f624

  // f626
  logic [0:0] f626_wen;
  logic [31:0] f626_wdata;
  logic [0:0] f626_clk;
  logic [0:0] f626_rst;
  logic [31:0] f626_rdata;
  sr_buffer_32_1 f626(.wen(f626_wen), .wdata(f626_wdata), .clk(f626_clk), .rst(f626_rst), .rdata(f626_rdata));
  assign f626_clk = clk;
  assign f626_rst = rst;
  // Bindings to f626

  // f628
  logic [0:0] f628_wen;
  logic [31:0] f628_wdata;
  logic [0:0] f628_clk;
  logic [0:0] f628_rst;
  logic [31:0] f628_rdata;
  sr_buffer_32_1 f628(.wen(f628_wen), .wdata(f628_wdata), .clk(f628_clk), .rst(f628_rst), .rdata(f628_rdata));
  assign f628_clk = clk;
  assign f628_rst = rst;
  // Bindings to f628

  // f630
  logic [0:0] f630_wen;
  logic [31:0] f630_wdata;
  logic [0:0] f630_clk;
  logic [0:0] f630_rst;
  logic [31:0] f630_rdata;
  sr_buffer_32_1 f630(.wen(f630_wen), .wdata(f630_wdata), .clk(f630_clk), .rst(f630_rst), .rdata(f630_rdata));
  assign f630_clk = clk;
  assign f630_rst = rst;
  // Bindings to f630

  // f632
  logic [0:0] f632_wen;
  logic [31:0] f632_wdata;
  logic [0:0] f632_clk;
  logic [0:0] f632_rst;
  logic [31:0] f632_rdata;
  sr_buffer_32_1 f632(.wen(f632_wen), .wdata(f632_wdata), .clk(f632_clk), .rst(f632_rst), .rdata(f632_rdata));
  assign f632_clk = clk;
  assign f632_rst = rst;
  // Bindings to f632

  // f634
  logic [0:0] f634_wen;
  logic [31:0] f634_wdata;
  logic [0:0] f634_clk;
  logic [0:0] f634_rst;
  logic [31:0] f634_rdata;
  sr_buffer_32_1 f634(.wen(f634_wen), .wdata(f634_wdata), .clk(f634_clk), .rst(f634_rst), .rdata(f634_rdata));
  assign f634_clk = clk;
  assign f634_rst = rst;
  // Bindings to f634

  // f636
  logic [0:0] f636_wen;
  logic [31:0] f636_wdata;
  logic [0:0] f636_clk;
  logic [0:0] f636_rst;
  logic [31:0] f636_rdata;
  sr_buffer_32_1 f636(.wen(f636_wen), .wdata(f636_wdata), .clk(f636_clk), .rst(f636_rst), .rdata(f636_rdata));
  assign f636_clk = clk;
  assign f636_rst = rst;
  // Bindings to f636

  // f638
  logic [0:0] f638_wen;
  logic [31:0] f638_wdata;
  logic [0:0] f638_clk;
  logic [0:0] f638_rst;
  logic [31:0] f638_rdata;
  sr_buffer_32_1 f638(.wen(f638_wen), .wdata(f638_wdata), .clk(f638_clk), .rst(f638_rst), .rdata(f638_rdata));
  assign f638_clk = clk;
  assign f638_rst = rst;
  // Bindings to f638

  // f640
  logic [0:0] f640_wen;
  logic [31:0] f640_wdata;
  logic [0:0] f640_clk;
  logic [0:0] f640_rst;
  logic [31:0] f640_rdata;
  sr_buffer_32_1 f640(.wen(f640_wen), .wdata(f640_wdata), .clk(f640_clk), .rst(f640_rst), .rdata(f640_rdata));
  assign f640_clk = clk;
  assign f640_rst = rst;
  // Bindings to f640

  // f642
  logic [0:0] f642_wen;
  logic [31:0] f642_wdata;
  logic [0:0] f642_clk;
  logic [0:0] f642_rst;
  logic [31:0] f642_rdata;
  sr_buffer_32_1 f642(.wen(f642_wen), .wdata(f642_wdata), .clk(f642_clk), .rst(f642_rst), .rdata(f642_rdata));
  assign f642_clk = clk;
  assign f642_rst = rst;
  // Bindings to f642

  // f644
  logic [0:0] f644_wen;
  logic [31:0] f644_wdata;
  logic [0:0] f644_clk;
  logic [0:0] f644_rst;
  logic [31:0] f644_rdata;
  sr_buffer_32_1 f644(.wen(f644_wen), .wdata(f644_wdata), .clk(f644_clk), .rst(f644_rst), .rdata(f644_rdata));
  assign f644_clk = clk;
  assign f644_rst = rst;
  // Bindings to f644

  // f646
  logic [0:0] f646_wen;
  logic [31:0] f646_wdata;
  logic [0:0] f646_clk;
  logic [0:0] f646_rst;
  logic [31:0] f646_rdata;
  sr_buffer_32_1 f646(.wen(f646_wen), .wdata(f646_wdata), .clk(f646_clk), .rst(f646_rst), .rdata(f646_rdata));
  assign f646_clk = clk;
  assign f646_rst = rst;
  // Bindings to f646

  // f648
  logic [0:0] f648_wen;
  logic [31:0] f648_wdata;
  logic [0:0] f648_clk;
  logic [0:0] f648_rst;
  logic [31:0] f648_rdata;
  sr_buffer_32_1 f648(.wen(f648_wen), .wdata(f648_wdata), .clk(f648_clk), .rst(f648_rst), .rdata(f648_rdata));
  assign f648_clk = clk;
  assign f648_rst = rst;
  // Bindings to f648

  // f650
  logic [0:0] f650_wen;
  logic [31:0] f650_wdata;
  logic [0:0] f650_clk;
  logic [0:0] f650_rst;
  logic [31:0] f650_rdata;
  sr_buffer_32_1 f650(.wen(f650_wen), .wdata(f650_wdata), .clk(f650_clk), .rst(f650_rst), .rdata(f650_rdata));
  assign f650_clk = clk;
  assign f650_rst = rst;
  // Bindings to f650

  // f652
  logic [0:0] f652_wen;
  logic [31:0] f652_wdata;
  logic [0:0] f652_clk;
  logic [0:0] f652_rst;
  logic [31:0] f652_rdata;
  sr_buffer_32_1 f652(.wen(f652_wen), .wdata(f652_wdata), .clk(f652_clk), .rst(f652_rst), .rdata(f652_rdata));
  assign f652_clk = clk;
  assign f652_rst = rst;
  // Bindings to f652

  // f654
  logic [0:0] f654_wen;
  logic [31:0] f654_wdata;
  logic [0:0] f654_clk;
  logic [0:0] f654_rst;
  logic [31:0] f654_rdata;
  sr_buffer_32_1 f654(.wen(f654_wen), .wdata(f654_wdata), .clk(f654_clk), .rst(f654_rst), .rdata(f654_rdata));
  assign f654_clk = clk;
  assign f654_rst = rst;
  // Bindings to f654

  // f656
  logic [0:0] f656_wen;
  logic [31:0] f656_wdata;
  logic [0:0] f656_clk;
  logic [0:0] f656_rst;
  logic [31:0] f656_rdata;
  sr_buffer_32_1 f656(.wen(f656_wen), .wdata(f656_wdata), .clk(f656_clk), .rst(f656_rst), .rdata(f656_rdata));
  assign f656_clk = clk;
  assign f656_rst = rst;
  // Bindings to f656

  // f658
  logic [0:0] f658_wen;
  logic [31:0] f658_wdata;
  logic [0:0] f658_clk;
  logic [0:0] f658_rst;
  logic [31:0] f658_rdata;
  sr_buffer_32_1 f658(.wen(f658_wen), .wdata(f658_wdata), .clk(f658_clk), .rst(f658_rst), .rdata(f658_rdata));
  assign f658_clk = clk;
  assign f658_rst = rst;
  // Bindings to f658

  // f660
  logic [0:0] f660_wen;
  logic [31:0] f660_wdata;
  logic [0:0] f660_clk;
  logic [0:0] f660_rst;
  logic [31:0] f660_rdata;
  sr_buffer_32_1 f660(.wen(f660_wen), .wdata(f660_wdata), .clk(f660_clk), .rst(f660_rst), .rdata(f660_rdata));
  assign f660_clk = clk;
  assign f660_rst = rst;
  // Bindings to f660

  // f662
  logic [0:0] f662_wen;
  logic [31:0] f662_wdata;
  logic [0:0] f662_clk;
  logic [0:0] f662_rst;
  logic [31:0] f662_rdata;
  sr_buffer_32_1 f662(.wen(f662_wen), .wdata(f662_wdata), .clk(f662_clk), .rst(f662_rst), .rdata(f662_rdata));
  assign f662_clk = clk;
  assign f662_rst = rst;
  // Bindings to f662

  // f664
  logic [0:0] f664_wen;
  logic [31:0] f664_wdata;
  logic [0:0] f664_clk;
  logic [0:0] f664_rst;
  logic [31:0] f664_rdata;
  sr_buffer_32_1 f664(.wen(f664_wen), .wdata(f664_wdata), .clk(f664_clk), .rst(f664_rst), .rdata(f664_rdata));
  assign f664_clk = clk;
  assign f664_rst = rst;
  // Bindings to f664

  // f666
  logic [0:0] f666_wen;
  logic [31:0] f666_wdata;
  logic [0:0] f666_clk;
  logic [0:0] f666_rst;
  logic [31:0] f666_rdata;
  sr_buffer_32_1 f666(.wen(f666_wen), .wdata(f666_wdata), .clk(f666_clk), .rst(f666_rst), .rdata(f666_rdata));
  assign f666_clk = clk;
  assign f666_rst = rst;
  // Bindings to f666

  // f668
  logic [0:0] f668_wen;
  logic [31:0] f668_wdata;
  logic [0:0] f668_clk;
  logic [0:0] f668_rst;
  logic [31:0] f668_rdata;
  sr_buffer_32_1 f668(.wen(f668_wen), .wdata(f668_wdata), .clk(f668_clk), .rst(f668_rst), .rdata(f668_rdata));
  assign f668_clk = clk;
  assign f668_rst = rst;
  // Bindings to f668

  // f670
  logic [0:0] f670_wen;
  logic [31:0] f670_wdata;
  logic [0:0] f670_clk;
  logic [0:0] f670_rst;
  logic [31:0] f670_rdata;
  sr_buffer_32_1 f670(.wen(f670_wen), .wdata(f670_wdata), .clk(f670_clk), .rst(f670_rst), .rdata(f670_rdata));
  assign f670_clk = clk;
  assign f670_rst = rst;
  // Bindings to f670

  // f672
  logic [0:0] f672_wen;
  logic [31:0] f672_wdata;
  logic [0:0] f672_clk;
  logic [0:0] f672_rst;
  logic [31:0] f672_rdata;
  sr_buffer_32_1 f672(.wen(f672_wen), .wdata(f672_wdata), .clk(f672_clk), .rst(f672_rst), .rdata(f672_rdata));
  assign f672_clk = clk;
  assign f672_rst = rst;
  // Bindings to f672

  // f674
  logic [0:0] f674_wen;
  logic [31:0] f674_wdata;
  logic [0:0] f674_clk;
  logic [0:0] f674_rst;
  logic [31:0] f674_rdata;
  sr_buffer_32_1 f674(.wen(f674_wen), .wdata(f674_wdata), .clk(f674_clk), .rst(f674_rst), .rdata(f674_rdata));
  assign f674_clk = clk;
  assign f674_rst = rst;
  // Bindings to f674

  // f676
  logic [0:0] f676_wen;
  logic [31:0] f676_wdata;
  logic [0:0] f676_clk;
  logic [0:0] f676_rst;
  logic [31:0] f676_rdata;
  sr_buffer_32_1 f676(.wen(f676_wen), .wdata(f676_wdata), .clk(f676_clk), .rst(f676_rst), .rdata(f676_rdata));
  assign f676_clk = clk;
  assign f676_rst = rst;
  // Bindings to f676

  // f678
  logic [0:0] f678_wen;
  logic [31:0] f678_wdata;
  logic [0:0] f678_clk;
  logic [0:0] f678_rst;
  logic [31:0] f678_rdata;
  sr_buffer_32_1 f678(.wen(f678_wen), .wdata(f678_wdata), .clk(f678_clk), .rst(f678_rst), .rdata(f678_rdata));
  assign f678_clk = clk;
  assign f678_rst = rst;
  // Bindings to f678

  // f680
  logic [0:0] f680_wen;
  logic [31:0] f680_wdata;
  logic [0:0] f680_clk;
  logic [0:0] f680_rst;
  logic [31:0] f680_rdata;
  sr_buffer_32_1 f680(.wen(f680_wen), .wdata(f680_wdata), .clk(f680_clk), .rst(f680_rst), .rdata(f680_rdata));
  assign f680_clk = clk;
  assign f680_rst = rst;
  // Bindings to f680

  // f682
  logic [0:0] f682_wen;
  logic [31:0] f682_wdata;
  logic [0:0] f682_clk;
  logic [0:0] f682_rst;
  logic [31:0] f682_rdata;
  sr_buffer_32_1 f682(.wen(f682_wen), .wdata(f682_wdata), .clk(f682_clk), .rst(f682_rst), .rdata(f682_rdata));
  assign f682_clk = clk;
  assign f682_rst = rst;
  // Bindings to f682

  // f684
  logic [0:0] f684_wen;
  logic [31:0] f684_wdata;
  logic [0:0] f684_clk;
  logic [0:0] f684_rst;
  logic [31:0] f684_rdata;
  sr_buffer_32_1 f684(.wen(f684_wen), .wdata(f684_wdata), .clk(f684_clk), .rst(f684_rst), .rdata(f684_rdata));
  assign f684_clk = clk;
  assign f684_rst = rst;
  // Bindings to f684

  // f686
  logic [0:0] f686_wen;
  logic [31:0] f686_wdata;
  logic [0:0] f686_clk;
  logic [0:0] f686_rst;
  logic [31:0] f686_rdata;
  sr_buffer_32_1 f686(.wen(f686_wen), .wdata(f686_wdata), .clk(f686_clk), .rst(f686_rst), .rdata(f686_rdata));
  assign f686_clk = clk;
  assign f686_rst = rst;
  // Bindings to f686

  // f688
  logic [0:0] f688_wen;
  logic [31:0] f688_wdata;
  logic [0:0] f688_clk;
  logic [0:0] f688_rst;
  logic [31:0] f688_rdata;
  sr_buffer_32_1 f688(.wen(f688_wen), .wdata(f688_wdata), .clk(f688_clk), .rst(f688_rst), .rdata(f688_rdata));
  assign f688_clk = clk;
  assign f688_rst = rst;
  // Bindings to f688

  // f690
  logic [0:0] f690_wen;
  logic [31:0] f690_wdata;
  logic [0:0] f690_clk;
  logic [0:0] f690_rst;
  logic [31:0] f690_rdata;
  sr_buffer_32_1 f690(.wen(f690_wen), .wdata(f690_wdata), .clk(f690_clk), .rst(f690_rst), .rdata(f690_rdata));
  assign f690_clk = clk;
  assign f690_rst = rst;
  // Bindings to f690

  // f692
  logic [0:0] f692_wen;
  logic [31:0] f692_wdata;
  logic [0:0] f692_clk;
  logic [0:0] f692_rst;
  logic [31:0] f692_rdata;
  sr_buffer_32_1 f692(.wen(f692_wen), .wdata(f692_wdata), .clk(f692_clk), .rst(f692_rst), .rdata(f692_rdata));
  assign f692_clk = clk;
  assign f692_rst = rst;
  // Bindings to f692

  // f694
  logic [0:0] f694_wen;
  logic [31:0] f694_wdata;
  logic [0:0] f694_clk;
  logic [0:0] f694_rst;
  logic [31:0] f694_rdata;
  sr_buffer_32_1 f694(.wen(f694_wen), .wdata(f694_wdata), .clk(f694_clk), .rst(f694_rst), .rdata(f694_rdata));
  assign f694_clk = clk;
  assign f694_rst = rst;
  // Bindings to f694

  // f696
  logic [0:0] f696_wen;
  logic [31:0] f696_wdata;
  logic [0:0] f696_clk;
  logic [0:0] f696_rst;
  logic [31:0] f696_rdata;
  sr_buffer_32_1 f696(.wen(f696_wen), .wdata(f696_wdata), .clk(f696_clk), .rst(f696_rst), .rdata(f696_rdata));
  assign f696_clk = clk;
  assign f696_rst = rst;
  // Bindings to f696

  // f698
  logic [0:0] f698_wen;
  logic [31:0] f698_wdata;
  logic [0:0] f698_clk;
  logic [0:0] f698_rst;
  logic [31:0] f698_rdata;
  sr_buffer_32_1 f698(.wen(f698_wen), .wdata(f698_wdata), .clk(f698_clk), .rst(f698_rst), .rdata(f698_rdata));
  assign f698_clk = clk;
  assign f698_rst = rst;
  // Bindings to f698

  // f700
  logic [0:0] f700_wen;
  logic [31:0] f700_wdata;
  logic [0:0] f700_clk;
  logic [0:0] f700_rst;
  logic [31:0] f700_rdata;
  sr_buffer_32_1 f700(.wen(f700_wen), .wdata(f700_wdata), .clk(f700_clk), .rst(f700_rst), .rdata(f700_rdata));
  assign f700_clk = clk;
  assign f700_rst = rst;
  // Bindings to f700

  // f702
  logic [0:0] f702_wen;
  logic [31:0] f702_wdata;
  logic [0:0] f702_clk;
  logic [0:0] f702_rst;
  logic [31:0] f702_rdata;
  sr_buffer_32_1 f702(.wen(f702_wen), .wdata(f702_wdata), .clk(f702_clk), .rst(f702_rst), .rdata(f702_rdata));
  assign f702_clk = clk;
  assign f702_rst = rst;
  // Bindings to f702

  // f704
  logic [0:0] f704_wen;
  logic [31:0] f704_wdata;
  logic [0:0] f704_clk;
  logic [0:0] f704_rst;
  logic [31:0] f704_rdata;
  sr_buffer_32_1 f704(.wen(f704_wen), .wdata(f704_wdata), .clk(f704_clk), .rst(f704_rst), .rdata(f704_rdata));
  assign f704_clk = clk;
  assign f704_rst = rst;
  // Bindings to f704

  // f706
  logic [0:0] f706_wen;
  logic [31:0] f706_wdata;
  logic [0:0] f706_clk;
  logic [0:0] f706_rst;
  logic [31:0] f706_rdata;
  sr_buffer_32_1 f706(.wen(f706_wen), .wdata(f706_wdata), .clk(f706_clk), .rst(f706_rst), .rdata(f706_rdata));
  assign f706_clk = clk;
  assign f706_rst = rst;
  // Bindings to f706

  // f708
  logic [0:0] f708_wen;
  logic [31:0] f708_wdata;
  logic [0:0] f708_clk;
  logic [0:0] f708_rst;
  logic [31:0] f708_rdata;
  sr_buffer_32_1 f708(.wen(f708_wen), .wdata(f708_wdata), .clk(f708_clk), .rst(f708_rst), .rdata(f708_rdata));
  assign f708_clk = clk;
  assign f708_rst = rst;
  // Bindings to f708

  // f710
  logic [0:0] f710_wen;
  logic [31:0] f710_wdata;
  logic [0:0] f710_clk;
  logic [0:0] f710_rst;
  logic [31:0] f710_rdata;
  sr_buffer_32_1 f710(.wen(f710_wen), .wdata(f710_wdata), .clk(f710_clk), .rst(f710_rst), .rdata(f710_rdata));
  assign f710_clk = clk;
  assign f710_rst = rst;
  // Bindings to f710

  // f712
  logic [0:0] f712_wen;
  logic [31:0] f712_wdata;
  logic [0:0] f712_clk;
  logic [0:0] f712_rst;
  logic [31:0] f712_rdata;
  sr_buffer_32_1 f712(.wen(f712_wen), .wdata(f712_wdata), .clk(f712_clk), .rst(f712_rst), .rdata(f712_rdata));
  assign f712_clk = clk;
  assign f712_rst = rst;
  // Bindings to f712

  // f714
  logic [0:0] f714_wen;
  logic [31:0] f714_wdata;
  logic [0:0] f714_clk;
  logic [0:0] f714_rst;
  logic [31:0] f714_rdata;
  sr_buffer_32_1 f714(.wen(f714_wen), .wdata(f714_wdata), .clk(f714_clk), .rst(f714_rst), .rdata(f714_rdata));
  assign f714_clk = clk;
  assign f714_rst = rst;
  // Bindings to f714

  // f716
  logic [0:0] f716_wen;
  logic [31:0] f716_wdata;
  logic [0:0] f716_clk;
  logic [0:0] f716_rst;
  logic [31:0] f716_rdata;
  sr_buffer_32_1 f716(.wen(f716_wen), .wdata(f716_wdata), .clk(f716_clk), .rst(f716_rst), .rdata(f716_rdata));
  assign f716_clk = clk;
  assign f716_rst = rst;
  // Bindings to f716

  // f718
  logic [0:0] f718_wen;
  logic [31:0] f718_wdata;
  logic [0:0] f718_clk;
  logic [0:0] f718_rst;
  logic [31:0] f718_rdata;
  sr_buffer_32_1 f718(.wen(f718_wen), .wdata(f718_wdata), .clk(f718_clk), .rst(f718_rst), .rdata(f718_rdata));
  assign f718_clk = clk;
  assign f718_rst = rst;
  // Bindings to f718

  // f720
  logic [0:0] f720_wen;
  logic [31:0] f720_wdata;
  logic [0:0] f720_clk;
  logic [0:0] f720_rst;
  logic [31:0] f720_rdata;
  sr_buffer_32_1 f720(.wen(f720_wen), .wdata(f720_wdata), .clk(f720_clk), .rst(f720_rst), .rdata(f720_rdata));
  assign f720_clk = clk;
  assign f720_rst = rst;
  // Bindings to f720

  // f722
  logic [0:0] f722_wen;
  logic [31:0] f722_wdata;
  logic [0:0] f722_clk;
  logic [0:0] f722_rst;
  logic [31:0] f722_rdata;
  sr_buffer_32_1 f722(.wen(f722_wen), .wdata(f722_wdata), .clk(f722_clk), .rst(f722_rst), .rdata(f722_rdata));
  assign f722_clk = clk;
  assign f722_rst = rst;
  // Bindings to f722

  // f724
  logic [0:0] f724_wen;
  logic [31:0] f724_wdata;
  logic [0:0] f724_clk;
  logic [0:0] f724_rst;
  logic [31:0] f724_rdata;
  sr_buffer_32_1 f724(.wen(f724_wen), .wdata(f724_wdata), .clk(f724_clk), .rst(f724_rst), .rdata(f724_rdata));
  assign f724_clk = clk;
  assign f724_rst = rst;
  // Bindings to f724

  // f726
  logic [0:0] f726_wen;
  logic [31:0] f726_wdata;
  logic [0:0] f726_clk;
  logic [0:0] f726_rst;
  logic [31:0] f726_rdata;
  sr_buffer_32_1 f726(.wen(f726_wen), .wdata(f726_wdata), .clk(f726_clk), .rst(f726_rst), .rdata(f726_rdata));
  assign f726_clk = clk;
  assign f726_rst = rst;
  // Bindings to f726

  // f728
  logic [0:0] f728_wen;
  logic [31:0] f728_wdata;
  logic [0:0] f728_clk;
  logic [0:0] f728_rst;
  logic [31:0] f728_rdata;
  sr_buffer_32_1 f728(.wen(f728_wen), .wdata(f728_wdata), .clk(f728_clk), .rst(f728_rst), .rdata(f728_rdata));
  assign f728_clk = clk;
  assign f728_rst = rst;
  // Bindings to f728

  // f730
  logic [0:0] f730_wen;
  logic [31:0] f730_wdata;
  logic [0:0] f730_clk;
  logic [0:0] f730_rst;
  logic [31:0] f730_rdata;
  sr_buffer_32_1 f730(.wen(f730_wen), .wdata(f730_wdata), .clk(f730_clk), .rst(f730_rst), .rdata(f730_rdata));
  assign f730_clk = clk;
  assign f730_rst = rst;
  // Bindings to f730

  // f732
  logic [0:0] f732_wen;
  logic [31:0] f732_wdata;
  logic [0:0] f732_clk;
  logic [0:0] f732_rst;
  logic [31:0] f732_rdata;
  sr_buffer_32_1 f732(.wen(f732_wen), .wdata(f732_wdata), .clk(f732_clk), .rst(f732_rst), .rdata(f732_rdata));
  assign f732_clk = clk;
  assign f732_rst = rst;
  // Bindings to f732

  // f734
  logic [0:0] f734_wen;
  logic [31:0] f734_wdata;
  logic [0:0] f734_clk;
  logic [0:0] f734_rst;
  logic [31:0] f734_rdata;
  sr_buffer_32_1 f734(.wen(f734_wen), .wdata(f734_wdata), .clk(f734_clk), .rst(f734_rst), .rdata(f734_rdata));
  assign f734_clk = clk;
  assign f734_rst = rst;
  // Bindings to f734

  // f736
  logic [0:0] f736_wen;
  logic [31:0] f736_wdata;
  logic [0:0] f736_clk;
  logic [0:0] f736_rst;
  logic [31:0] f736_rdata;
  sr_buffer_32_1 f736(.wen(f736_wen), .wdata(f736_wdata), .clk(f736_clk), .rst(f736_rst), .rdata(f736_rdata));
  assign f736_clk = clk;
  assign f736_rst = rst;
  // Bindings to f736

  // f738
  logic [0:0] f738_wen;
  logic [31:0] f738_wdata;
  logic [0:0] f738_clk;
  logic [0:0] f738_rst;
  logic [31:0] f738_rdata;
  sr_buffer_32_1 f738(.wen(f738_wen), .wdata(f738_wdata), .clk(f738_clk), .rst(f738_rst), .rdata(f738_rdata));
  assign f738_clk = clk;
  assign f738_rst = rst;
  // Bindings to f738

  // f740
  logic [0:0] f740_wen;
  logic [31:0] f740_wdata;
  logic [0:0] f740_clk;
  logic [0:0] f740_rst;
  logic [31:0] f740_rdata;
  sr_buffer_32_1 f740(.wen(f740_wen), .wdata(f740_wdata), .clk(f740_clk), .rst(f740_rst), .rdata(f740_rdata));
  assign f740_clk = clk;
  assign f740_rst = rst;
  // Bindings to f740

  // f742
  logic [0:0] f742_wen;
  logic [31:0] f742_wdata;
  logic [0:0] f742_clk;
  logic [0:0] f742_rst;
  logic [31:0] f742_rdata;
  sr_buffer_32_1 f742(.wen(f742_wen), .wdata(f742_wdata), .clk(f742_clk), .rst(f742_rst), .rdata(f742_rdata));
  assign f742_clk = clk;
  assign f742_rst = rst;
  // Bindings to f742

  // f744
  logic [0:0] f744_wen;
  logic [31:0] f744_wdata;
  logic [0:0] f744_clk;
  logic [0:0] f744_rst;
  logic [31:0] f744_rdata;
  sr_buffer_32_1 f744(.wen(f744_wen), .wdata(f744_wdata), .clk(f744_clk), .rst(f744_rst), .rdata(f744_rdata));
  assign f744_clk = clk;
  assign f744_rst = rst;
  // Bindings to f744

  // f746
  logic [0:0] f746_wen;
  logic [31:0] f746_wdata;
  logic [0:0] f746_clk;
  logic [0:0] f746_rst;
  logic [31:0] f746_rdata;
  sr_buffer_32_1 f746(.wen(f746_wen), .wdata(f746_wdata), .clk(f746_clk), .rst(f746_rst), .rdata(f746_rdata));
  assign f746_clk = clk;
  assign f746_rst = rst;
  // Bindings to f746

  // f748
  logic [0:0] f748_wen;
  logic [31:0] f748_wdata;
  logic [0:0] f748_clk;
  logic [0:0] f748_rst;
  logic [31:0] f748_rdata;
  sr_buffer_32_1 f748(.wen(f748_wen), .wdata(f748_wdata), .clk(f748_clk), .rst(f748_rst), .rdata(f748_rdata));
  assign f748_clk = clk;
  assign f748_rst = rst;
  // Bindings to f748

  // f750
  logic [0:0] f750_wen;
  logic [31:0] f750_wdata;
  logic [0:0] f750_clk;
  logic [0:0] f750_rst;
  logic [31:0] f750_rdata;
  sr_buffer_32_1 f750(.wen(f750_wen), .wdata(f750_wdata), .clk(f750_clk), .rst(f750_rst), .rdata(f750_rdata));
  assign f750_clk = clk;
  assign f750_rst = rst;
  // Bindings to f750

  // f752
  logic [0:0] f752_wen;
  logic [31:0] f752_wdata;
  logic [0:0] f752_clk;
  logic [0:0] f752_rst;
  logic [31:0] f752_rdata;
  sr_buffer_32_1 f752(.wen(f752_wen), .wdata(f752_wdata), .clk(f752_clk), .rst(f752_rst), .rdata(f752_rdata));
  assign f752_clk = clk;
  assign f752_rst = rst;
  // Bindings to f752

  // f754
  logic [0:0] f754_wen;
  logic [31:0] f754_wdata;
  logic [0:0] f754_clk;
  logic [0:0] f754_rst;
  logic [31:0] f754_rdata;
  sr_buffer_32_1 f754(.wen(f754_wen), .wdata(f754_wdata), .clk(f754_clk), .rst(f754_rst), .rdata(f754_rdata));
  assign f754_clk = clk;
  assign f754_rst = rst;
  // Bindings to f754

  // f756
  logic [0:0] f756_wen;
  logic [31:0] f756_wdata;
  logic [0:0] f756_clk;
  logic [0:0] f756_rst;
  logic [31:0] f756_rdata;
  sr_buffer_32_1 f756(.wen(f756_wen), .wdata(f756_wdata), .clk(f756_clk), .rst(f756_rst), .rdata(f756_rdata));
  assign f756_clk = clk;
  assign f756_rst = rst;
  // Bindings to f756

  // f758
  logic [0:0] f758_wen;
  logic [31:0] f758_wdata;
  logic [0:0] f758_clk;
  logic [0:0] f758_rst;
  logic [31:0] f758_rdata;
  sr_buffer_32_1 f758(.wen(f758_wen), .wdata(f758_wdata), .clk(f758_clk), .rst(f758_rst), .rdata(f758_rdata));
  assign f758_clk = clk;
  assign f758_rst = rst;
  // Bindings to f758

  // f760
  logic [0:0] f760_wen;
  logic [31:0] f760_wdata;
  logic [0:0] f760_clk;
  logic [0:0] f760_rst;
  logic [31:0] f760_rdata;
  sr_buffer_32_1 f760(.wen(f760_wen), .wdata(f760_wdata), .clk(f760_clk), .rst(f760_rst), .rdata(f760_rdata));
  assign f760_clk = clk;
  assign f760_rst = rst;
  // Bindings to f760

  // f762
  logic [0:0] f762_wen;
  logic [31:0] f762_wdata;
  logic [0:0] f762_clk;
  logic [0:0] f762_rst;
  logic [31:0] f762_rdata;
  sr_buffer_32_1 f762(.wen(f762_wen), .wdata(f762_wdata), .clk(f762_clk), .rst(f762_rst), .rdata(f762_rdata));
  assign f762_clk = clk;
  assign f762_rst = rst;
  // Bindings to f762

  // f764
  logic [0:0] f764_wen;
  logic [31:0] f764_wdata;
  logic [0:0] f764_clk;
  logic [0:0] f764_rst;
  logic [31:0] f764_rdata;
  sr_buffer_32_1 f764(.wen(f764_wen), .wdata(f764_wdata), .clk(f764_clk), .rst(f764_rst), .rdata(f764_rdata));
  assign f764_clk = clk;
  assign f764_rst = rst;
  // Bindings to f764

  // f766
  logic [0:0] f766_wen;
  logic [31:0] f766_wdata;
  logic [0:0] f766_clk;
  logic [0:0] f766_rst;
  logic [31:0] f766_rdata;
  sr_buffer_32_1 f766(.wen(f766_wen), .wdata(f766_wdata), .clk(f766_clk), .rst(f766_rst), .rdata(f766_rdata));
  assign f766_clk = clk;
  assign f766_rst = rst;
  // Bindings to f766

  // f768
  logic [0:0] f768_wen;
  logic [31:0] f768_wdata;
  logic [0:0] f768_clk;
  logic [0:0] f768_rst;
  logic [31:0] f768_rdata;
  sr_buffer_32_1 f768(.wen(f768_wen), .wdata(f768_wdata), .clk(f768_clk), .rst(f768_rst), .rdata(f768_rdata));
  assign f768_clk = clk;
  assign f768_rst = rst;
  // Bindings to f768

  // f770
  logic [0:0] f770_wen;
  logic [31:0] f770_wdata;
  logic [0:0] f770_clk;
  logic [0:0] f770_rst;
  logic [31:0] f770_rdata;
  sr_buffer_32_1 f770(.wen(f770_wen), .wdata(f770_wdata), .clk(f770_clk), .rst(f770_rst), .rdata(f770_rdata));
  assign f770_clk = clk;
  assign f770_rst = rst;
  // Bindings to f770

  // f1034
  logic [0:0] f1034_wen;
  logic [31:0] f1034_wdata;
  logic [0:0] f1034_clk;
  logic [0:0] f1034_rst;
  logic [31:0] f1034_rdata;
  sr_buffer_32_1 f1034(.wen(f1034_wen), .wdata(f1034_wdata), .clk(f1034_clk), .rst(f1034_rst), .rdata(f1034_rdata));
  assign f1034_clk = clk;
  assign f1034_rst = rst;
  // Bindings to f1034

  // f1026
  logic [0:0] f1026_wen;
  logic [31:0] f1026_wdata;
  logic [0:0] f1026_clk;
  logic [0:0] f1026_rst;
  logic [31:0] f1026_rdata;
  sr_buffer_32_1 f1026(.wen(f1026_wen), .wdata(f1026_wdata), .clk(f1026_clk), .rst(f1026_rst), .rdata(f1026_rdata));
  assign f1026_clk = clk;
  assign f1026_rst = rst;
  // Bindings to f1026

  // f1020
  logic [0:0] f1020_wen;
  logic [31:0] f1020_wdata;
  logic [0:0] f1020_clk;
  logic [0:0] f1020_rst;
  logic [31:0] f1020_rdata;
  sr_buffer_32_1 f1020(.wen(f1020_wen), .wdata(f1020_wdata), .clk(f1020_clk), .rst(f1020_rst), .rdata(f1020_rdata));
  assign f1020_clk = clk;
  assign f1020_rst = rst;
  // Bindings to f1020

  // f1006
  logic [0:0] f1006_wen;
  logic [31:0] f1006_wdata;
  logic [0:0] f1006_clk;
  logic [0:0] f1006_rst;
  logic [31:0] f1006_rdata;
  sr_buffer_32_1 f1006(.wen(f1006_wen), .wdata(f1006_wdata), .clk(f1006_clk), .rst(f1006_rst), .rdata(f1006_rdata));
  assign f1006_clk = clk;
  assign f1006_rst = rst;
  // Bindings to f1006

  // f970
  logic [0:0] f970_wen;
  logic [31:0] f970_wdata;
  logic [0:0] f970_clk;
  logic [0:0] f970_rst;
  logic [31:0] f970_rdata;
  sr_buffer_32_1 f970(.wen(f970_wen), .wdata(f970_wdata), .clk(f970_clk), .rst(f970_rst), .rdata(f970_rdata));
  assign f970_clk = clk;
  assign f970_rst = rst;
  // Bindings to f970

  // f1032
  logic [0:0] f1032_wen;
  logic [31:0] f1032_wdata;
  logic [0:0] f1032_clk;
  logic [0:0] f1032_rst;
  logic [31:0] f1032_rdata;
  sr_buffer_32_1 f1032(.wen(f1032_wen), .wdata(f1032_wdata), .clk(f1032_clk), .rst(f1032_rst), .rdata(f1032_rdata));
  assign f1032_clk = clk;
  assign f1032_rst = rst;
  // Bindings to f1032

  // f1030
  logic [0:0] f1030_wen;
  logic [31:0] f1030_wdata;
  logic [0:0] f1030_clk;
  logic [0:0] f1030_rst;
  logic [31:0] f1030_rdata;
  sr_buffer_32_1 f1030(.wen(f1030_wen), .wdata(f1030_wdata), .clk(f1030_clk), .rst(f1030_rst), .rdata(f1030_rdata));
  assign f1030_clk = clk;
  assign f1030_rst = rst;
  // Bindings to f1030

  // f1028
  logic [0:0] f1028_wen;
  logic [31:0] f1028_wdata;
  logic [0:0] f1028_clk;
  logic [0:0] f1028_rst;
  logic [31:0] f1028_rdata;
  sr_buffer_32_1 f1028(.wen(f1028_wen), .wdata(f1028_wdata), .clk(f1028_clk), .rst(f1028_rst), .rdata(f1028_rdata));
  assign f1028_clk = clk;
  assign f1028_rst = rst;
  // Bindings to f1028

  // f1022
  logic [0:0] f1022_wen;
  logic [31:0] f1022_wdata;
  logic [0:0] f1022_clk;
  logic [0:0] f1022_rst;
  logic [31:0] f1022_rdata;
  sr_buffer_32_1 f1022(.wen(f1022_wen), .wdata(f1022_wdata), .clk(f1022_clk), .rst(f1022_rst), .rdata(f1022_rdata));
  assign f1022_clk = clk;
  assign f1022_rst = rst;
  // Bindings to f1022

  // f1024
  logic [0:0] f1024_wen;
  logic [31:0] f1024_wdata;
  logic [0:0] f1024_clk;
  logic [0:0] f1024_rst;
  logic [31:0] f1024_rdata;
  sr_buffer_32_1 f1024(.wen(f1024_wen), .wdata(f1024_wdata), .clk(f1024_clk), .rst(f1024_rst), .rdata(f1024_rdata));
  assign f1024_clk = clk;
  assign f1024_rst = rst;
  // Bindings to f1024

  // f1018
  logic [0:0] f1018_wen;
  logic [31:0] f1018_wdata;
  logic [0:0] f1018_clk;
  logic [0:0] f1018_rst;
  logic [31:0] f1018_rdata;
  sr_buffer_32_1 f1018(.wen(f1018_wen), .wdata(f1018_wdata), .clk(f1018_clk), .rst(f1018_rst), .rdata(f1018_rdata));
  assign f1018_clk = clk;
  assign f1018_rst = rst;
  // Bindings to f1018

  // f1010
  logic [0:0] f1010_wen;
  logic [31:0] f1010_wdata;
  logic [0:0] f1010_clk;
  logic [0:0] f1010_rst;
  logic [31:0] f1010_rdata;
  sr_buffer_32_1 f1010(.wen(f1010_wen), .wdata(f1010_wdata), .clk(f1010_clk), .rst(f1010_rst), .rdata(f1010_rdata));
  assign f1010_clk = clk;
  assign f1010_rst = rst;
  // Bindings to f1010

  // f1016
  logic [0:0] f1016_wen;
  logic [31:0] f1016_wdata;
  logic [0:0] f1016_clk;
  logic [0:0] f1016_rst;
  logic [31:0] f1016_rdata;
  sr_buffer_32_1 f1016(.wen(f1016_wen), .wdata(f1016_wdata), .clk(f1016_clk), .rst(f1016_rst), .rdata(f1016_rdata));
  assign f1016_clk = clk;
  assign f1016_rst = rst;
  // Bindings to f1016

  // f1014
  logic [0:0] f1014_wen;
  logic [31:0] f1014_wdata;
  logic [0:0] f1014_clk;
  logic [0:0] f1014_rst;
  logic [31:0] f1014_rdata;
  sr_buffer_32_1 f1014(.wen(f1014_wen), .wdata(f1014_wdata), .clk(f1014_clk), .rst(f1014_rst), .rdata(f1014_rdata));
  assign f1014_clk = clk;
  assign f1014_rst = rst;
  // Bindings to f1014

  // f1012
  logic [0:0] f1012_wen;
  logic [31:0] f1012_wdata;
  logic [0:0] f1012_clk;
  logic [0:0] f1012_rst;
  logic [31:0] f1012_rdata;
  sr_buffer_32_1 f1012(.wen(f1012_wen), .wdata(f1012_wdata), .clk(f1012_clk), .rst(f1012_rst), .rdata(f1012_rdata));
  assign f1012_clk = clk;
  assign f1012_rst = rst;
  // Bindings to f1012

  // f1008
  logic [0:0] f1008_wen;
  logic [31:0] f1008_wdata;
  logic [0:0] f1008_clk;
  logic [0:0] f1008_rst;
  logic [31:0] f1008_rdata;
  sr_buffer_32_1 f1008(.wen(f1008_wen), .wdata(f1008_wdata), .clk(f1008_clk), .rst(f1008_rst), .rdata(f1008_rdata));
  assign f1008_clk = clk;
  assign f1008_rst = rst;
  // Bindings to f1008

  // f994
  logic [0:0] f994_wen;
  logic [31:0] f994_wdata;
  logic [0:0] f994_clk;
  logic [0:0] f994_rst;
  logic [31:0] f994_rdata;
  sr_buffer_32_1 f994(.wen(f994_wen), .wdata(f994_wdata), .clk(f994_clk), .rst(f994_rst), .rdata(f994_rdata));
  assign f994_clk = clk;
  assign f994_rst = rst;
  // Bindings to f994

  // f996
  logic [0:0] f996_wen;
  logic [31:0] f996_wdata;
  logic [0:0] f996_clk;
  logic [0:0] f996_rst;
  logic [31:0] f996_rdata;
  sr_buffer_32_1 f996(.wen(f996_wen), .wdata(f996_wdata), .clk(f996_clk), .rst(f996_rst), .rdata(f996_rdata));
  assign f996_clk = clk;
  assign f996_rst = rst;
  // Bindings to f996

  // f998
  logic [0:0] f998_wen;
  logic [31:0] f998_wdata;
  logic [0:0] f998_clk;
  logic [0:0] f998_rst;
  logic [31:0] f998_rdata;
  sr_buffer_32_1 f998(.wen(f998_wen), .wdata(f998_wdata), .clk(f998_clk), .rst(f998_rst), .rdata(f998_rdata));
  assign f998_clk = clk;
  assign f998_rst = rst;
  // Bindings to f998

  // f1004
  logic [0:0] f1004_wen;
  logic [31:0] f1004_wdata;
  logic [0:0] f1004_clk;
  logic [0:0] f1004_rst;
  logic [31:0] f1004_rdata;
  sr_buffer_32_1 f1004(.wen(f1004_wen), .wdata(f1004_wdata), .clk(f1004_clk), .rst(f1004_rst), .rdata(f1004_rdata));
  assign f1004_clk = clk;
  assign f1004_rst = rst;
  // Bindings to f1004

  // f966
  logic [0:0] f966_wen;
  logic [31:0] f966_wdata;
  logic [0:0] f966_clk;
  logic [0:0] f966_rst;
  logic [31:0] f966_rdata;
  sr_buffer_32_1 f966(.wen(f966_wen), .wdata(f966_wdata), .clk(f966_clk), .rst(f966_rst), .rdata(f966_rdata));
  assign f966_clk = clk;
  assign f966_rst = rst;
  // Bindings to f966

  // f1000
  logic [0:0] f1000_wen;
  logic [31:0] f1000_wdata;
  logic [0:0] f1000_clk;
  logic [0:0] f1000_rst;
  logic [31:0] f1000_rdata;
  sr_buffer_32_1 f1000(.wen(f1000_wen), .wdata(f1000_wdata), .clk(f1000_clk), .rst(f1000_rst), .rdata(f1000_rdata));
  assign f1000_clk = clk;
  assign f1000_rst = rst;
  // Bindings to f1000

  // f964
  logic [0:0] f964_wen;
  logic [31:0] f964_wdata;
  logic [0:0] f964_clk;
  logic [0:0] f964_rst;
  logic [31:0] f964_rdata;
  sr_buffer_32_1 f964(.wen(f964_wen), .wdata(f964_wdata), .clk(f964_clk), .rst(f964_rst), .rdata(f964_rdata));
  assign f964_clk = clk;
  assign f964_rst = rst;
  // Bindings to f964

  // f968
  logic [0:0] f968_wen;
  logic [31:0] f968_wdata;
  logic [0:0] f968_clk;
  logic [0:0] f968_rst;
  logic [31:0] f968_rdata;
  sr_buffer_32_1 f968(.wen(f968_wen), .wdata(f968_wdata), .clk(f968_clk), .rst(f968_rst), .rdata(f968_rdata));
  assign f968_clk = clk;
  assign f968_rst = rst;
  // Bindings to f968

  // f978
  logic [0:0] f978_wen;
  logic [31:0] f978_wdata;
  logic [0:0] f978_clk;
  logic [0:0] f978_rst;
  logic [31:0] f978_rdata;
  sr_buffer_32_1 f978(.wen(f978_wen), .wdata(f978_wdata), .clk(f978_clk), .rst(f978_rst), .rdata(f978_rdata));
  assign f978_clk = clk;
  assign f978_rst = rst;
  // Bindings to f978

  // f984
  logic [0:0] f984_wen;
  logic [31:0] f984_wdata;
  logic [0:0] f984_clk;
  logic [0:0] f984_rst;
  logic [31:0] f984_rdata;
  sr_buffer_32_1 f984(.wen(f984_wen), .wdata(f984_wdata), .clk(f984_clk), .rst(f984_rst), .rdata(f984_rdata));
  assign f984_clk = clk;
  assign f984_rst = rst;
  // Bindings to f984

  // f982
  logic [0:0] f982_wen;
  logic [31:0] f982_wdata;
  logic [0:0] f982_clk;
  logic [0:0] f982_rst;
  logic [31:0] f982_rdata;
  sr_buffer_32_1 f982(.wen(f982_wen), .wdata(f982_wdata), .clk(f982_clk), .rst(f982_rst), .rdata(f982_rdata));
  assign f982_clk = clk;
  assign f982_rst = rst;
  // Bindings to f982

  // f972
  logic [0:0] f972_wen;
  logic [31:0] f972_wdata;
  logic [0:0] f972_clk;
  logic [0:0] f972_rst;
  logic [31:0] f972_rdata;
  sr_buffer_32_1 f972(.wen(f972_wen), .wdata(f972_wdata), .clk(f972_clk), .rst(f972_rst), .rdata(f972_rdata));
  assign f972_clk = clk;
  assign f972_rst = rst;
  // Bindings to f972

  // f990
  logic [0:0] f990_wen;
  logic [31:0] f990_wdata;
  logic [0:0] f990_clk;
  logic [0:0] f990_rst;
  logic [31:0] f990_rdata;
  sr_buffer_32_1 f990(.wen(f990_wen), .wdata(f990_wdata), .clk(f990_clk), .rst(f990_rst), .rdata(f990_rdata));
  assign f990_clk = clk;
  assign f990_rst = rst;
  // Bindings to f990

  // f1002
  logic [0:0] f1002_wen;
  logic [31:0] f1002_wdata;
  logic [0:0] f1002_clk;
  logic [0:0] f1002_rst;
  logic [31:0] f1002_rdata;
  sr_buffer_32_1 f1002(.wen(f1002_wen), .wdata(f1002_wdata), .clk(f1002_clk), .rst(f1002_rst), .rdata(f1002_rdata));
  assign f1002_clk = clk;
  assign f1002_rst = rst;
  // Bindings to f1002

  // f976
  logic [0:0] f976_wen;
  logic [31:0] f976_wdata;
  logic [0:0] f976_clk;
  logic [0:0] f976_rst;
  logic [31:0] f976_rdata;
  sr_buffer_32_1 f976(.wen(f976_wen), .wdata(f976_wdata), .clk(f976_clk), .rst(f976_rst), .rdata(f976_rdata));
  assign f976_clk = clk;
  assign f976_rst = rst;
  // Bindings to f976

  // f974
  logic [0:0] f974_wen;
  logic [31:0] f974_wdata;
  logic [0:0] f974_clk;
  logic [0:0] f974_rst;
  logic [31:0] f974_rdata;
  sr_buffer_32_1 f974(.wen(f974_wen), .wdata(f974_wdata), .clk(f974_clk), .rst(f974_rst), .rdata(f974_rdata));
  assign f974_clk = clk;
  assign f974_rst = rst;
  // Bindings to f974

  // f992
  logic [0:0] f992_wen;
  logic [31:0] f992_wdata;
  logic [0:0] f992_clk;
  logic [0:0] f992_rst;
  logic [31:0] f992_rdata;
  sr_buffer_32_1 f992(.wen(f992_wen), .wdata(f992_wdata), .clk(f992_clk), .rst(f992_rst), .rdata(f992_rdata));
  assign f992_clk = clk;
  assign f992_rst = rst;
  // Bindings to f992

  // f986
  logic [0:0] f986_wen;
  logic [31:0] f986_wdata;
  logic [0:0] f986_clk;
  logic [0:0] f986_rst;
  logic [31:0] f986_rdata;
  sr_buffer_32_1 f986(.wen(f986_wen), .wdata(f986_wdata), .clk(f986_clk), .rst(f986_rst), .rdata(f986_rdata));
  assign f986_clk = clk;
  assign f986_rst = rst;
  // Bindings to f986

  // f988
  logic [0:0] f988_wen;
  logic [31:0] f988_wdata;
  logic [0:0] f988_clk;
  logic [0:0] f988_rst;
  logic [31:0] f988_rdata;
  sr_buffer_32_1 f988(.wen(f988_wen), .wdata(f988_wdata), .clk(f988_clk), .rst(f988_rst), .rdata(f988_rdata));
  assign f988_clk = clk;
  assign f988_rst = rst;
  // Bindings to f988

  // f962
  logic [0:0] f962_wen;
  logic [31:0] f962_wdata;
  logic [0:0] f962_clk;
  logic [0:0] f962_rst;
  logic [31:0] f962_rdata;
  sr_buffer_32_1 f962(.wen(f962_wen), .wdata(f962_wdata), .clk(f962_clk), .rst(f962_rst), .rdata(f962_rdata));
  assign f962_clk = clk;
  assign f962_rst = rst;
  // Bindings to f962

  // f1036
  logic [0:0] f1036_wen;
  logic [31:0] f1036_wdata;
  logic [0:0] f1036_clk;
  logic [0:0] f1036_rst;
  logic [31:0] f1036_rdata;
  sr_buffer_32_1 f1036(.wen(f1036_wen), .wdata(f1036_wdata), .clk(f1036_clk), .rst(f1036_rst), .rdata(f1036_rdata));
  assign f1036_clk = clk;
  assign f1036_rst = rst;
  // Bindings to f1036

  // f1038
  logic [0:0] f1038_wen;
  logic [31:0] f1038_wdata;
  logic [0:0] f1038_clk;
  logic [0:0] f1038_rst;
  logic [31:0] f1038_rdata;
  sr_buffer_32_1 f1038(.wen(f1038_wen), .wdata(f1038_wdata), .clk(f1038_clk), .rst(f1038_rst), .rdata(f1038_rdata));
  assign f1038_clk = clk;
  assign f1038_rst = rst;
  // Bindings to f1038

  // f1040
  logic [0:0] f1040_wen;
  logic [31:0] f1040_wdata;
  logic [0:0] f1040_clk;
  logic [0:0] f1040_rst;
  logic [31:0] f1040_rdata;
  sr_buffer_32_1 f1040(.wen(f1040_wen), .wdata(f1040_wdata), .clk(f1040_clk), .rst(f1040_rst), .rdata(f1040_rdata));
  assign f1040_clk = clk;
  assign f1040_rst = rst;
  // Bindings to f1040

  // f1042
  logic [0:0] f1042_wen;
  logic [31:0] f1042_wdata;
  logic [0:0] f1042_clk;
  logic [0:0] f1042_rst;
  logic [31:0] f1042_rdata;
  sr_buffer_32_1 f1042(.wen(f1042_wen), .wdata(f1042_wdata), .clk(f1042_clk), .rst(f1042_rst), .rdata(f1042_rdata));
  assign f1042_clk = clk;
  assign f1042_rst = rst;
  // Bindings to f1042

  // f1044
  logic [0:0] f1044_wen;
  logic [31:0] f1044_wdata;
  logic [0:0] f1044_clk;
  logic [0:0] f1044_rst;
  logic [31:0] f1044_rdata;
  sr_buffer_32_1 f1044(.wen(f1044_wen), .wdata(f1044_wdata), .clk(f1044_clk), .rst(f1044_rst), .rdata(f1044_rdata));
  assign f1044_clk = clk;
  assign f1044_rst = rst;
  // Bindings to f1044

  // f1046
  logic [0:0] f1046_wen;
  logic [31:0] f1046_wdata;
  logic [0:0] f1046_clk;
  logic [0:0] f1046_rst;
  logic [31:0] f1046_rdata;
  sr_buffer_32_1 f1046(.wen(f1046_wen), .wdata(f1046_wdata), .clk(f1046_clk), .rst(f1046_rst), .rdata(f1046_rdata));
  assign f1046_clk = clk;
  assign f1046_rst = rst;
  // Bindings to f1046

  // f1048
  logic [0:0] f1048_wen;
  logic [31:0] f1048_wdata;
  logic [0:0] f1048_clk;
  logic [0:0] f1048_rst;
  logic [31:0] f1048_rdata;
  sr_buffer_32_1 f1048(.wen(f1048_wen), .wdata(f1048_wdata), .clk(f1048_clk), .rst(f1048_rst), .rdata(f1048_rdata));
  assign f1048_clk = clk;
  assign f1048_rst = rst;
  // Bindings to f1048

  // f1050
  logic [0:0] f1050_wen;
  logic [31:0] f1050_wdata;
  logic [0:0] f1050_clk;
  logic [0:0] f1050_rst;
  logic [31:0] f1050_rdata;
  sr_buffer_32_1 f1050(.wen(f1050_wen), .wdata(f1050_wdata), .clk(f1050_clk), .rst(f1050_rst), .rdata(f1050_rdata));
  assign f1050_clk = clk;
  assign f1050_rst = rst;
  // Bindings to f1050

  // f1052
  logic [0:0] f1052_wen;
  logic [31:0] f1052_wdata;
  logic [0:0] f1052_clk;
  logic [0:0] f1052_rst;
  logic [31:0] f1052_rdata;
  sr_buffer_32_1 f1052(.wen(f1052_wen), .wdata(f1052_wdata), .clk(f1052_clk), .rst(f1052_rst), .rdata(f1052_rdata));
  assign f1052_clk = clk;
  assign f1052_rst = rst;
  // Bindings to f1052

  // f1054
  logic [0:0] f1054_wen;
  logic [31:0] f1054_wdata;
  logic [0:0] f1054_clk;
  logic [0:0] f1054_rst;
  logic [31:0] f1054_rdata;
  sr_buffer_32_1 f1054(.wen(f1054_wen), .wdata(f1054_wdata), .clk(f1054_clk), .rst(f1054_rst), .rdata(f1054_rdata));
  assign f1054_clk = clk;
  assign f1054_rst = rst;
  // Bindings to f1054

  // f1056
  logic [0:0] f1056_wen;
  logic [31:0] f1056_wdata;
  logic [0:0] f1056_clk;
  logic [0:0] f1056_rst;
  logic [31:0] f1056_rdata;
  sr_buffer_32_1 f1056(.wen(f1056_wen), .wdata(f1056_wdata), .clk(f1056_clk), .rst(f1056_rst), .rdata(f1056_rdata));
  assign f1056_clk = clk;
  assign f1056_rst = rst;
  // Bindings to f1056

  // f1058
  logic [0:0] f1058_wen;
  logic [31:0] f1058_wdata;
  logic [0:0] f1058_clk;
  logic [0:0] f1058_rst;
  logic [31:0] f1058_rdata;
  sr_buffer_32_1 f1058(.wen(f1058_wen), .wdata(f1058_wdata), .clk(f1058_clk), .rst(f1058_rst), .rdata(f1058_rdata));
  assign f1058_clk = clk;
  assign f1058_rst = rst;
  // Bindings to f1058

  // f1060
  logic [0:0] f1060_wen;
  logic [31:0] f1060_wdata;
  logic [0:0] f1060_clk;
  logic [0:0] f1060_rst;
  logic [31:0] f1060_rdata;
  sr_buffer_32_1 f1060(.wen(f1060_wen), .wdata(f1060_wdata), .clk(f1060_clk), .rst(f1060_rst), .rdata(f1060_rdata));
  assign f1060_clk = clk;
  assign f1060_rst = rst;
  // Bindings to f1060

  // f1062
  logic [0:0] f1062_wen;
  logic [31:0] f1062_wdata;
  logic [0:0] f1062_clk;
  logic [0:0] f1062_rst;
  logic [31:0] f1062_rdata;
  sr_buffer_32_1 f1062(.wen(f1062_wen), .wdata(f1062_wdata), .clk(f1062_clk), .rst(f1062_rst), .rdata(f1062_rdata));
  assign f1062_clk = clk;
  assign f1062_rst = rst;
  // Bindings to f1062

  // f1064
  logic [0:0] f1064_wen;
  logic [31:0] f1064_wdata;
  logic [0:0] f1064_clk;
  logic [0:0] f1064_rst;
  logic [31:0] f1064_rdata;
  sr_buffer_32_1 f1064(.wen(f1064_wen), .wdata(f1064_wdata), .clk(f1064_clk), .rst(f1064_rst), .rdata(f1064_rdata));
  assign f1064_clk = clk;
  assign f1064_rst = rst;
  // Bindings to f1064

  // f1066
  logic [0:0] f1066_wen;
  logic [31:0] f1066_wdata;
  logic [0:0] f1066_clk;
  logic [0:0] f1066_rst;
  logic [31:0] f1066_rdata;
  sr_buffer_32_1 f1066(.wen(f1066_wen), .wdata(f1066_wdata), .clk(f1066_clk), .rst(f1066_rst), .rdata(f1066_rdata));
  assign f1066_clk = clk;
  assign f1066_rst = rst;
  // Bindings to f1066

  // f1068
  logic [0:0] f1068_wen;
  logic [31:0] f1068_wdata;
  logic [0:0] f1068_clk;
  logic [0:0] f1068_rst;
  logic [31:0] f1068_rdata;
  sr_buffer_32_1 f1068(.wen(f1068_wen), .wdata(f1068_wdata), .clk(f1068_clk), .rst(f1068_rst), .rdata(f1068_rdata));
  assign f1068_clk = clk;
  assign f1068_rst = rst;
  // Bindings to f1068

  // f1070
  logic [0:0] f1070_wen;
  logic [31:0] f1070_wdata;
  logic [0:0] f1070_clk;
  logic [0:0] f1070_rst;
  logic [31:0] f1070_rdata;
  sr_buffer_32_1 f1070(.wen(f1070_wen), .wdata(f1070_wdata), .clk(f1070_clk), .rst(f1070_rst), .rdata(f1070_rdata));
  assign f1070_clk = clk;
  assign f1070_rst = rst;
  // Bindings to f1070

  // f1072
  logic [0:0] f1072_wen;
  logic [31:0] f1072_wdata;
  logic [0:0] f1072_clk;
  logic [0:0] f1072_rst;
  logic [31:0] f1072_rdata;
  sr_buffer_32_1 f1072(.wen(f1072_wen), .wdata(f1072_wdata), .clk(f1072_clk), .rst(f1072_rst), .rdata(f1072_rdata));
  assign f1072_clk = clk;
  assign f1072_rst = rst;
  // Bindings to f1072

  // f1074
  logic [0:0] f1074_wen;
  logic [31:0] f1074_wdata;
  logic [0:0] f1074_clk;
  logic [0:0] f1074_rst;
  logic [31:0] f1074_rdata;
  sr_buffer_32_1 f1074(.wen(f1074_wen), .wdata(f1074_wdata), .clk(f1074_clk), .rst(f1074_rst), .rdata(f1074_rdata));
  assign f1074_clk = clk;
  assign f1074_rst = rst;
  // Bindings to f1074

  // f1076
  logic [0:0] f1076_wen;
  logic [31:0] f1076_wdata;
  logic [0:0] f1076_clk;
  logic [0:0] f1076_rst;
  logic [31:0] f1076_rdata;
  sr_buffer_32_1 f1076(.wen(f1076_wen), .wdata(f1076_wdata), .clk(f1076_clk), .rst(f1076_rst), .rdata(f1076_rdata));
  assign f1076_clk = clk;
  assign f1076_rst = rst;
  // Bindings to f1076

  // f1078
  logic [0:0] f1078_wen;
  logic [31:0] f1078_wdata;
  logic [0:0] f1078_clk;
  logic [0:0] f1078_rst;
  logic [31:0] f1078_rdata;
  sr_buffer_32_1 f1078(.wen(f1078_wen), .wdata(f1078_wdata), .clk(f1078_clk), .rst(f1078_rst), .rdata(f1078_rdata));
  assign f1078_clk = clk;
  assign f1078_rst = rst;
  // Bindings to f1078

  // f1080
  logic [0:0] f1080_wen;
  logic [31:0] f1080_wdata;
  logic [0:0] f1080_clk;
  logic [0:0] f1080_rst;
  logic [31:0] f1080_rdata;
  sr_buffer_32_1 f1080(.wen(f1080_wen), .wdata(f1080_wdata), .clk(f1080_clk), .rst(f1080_rst), .rdata(f1080_rdata));
  assign f1080_clk = clk;
  assign f1080_rst = rst;
  // Bindings to f1080

  // f1082
  logic [0:0] f1082_wen;
  logic [31:0] f1082_wdata;
  logic [0:0] f1082_clk;
  logic [0:0] f1082_rst;
  logic [31:0] f1082_rdata;
  sr_buffer_32_1 f1082(.wen(f1082_wen), .wdata(f1082_wdata), .clk(f1082_clk), .rst(f1082_rst), .rdata(f1082_rdata));
  assign f1082_clk = clk;
  assign f1082_rst = rst;
  // Bindings to f1082

  // f1084
  logic [0:0] f1084_wen;
  logic [31:0] f1084_wdata;
  logic [0:0] f1084_clk;
  logic [0:0] f1084_rst;
  logic [31:0] f1084_rdata;
  sr_buffer_32_1 f1084(.wen(f1084_wen), .wdata(f1084_wdata), .clk(f1084_clk), .rst(f1084_rst), .rdata(f1084_rdata));
  assign f1084_clk = clk;
  assign f1084_rst = rst;
  // Bindings to f1084

  // f1086
  logic [0:0] f1086_wen;
  logic [31:0] f1086_wdata;
  logic [0:0] f1086_clk;
  logic [0:0] f1086_rst;
  logic [31:0] f1086_rdata;
  sr_buffer_32_1 f1086(.wen(f1086_wen), .wdata(f1086_wdata), .clk(f1086_clk), .rst(f1086_rst), .rdata(f1086_rdata));
  assign f1086_clk = clk;
  assign f1086_rst = rst;
  // Bindings to f1086

  // f1088
  logic [0:0] f1088_wen;
  logic [31:0] f1088_wdata;
  logic [0:0] f1088_clk;
  logic [0:0] f1088_rst;
  logic [31:0] f1088_rdata;
  sr_buffer_32_1 f1088(.wen(f1088_wen), .wdata(f1088_wdata), .clk(f1088_clk), .rst(f1088_rst), .rdata(f1088_rdata));
  assign f1088_clk = clk;
  assign f1088_rst = rst;
  // Bindings to f1088

  // f1090
  logic [0:0] f1090_wen;
  logic [31:0] f1090_wdata;
  logic [0:0] f1090_clk;
  logic [0:0] f1090_rst;
  logic [31:0] f1090_rdata;
  sr_buffer_32_1 f1090(.wen(f1090_wen), .wdata(f1090_wdata), .clk(f1090_clk), .rst(f1090_rst), .rdata(f1090_rdata));
  assign f1090_clk = clk;
  assign f1090_rst = rst;
  // Bindings to f1090

  // f1092
  logic [0:0] f1092_wen;
  logic [31:0] f1092_wdata;
  logic [0:0] f1092_clk;
  logic [0:0] f1092_rst;
  logic [31:0] f1092_rdata;
  sr_buffer_32_1 f1092(.wen(f1092_wen), .wdata(f1092_wdata), .clk(f1092_clk), .rst(f1092_rst), .rdata(f1092_rdata));
  assign f1092_clk = clk;
  assign f1092_rst = rst;
  // Bindings to f1092

  // f1094
  logic [0:0] f1094_wen;
  logic [31:0] f1094_wdata;
  logic [0:0] f1094_clk;
  logic [0:0] f1094_rst;
  logic [31:0] f1094_rdata;
  sr_buffer_32_1 f1094(.wen(f1094_wen), .wdata(f1094_wdata), .clk(f1094_clk), .rst(f1094_rst), .rdata(f1094_rdata));
  assign f1094_clk = clk;
  assign f1094_rst = rst;
  // Bindings to f1094

  // f1096
  logic [0:0] f1096_wen;
  logic [31:0] f1096_wdata;
  logic [0:0] f1096_clk;
  logic [0:0] f1096_rst;
  logic [31:0] f1096_rdata;
  sr_buffer_32_1 f1096(.wen(f1096_wen), .wdata(f1096_wdata), .clk(f1096_clk), .rst(f1096_rst), .rdata(f1096_rdata));
  assign f1096_clk = clk;
  assign f1096_rst = rst;
  // Bindings to f1096

  // f1098
  logic [0:0] f1098_wen;
  logic [31:0] f1098_wdata;
  logic [0:0] f1098_clk;
  logic [0:0] f1098_rst;
  logic [31:0] f1098_rdata;
  sr_buffer_32_1 f1098(.wen(f1098_wen), .wdata(f1098_wdata), .clk(f1098_clk), .rst(f1098_rst), .rdata(f1098_rdata));
  assign f1098_clk = clk;
  assign f1098_rst = rst;
  // Bindings to f1098

  // f1100
  logic [0:0] f1100_wen;
  logic [31:0] f1100_wdata;
  logic [0:0] f1100_clk;
  logic [0:0] f1100_rst;
  logic [31:0] f1100_rdata;
  sr_buffer_32_1 f1100(.wen(f1100_wen), .wdata(f1100_wdata), .clk(f1100_clk), .rst(f1100_rst), .rdata(f1100_rdata));
  assign f1100_clk = clk;
  assign f1100_rst = rst;
  // Bindings to f1100

  // f1102
  logic [0:0] f1102_wen;
  logic [31:0] f1102_wdata;
  logic [0:0] f1102_clk;
  logic [0:0] f1102_rst;
  logic [31:0] f1102_rdata;
  sr_buffer_32_1 f1102(.wen(f1102_wen), .wdata(f1102_wdata), .clk(f1102_clk), .rst(f1102_rst), .rdata(f1102_rdata));
  assign f1102_clk = clk;
  assign f1102_rst = rst;
  // Bindings to f1102

  // f1104
  logic [0:0] f1104_wen;
  logic [31:0] f1104_wdata;
  logic [0:0] f1104_clk;
  logic [0:0] f1104_rst;
  logic [31:0] f1104_rdata;
  sr_buffer_32_1 f1104(.wen(f1104_wen), .wdata(f1104_wdata), .clk(f1104_clk), .rst(f1104_rst), .rdata(f1104_rdata));
  assign f1104_clk = clk;
  assign f1104_rst = rst;
  // Bindings to f1104

  // f1106
  logic [0:0] f1106_wen;
  logic [31:0] f1106_wdata;
  logic [0:0] f1106_clk;
  logic [0:0] f1106_rst;
  logic [31:0] f1106_rdata;
  sr_buffer_32_1 f1106(.wen(f1106_wen), .wdata(f1106_wdata), .clk(f1106_clk), .rst(f1106_rst), .rdata(f1106_rdata));
  assign f1106_clk = clk;
  assign f1106_rst = rst;
  // Bindings to f1106

  // f1108
  logic [0:0] f1108_wen;
  logic [31:0] f1108_wdata;
  logic [0:0] f1108_clk;
  logic [0:0] f1108_rst;
  logic [31:0] f1108_rdata;
  sr_buffer_32_1 f1108(.wen(f1108_wen), .wdata(f1108_wdata), .clk(f1108_clk), .rst(f1108_rst), .rdata(f1108_rdata));
  assign f1108_clk = clk;
  assign f1108_rst = rst;
  // Bindings to f1108

  // f1110
  logic [0:0] f1110_wen;
  logic [31:0] f1110_wdata;
  logic [0:0] f1110_clk;
  logic [0:0] f1110_rst;
  logic [31:0] f1110_rdata;
  sr_buffer_32_1 f1110(.wen(f1110_wen), .wdata(f1110_wdata), .clk(f1110_clk), .rst(f1110_rst), .rdata(f1110_rdata));
  assign f1110_clk = clk;
  assign f1110_rst = rst;
  // Bindings to f1110

  // f1112
  logic [0:0] f1112_wen;
  logic [31:0] f1112_wdata;
  logic [0:0] f1112_clk;
  logic [0:0] f1112_rst;
  logic [31:0] f1112_rdata;
  sr_buffer_32_1 f1112(.wen(f1112_wen), .wdata(f1112_wdata), .clk(f1112_clk), .rst(f1112_rst), .rdata(f1112_rdata));
  assign f1112_clk = clk;
  assign f1112_rst = rst;
  // Bindings to f1112

  // f1114
  logic [0:0] f1114_wen;
  logic [31:0] f1114_wdata;
  logic [0:0] f1114_clk;
  logic [0:0] f1114_rst;
  logic [31:0] f1114_rdata;
  sr_buffer_32_1 f1114(.wen(f1114_wen), .wdata(f1114_wdata), .clk(f1114_clk), .rst(f1114_rst), .rdata(f1114_rdata));
  assign f1114_clk = clk;
  assign f1114_rst = rst;
  // Bindings to f1114

  // f1116
  logic [0:0] f1116_wen;
  logic [31:0] f1116_wdata;
  logic [0:0] f1116_clk;
  logic [0:0] f1116_rst;
  logic [31:0] f1116_rdata;
  sr_buffer_32_1 f1116(.wen(f1116_wen), .wdata(f1116_wdata), .clk(f1116_clk), .rst(f1116_rst), .rdata(f1116_rdata));
  assign f1116_clk = clk;
  assign f1116_rst = rst;
  // Bindings to f1116

  // f1118
  logic [0:0] f1118_wen;
  logic [31:0] f1118_wdata;
  logic [0:0] f1118_clk;
  logic [0:0] f1118_rst;
  logic [31:0] f1118_rdata;
  sr_buffer_32_1 f1118(.wen(f1118_wen), .wdata(f1118_wdata), .clk(f1118_clk), .rst(f1118_rst), .rdata(f1118_rdata));
  assign f1118_clk = clk;
  assign f1118_rst = rst;
  // Bindings to f1118

  // f1120
  logic [0:0] f1120_wen;
  logic [31:0] f1120_wdata;
  logic [0:0] f1120_clk;
  logic [0:0] f1120_rst;
  logic [31:0] f1120_rdata;
  sr_buffer_32_1 f1120(.wen(f1120_wen), .wdata(f1120_wdata), .clk(f1120_clk), .rst(f1120_rst), .rdata(f1120_rdata));
  assign f1120_clk = clk;
  assign f1120_rst = rst;
  // Bindings to f1120

  // f1122
  logic [0:0] f1122_wen;
  logic [31:0] f1122_wdata;
  logic [0:0] f1122_clk;
  logic [0:0] f1122_rst;
  logic [31:0] f1122_rdata;
  sr_buffer_32_1 f1122(.wen(f1122_wen), .wdata(f1122_wdata), .clk(f1122_clk), .rst(f1122_rst), .rdata(f1122_rdata));
  assign f1122_clk = clk;
  assign f1122_rst = rst;
  // Bindings to f1122

  // f1124
  logic [0:0] f1124_wen;
  logic [31:0] f1124_wdata;
  logic [0:0] f1124_clk;
  logic [0:0] f1124_rst;
  logic [31:0] f1124_rdata;
  sr_buffer_32_1 f1124(.wen(f1124_wen), .wdata(f1124_wdata), .clk(f1124_clk), .rst(f1124_rst), .rdata(f1124_rdata));
  assign f1124_clk = clk;
  assign f1124_rst = rst;
  // Bindings to f1124

  // f1126
  logic [0:0] f1126_wen;
  logic [31:0] f1126_wdata;
  logic [0:0] f1126_clk;
  logic [0:0] f1126_rst;
  logic [31:0] f1126_rdata;
  sr_buffer_32_1 f1126(.wen(f1126_wen), .wdata(f1126_wdata), .clk(f1126_clk), .rst(f1126_rst), .rdata(f1126_rdata));
  assign f1126_clk = clk;
  assign f1126_rst = rst;
  // Bindings to f1126

  // f1128
  logic [0:0] f1128_wen;
  logic [31:0] f1128_wdata;
  logic [0:0] f1128_clk;
  logic [0:0] f1128_rst;
  logic [31:0] f1128_rdata;
  sr_buffer_32_1 f1128(.wen(f1128_wen), .wdata(f1128_wdata), .clk(f1128_clk), .rst(f1128_rst), .rdata(f1128_rdata));
  assign f1128_clk = clk;
  assign f1128_rst = rst;
  // Bindings to f1128

  // f1130
  logic [0:0] f1130_wen;
  logic [31:0] f1130_wdata;
  logic [0:0] f1130_clk;
  logic [0:0] f1130_rst;
  logic [31:0] f1130_rdata;
  sr_buffer_32_1 f1130(.wen(f1130_wen), .wdata(f1130_wdata), .clk(f1130_clk), .rst(f1130_rst), .rdata(f1130_rdata));
  assign f1130_clk = clk;
  assign f1130_rst = rst;
  // Bindings to f1130

  // f1132
  logic [0:0] f1132_wen;
  logic [31:0] f1132_wdata;
  logic [0:0] f1132_clk;
  logic [0:0] f1132_rst;
  logic [31:0] f1132_rdata;
  sr_buffer_32_1 f1132(.wen(f1132_wen), .wdata(f1132_wdata), .clk(f1132_clk), .rst(f1132_rst), .rdata(f1132_rdata));
  assign f1132_clk = clk;
  assign f1132_rst = rst;
  // Bindings to f1132

  // f1134
  logic [0:0] f1134_wen;
  logic [31:0] f1134_wdata;
  logic [0:0] f1134_clk;
  logic [0:0] f1134_rst;
  logic [31:0] f1134_rdata;
  sr_buffer_32_1 f1134(.wen(f1134_wen), .wdata(f1134_wdata), .clk(f1134_clk), .rst(f1134_rst), .rdata(f1134_rdata));
  assign f1134_clk = clk;
  assign f1134_rst = rst;
  // Bindings to f1134

  // f1136
  logic [0:0] f1136_wen;
  logic [31:0] f1136_wdata;
  logic [0:0] f1136_clk;
  logic [0:0] f1136_rst;
  logic [31:0] f1136_rdata;
  sr_buffer_32_1 f1136(.wen(f1136_wen), .wdata(f1136_wdata), .clk(f1136_clk), .rst(f1136_rst), .rdata(f1136_rdata));
  assign f1136_clk = clk;
  assign f1136_rst = rst;
  // Bindings to f1136

  // f1138
  logic [0:0] f1138_wen;
  logic [31:0] f1138_wdata;
  logic [0:0] f1138_clk;
  logic [0:0] f1138_rst;
  logic [31:0] f1138_rdata;
  sr_buffer_32_1 f1138(.wen(f1138_wen), .wdata(f1138_wdata), .clk(f1138_clk), .rst(f1138_rst), .rdata(f1138_rdata));
  assign f1138_clk = clk;
  assign f1138_rst = rst;
  // Bindings to f1138

  // f1140
  logic [0:0] f1140_wen;
  logic [31:0] f1140_wdata;
  logic [0:0] f1140_clk;
  logic [0:0] f1140_rst;
  logic [31:0] f1140_rdata;
  sr_buffer_32_1 f1140(.wen(f1140_wen), .wdata(f1140_wdata), .clk(f1140_clk), .rst(f1140_rst), .rdata(f1140_rdata));
  assign f1140_clk = clk;
  assign f1140_rst = rst;
  // Bindings to f1140

  // f1142
  logic [0:0] f1142_wen;
  logic [31:0] f1142_wdata;
  logic [0:0] f1142_clk;
  logic [0:0] f1142_rst;
  logic [31:0] f1142_rdata;
  sr_buffer_32_1 f1142(.wen(f1142_wen), .wdata(f1142_wdata), .clk(f1142_clk), .rst(f1142_rst), .rdata(f1142_rdata));
  assign f1142_clk = clk;
  assign f1142_rst = rst;
  // Bindings to f1142

  // f1144
  logic [0:0] f1144_wen;
  logic [31:0] f1144_wdata;
  logic [0:0] f1144_clk;
  logic [0:0] f1144_rst;
  logic [31:0] f1144_rdata;
  sr_buffer_32_1 f1144(.wen(f1144_wen), .wdata(f1144_wdata), .clk(f1144_clk), .rst(f1144_rst), .rdata(f1144_rdata));
  assign f1144_clk = clk;
  assign f1144_rst = rst;
  // Bindings to f1144

  // f1146
  logic [0:0] f1146_wen;
  logic [31:0] f1146_wdata;
  logic [0:0] f1146_clk;
  logic [0:0] f1146_rst;
  logic [31:0] f1146_rdata;
  sr_buffer_32_1 f1146(.wen(f1146_wen), .wdata(f1146_wdata), .clk(f1146_clk), .rst(f1146_rst), .rdata(f1146_rdata));
  assign f1146_clk = clk;
  assign f1146_rst = rst;
  // Bindings to f1146

  // f1148
  logic [0:0] f1148_wen;
  logic [31:0] f1148_wdata;
  logic [0:0] f1148_clk;
  logic [0:0] f1148_rst;
  logic [31:0] f1148_rdata;
  sr_buffer_32_1 f1148(.wen(f1148_wen), .wdata(f1148_wdata), .clk(f1148_clk), .rst(f1148_rst), .rdata(f1148_rdata));
  assign f1148_clk = clk;
  assign f1148_rst = rst;
  // Bindings to f1148

  // f1150
  logic [0:0] f1150_wen;
  logic [31:0] f1150_wdata;
  logic [0:0] f1150_clk;
  logic [0:0] f1150_rst;
  logic [31:0] f1150_rdata;
  sr_buffer_32_1 f1150(.wen(f1150_wen), .wdata(f1150_wdata), .clk(f1150_clk), .rst(f1150_rst), .rdata(f1150_rdata));
  assign f1150_clk = clk;
  assign f1150_rst = rst;
  // Bindings to f1150

  // f1152
  logic [0:0] f1152_wen;
  logic [31:0] f1152_wdata;
  logic [0:0] f1152_clk;
  logic [0:0] f1152_rst;
  logic [31:0] f1152_rdata;
  sr_buffer_32_1 f1152(.wen(f1152_wen), .wdata(f1152_wdata), .clk(f1152_clk), .rst(f1152_rst), .rdata(f1152_rdata));
  assign f1152_clk = clk;
  assign f1152_rst = rst;
  // Bindings to f1152

  // f1154
  logic [0:0] f1154_wen;
  logic [31:0] f1154_wdata;
  logic [0:0] f1154_clk;
  logic [0:0] f1154_rst;
  logic [31:0] f1154_rdata;
  sr_buffer_32_1 f1154(.wen(f1154_wen), .wdata(f1154_wdata), .clk(f1154_clk), .rst(f1154_rst), .rdata(f1154_rdata));
  assign f1154_clk = clk;
  assign f1154_rst = rst;
  // Bindings to f1154

  // f1156
  logic [0:0] f1156_wen;
  logic [31:0] f1156_wdata;
  logic [0:0] f1156_clk;
  logic [0:0] f1156_rst;
  logic [31:0] f1156_rdata;
  sr_buffer_32_1 f1156(.wen(f1156_wen), .wdata(f1156_wdata), .clk(f1156_clk), .rst(f1156_rst), .rdata(f1156_rdata));
  assign f1156_clk = clk;
  assign f1156_rst = rst;
  // Bindings to f1156

  // f1158
  logic [0:0] f1158_wen;
  logic [31:0] f1158_wdata;
  logic [0:0] f1158_clk;
  logic [0:0] f1158_rst;
  logic [31:0] f1158_rdata;
  sr_buffer_32_1 f1158(.wen(f1158_wen), .wdata(f1158_wdata), .clk(f1158_clk), .rst(f1158_rst), .rdata(f1158_rdata));
  assign f1158_clk = clk;
  assign f1158_rst = rst;
  // Bindings to f1158

  // f1160
  logic [0:0] f1160_wen;
  logic [31:0] f1160_wdata;
  logic [0:0] f1160_clk;
  logic [0:0] f1160_rst;
  logic [31:0] f1160_rdata;
  sr_buffer_32_1 f1160(.wen(f1160_wen), .wdata(f1160_wdata), .clk(f1160_clk), .rst(f1160_rst), .rdata(f1160_rdata));
  assign f1160_clk = clk;
  assign f1160_rst = rst;
  // Bindings to f1160

  // f1162
  logic [0:0] f1162_wen;
  logic [31:0] f1162_wdata;
  logic [0:0] f1162_clk;
  logic [0:0] f1162_rst;
  logic [31:0] f1162_rdata;
  sr_buffer_32_1 f1162(.wen(f1162_wen), .wdata(f1162_wdata), .clk(f1162_clk), .rst(f1162_rst), .rdata(f1162_rdata));
  assign f1162_clk = clk;
  assign f1162_rst = rst;
  // Bindings to f1162

  // f1164
  logic [0:0] f1164_wen;
  logic [31:0] f1164_wdata;
  logic [0:0] f1164_clk;
  logic [0:0] f1164_rst;
  logic [31:0] f1164_rdata;
  sr_buffer_32_1 f1164(.wen(f1164_wen), .wdata(f1164_wdata), .clk(f1164_clk), .rst(f1164_rst), .rdata(f1164_rdata));
  assign f1164_clk = clk;
  assign f1164_rst = rst;
  // Bindings to f1164

  // f1166
  logic [0:0] f1166_wen;
  logic [31:0] f1166_wdata;
  logic [0:0] f1166_clk;
  logic [0:0] f1166_rst;
  logic [31:0] f1166_rdata;
  sr_buffer_32_1 f1166(.wen(f1166_wen), .wdata(f1166_wdata), .clk(f1166_clk), .rst(f1166_rst), .rdata(f1166_rdata));
  assign f1166_clk = clk;
  assign f1166_rst = rst;
  // Bindings to f1166

  // f1168
  logic [0:0] f1168_wen;
  logic [31:0] f1168_wdata;
  logic [0:0] f1168_clk;
  logic [0:0] f1168_rst;
  logic [31:0] f1168_rdata;
  sr_buffer_32_1 f1168(.wen(f1168_wen), .wdata(f1168_wdata), .clk(f1168_clk), .rst(f1168_rst), .rdata(f1168_rdata));
  assign f1168_clk = clk;
  assign f1168_rst = rst;
  // Bindings to f1168

  // f1170
  logic [0:0] f1170_wen;
  logic [31:0] f1170_wdata;
  logic [0:0] f1170_clk;
  logic [0:0] f1170_rst;
  logic [31:0] f1170_rdata;
  sr_buffer_32_1 f1170(.wen(f1170_wen), .wdata(f1170_wdata), .clk(f1170_clk), .rst(f1170_rst), .rdata(f1170_rdata));
  assign f1170_clk = clk;
  assign f1170_rst = rst;
  // Bindings to f1170

  // f1172
  logic [0:0] f1172_wen;
  logic [31:0] f1172_wdata;
  logic [0:0] f1172_clk;
  logic [0:0] f1172_rst;
  logic [31:0] f1172_rdata;
  sr_buffer_32_1 f1172(.wen(f1172_wen), .wdata(f1172_wdata), .clk(f1172_clk), .rst(f1172_rst), .rdata(f1172_rdata));
  assign f1172_clk = clk;
  assign f1172_rst = rst;
  // Bindings to f1172

  // f1174
  logic [0:0] f1174_wen;
  logic [31:0] f1174_wdata;
  logic [0:0] f1174_clk;
  logic [0:0] f1174_rst;
  logic [31:0] f1174_rdata;
  sr_buffer_32_1 f1174(.wen(f1174_wen), .wdata(f1174_wdata), .clk(f1174_clk), .rst(f1174_rst), .rdata(f1174_rdata));
  assign f1174_clk = clk;
  assign f1174_rst = rst;
  // Bindings to f1174

  // f1176
  logic [0:0] f1176_wen;
  logic [31:0] f1176_wdata;
  logic [0:0] f1176_clk;
  logic [0:0] f1176_rst;
  logic [31:0] f1176_rdata;
  sr_buffer_32_1 f1176(.wen(f1176_wen), .wdata(f1176_wdata), .clk(f1176_clk), .rst(f1176_rst), .rdata(f1176_rdata));
  assign f1176_clk = clk;
  assign f1176_rst = rst;
  // Bindings to f1176

  // f1178
  logic [0:0] f1178_wen;
  logic [31:0] f1178_wdata;
  logic [0:0] f1178_clk;
  logic [0:0] f1178_rst;
  logic [31:0] f1178_rdata;
  sr_buffer_32_1 f1178(.wen(f1178_wen), .wdata(f1178_wdata), .clk(f1178_clk), .rst(f1178_rst), .rdata(f1178_rdata));
  assign f1178_clk = clk;
  assign f1178_rst = rst;
  // Bindings to f1178

  // f1180
  logic [0:0] f1180_wen;
  logic [31:0] f1180_wdata;
  logic [0:0] f1180_clk;
  logic [0:0] f1180_rst;
  logic [31:0] f1180_rdata;
  sr_buffer_32_1 f1180(.wen(f1180_wen), .wdata(f1180_wdata), .clk(f1180_clk), .rst(f1180_rst), .rdata(f1180_rdata));
  assign f1180_clk = clk;
  assign f1180_rst = rst;
  // Bindings to f1180

  // f1182
  logic [0:0] f1182_wen;
  logic [31:0] f1182_wdata;
  logic [0:0] f1182_clk;
  logic [0:0] f1182_rst;
  logic [31:0] f1182_rdata;
  sr_buffer_32_1 f1182(.wen(f1182_wen), .wdata(f1182_wdata), .clk(f1182_clk), .rst(f1182_rst), .rdata(f1182_rdata));
  assign f1182_clk = clk;
  assign f1182_rst = rst;
  // Bindings to f1182

  // f1184
  logic [0:0] f1184_wen;
  logic [31:0] f1184_wdata;
  logic [0:0] f1184_clk;
  logic [0:0] f1184_rst;
  logic [31:0] f1184_rdata;
  sr_buffer_32_1 f1184(.wen(f1184_wen), .wdata(f1184_wdata), .clk(f1184_clk), .rst(f1184_rst), .rdata(f1184_rdata));
  assign f1184_clk = clk;
  assign f1184_rst = rst;
  // Bindings to f1184

  // f1186
  logic [0:0] f1186_wen;
  logic [31:0] f1186_wdata;
  logic [0:0] f1186_clk;
  logic [0:0] f1186_rst;
  logic [31:0] f1186_rdata;
  sr_buffer_32_1 f1186(.wen(f1186_wen), .wdata(f1186_wdata), .clk(f1186_clk), .rst(f1186_rst), .rdata(f1186_rdata));
  assign f1186_clk = clk;
  assign f1186_rst = rst;
  // Bindings to f1186

  // f1188
  logic [0:0] f1188_wen;
  logic [31:0] f1188_wdata;
  logic [0:0] f1188_clk;
  logic [0:0] f1188_rst;
  logic [31:0] f1188_rdata;
  sr_buffer_32_1 f1188(.wen(f1188_wen), .wdata(f1188_wdata), .clk(f1188_clk), .rst(f1188_rst), .rdata(f1188_rdata));
  assign f1188_clk = clk;
  assign f1188_rst = rst;
  // Bindings to f1188

  // f1190
  logic [0:0] f1190_wen;
  logic [31:0] f1190_wdata;
  logic [0:0] f1190_clk;
  logic [0:0] f1190_rst;
  logic [31:0] f1190_rdata;
  sr_buffer_32_1 f1190(.wen(f1190_wen), .wdata(f1190_wdata), .clk(f1190_clk), .rst(f1190_rst), .rdata(f1190_rdata));
  assign f1190_clk = clk;
  assign f1190_rst = rst;
  // Bindings to f1190

  // f1192
  logic [0:0] f1192_wen;
  logic [31:0] f1192_wdata;
  logic [0:0] f1192_clk;
  logic [0:0] f1192_rst;
  logic [31:0] f1192_rdata;
  sr_buffer_32_1 f1192(.wen(f1192_wen), .wdata(f1192_wdata), .clk(f1192_clk), .rst(f1192_rst), .rdata(f1192_rdata));
  assign f1192_clk = clk;
  assign f1192_rst = rst;
  // Bindings to f1192

  // f1194
  logic [0:0] f1194_wen;
  logic [31:0] f1194_wdata;
  logic [0:0] f1194_clk;
  logic [0:0] f1194_rst;
  logic [31:0] f1194_rdata;
  sr_buffer_32_1 f1194(.wen(f1194_wen), .wdata(f1194_wdata), .clk(f1194_clk), .rst(f1194_rst), .rdata(f1194_rdata));
  assign f1194_clk = clk;
  assign f1194_rst = rst;
  // Bindings to f1194

  // f1196
  logic [0:0] f1196_wen;
  logic [31:0] f1196_wdata;
  logic [0:0] f1196_clk;
  logic [0:0] f1196_rst;
  logic [31:0] f1196_rdata;
  sr_buffer_32_1 f1196(.wen(f1196_wen), .wdata(f1196_wdata), .clk(f1196_clk), .rst(f1196_rst), .rdata(f1196_rdata));
  assign f1196_clk = clk;
  assign f1196_rst = rst;
  // Bindings to f1196

  // f1198
  logic [0:0] f1198_wen;
  logic [31:0] f1198_wdata;
  logic [0:0] f1198_clk;
  logic [0:0] f1198_rst;
  logic [31:0] f1198_rdata;
  sr_buffer_32_1 f1198(.wen(f1198_wen), .wdata(f1198_wdata), .clk(f1198_clk), .rst(f1198_rst), .rdata(f1198_rdata));
  assign f1198_clk = clk;
  assign f1198_rst = rst;
  // Bindings to f1198

  // f1200
  logic [0:0] f1200_wen;
  logic [31:0] f1200_wdata;
  logic [0:0] f1200_clk;
  logic [0:0] f1200_rst;
  logic [31:0] f1200_rdata;
  sr_buffer_32_1 f1200(.wen(f1200_wen), .wdata(f1200_wdata), .clk(f1200_clk), .rst(f1200_rst), .rdata(f1200_rdata));
  assign f1200_clk = clk;
  assign f1200_rst = rst;
  // Bindings to f1200

  // f1202
  logic [0:0] f1202_wen;
  logic [31:0] f1202_wdata;
  logic [0:0] f1202_clk;
  logic [0:0] f1202_rst;
  logic [31:0] f1202_rdata;
  sr_buffer_32_1 f1202(.wen(f1202_wen), .wdata(f1202_wdata), .clk(f1202_clk), .rst(f1202_rst), .rdata(f1202_rdata));
  assign f1202_clk = clk;
  assign f1202_rst = rst;
  // Bindings to f1202

  // f1204
  logic [0:0] f1204_wen;
  logic [31:0] f1204_wdata;
  logic [0:0] f1204_clk;
  logic [0:0] f1204_rst;
  logic [31:0] f1204_rdata;
  sr_buffer_32_1 f1204(.wen(f1204_wen), .wdata(f1204_wdata), .clk(f1204_clk), .rst(f1204_rst), .rdata(f1204_rdata));
  assign f1204_clk = clk;
  assign f1204_rst = rst;
  // Bindings to f1204

  // f1206
  logic [0:0] f1206_wen;
  logic [31:0] f1206_wdata;
  logic [0:0] f1206_clk;
  logic [0:0] f1206_rst;
  logic [31:0] f1206_rdata;
  sr_buffer_32_1 f1206(.wen(f1206_wen), .wdata(f1206_wdata), .clk(f1206_clk), .rst(f1206_rst), .rdata(f1206_rdata));
  assign f1206_clk = clk;
  assign f1206_rst = rst;
  // Bindings to f1206

  // f1208
  logic [0:0] f1208_wen;
  logic [31:0] f1208_wdata;
  logic [0:0] f1208_clk;
  logic [0:0] f1208_rst;
  logic [31:0] f1208_rdata;
  sr_buffer_32_1 f1208(.wen(f1208_wen), .wdata(f1208_wdata), .clk(f1208_clk), .rst(f1208_rst), .rdata(f1208_rdata));
  assign f1208_clk = clk;
  assign f1208_rst = rst;
  // Bindings to f1208

  // f1210
  logic [0:0] f1210_wen;
  logic [31:0] f1210_wdata;
  logic [0:0] f1210_clk;
  logic [0:0] f1210_rst;
  logic [31:0] f1210_rdata;
  sr_buffer_32_1 f1210(.wen(f1210_wen), .wdata(f1210_wdata), .clk(f1210_clk), .rst(f1210_rst), .rdata(f1210_rdata));
  assign f1210_clk = clk;
  assign f1210_rst = rst;
  // Bindings to f1210

  // f1212
  logic [0:0] f1212_wen;
  logic [31:0] f1212_wdata;
  logic [0:0] f1212_clk;
  logic [0:0] f1212_rst;
  logic [31:0] f1212_rdata;
  sr_buffer_32_1 f1212(.wen(f1212_wen), .wdata(f1212_wdata), .clk(f1212_clk), .rst(f1212_rst), .rdata(f1212_rdata));
  assign f1212_clk = clk;
  assign f1212_rst = rst;
  // Bindings to f1212

  // f1214
  logic [0:0] f1214_wen;
  logic [31:0] f1214_wdata;
  logic [0:0] f1214_clk;
  logic [0:0] f1214_rst;
  logic [31:0] f1214_rdata;
  sr_buffer_32_1 f1214(.wen(f1214_wen), .wdata(f1214_wdata), .clk(f1214_clk), .rst(f1214_rst), .rdata(f1214_rdata));
  assign f1214_clk = clk;
  assign f1214_rst = rst;
  // Bindings to f1214

  // f1216
  logic [0:0] f1216_wen;
  logic [31:0] f1216_wdata;
  logic [0:0] f1216_clk;
  logic [0:0] f1216_rst;
  logic [31:0] f1216_rdata;
  sr_buffer_32_1 f1216(.wen(f1216_wen), .wdata(f1216_wdata), .clk(f1216_clk), .rst(f1216_rst), .rdata(f1216_rdata));
  assign f1216_clk = clk;
  assign f1216_rst = rst;
  // Bindings to f1216

  // f1218
  logic [0:0] f1218_wen;
  logic [31:0] f1218_wdata;
  logic [0:0] f1218_clk;
  logic [0:0] f1218_rst;
  logic [31:0] f1218_rdata;
  sr_buffer_32_1 f1218(.wen(f1218_wen), .wdata(f1218_wdata), .clk(f1218_clk), .rst(f1218_rst), .rdata(f1218_rdata));
  assign f1218_clk = clk;
  assign f1218_rst = rst;
  // Bindings to f1218

  // f1220
  logic [0:0] f1220_wen;
  logic [31:0] f1220_wdata;
  logic [0:0] f1220_clk;
  logic [0:0] f1220_rst;
  logic [31:0] f1220_rdata;
  sr_buffer_32_1 f1220(.wen(f1220_wen), .wdata(f1220_wdata), .clk(f1220_clk), .rst(f1220_rst), .rdata(f1220_rdata));
  assign f1220_clk = clk;
  assign f1220_rst = rst;
  // Bindings to f1220

  // f1222
  logic [0:0] f1222_wen;
  logic [31:0] f1222_wdata;
  logic [0:0] f1222_clk;
  logic [0:0] f1222_rst;
  logic [31:0] f1222_rdata;
  sr_buffer_32_1 f1222(.wen(f1222_wen), .wdata(f1222_wdata), .clk(f1222_clk), .rst(f1222_rst), .rdata(f1222_rdata));
  assign f1222_clk = clk;
  assign f1222_rst = rst;
  // Bindings to f1222

  // f1224
  logic [0:0] f1224_wen;
  logic [31:0] f1224_wdata;
  logic [0:0] f1224_clk;
  logic [0:0] f1224_rst;
  logic [31:0] f1224_rdata;
  sr_buffer_32_1 f1224(.wen(f1224_wen), .wdata(f1224_wdata), .clk(f1224_clk), .rst(f1224_rst), .rdata(f1224_rdata));
  assign f1224_clk = clk;
  assign f1224_rst = rst;
  // Bindings to f1224

  // f1226
  logic [0:0] f1226_wen;
  logic [31:0] f1226_wdata;
  logic [0:0] f1226_clk;
  logic [0:0] f1226_rst;
  logic [31:0] f1226_rdata;
  sr_buffer_32_1 f1226(.wen(f1226_wen), .wdata(f1226_wdata), .clk(f1226_clk), .rst(f1226_rst), .rdata(f1226_rdata));
  assign f1226_clk = clk;
  assign f1226_rst = rst;
  // Bindings to f1226

  // f1228
  logic [0:0] f1228_wen;
  logic [31:0] f1228_wdata;
  logic [0:0] f1228_clk;
  logic [0:0] f1228_rst;
  logic [31:0] f1228_rdata;
  sr_buffer_32_1 f1228(.wen(f1228_wen), .wdata(f1228_wdata), .clk(f1228_clk), .rst(f1228_rst), .rdata(f1228_rdata));
  assign f1228_clk = clk;
  assign f1228_rst = rst;
  // Bindings to f1228

  // f1230
  logic [0:0] f1230_wen;
  logic [31:0] f1230_wdata;
  logic [0:0] f1230_clk;
  logic [0:0] f1230_rst;
  logic [31:0] f1230_rdata;
  sr_buffer_32_1 f1230(.wen(f1230_wen), .wdata(f1230_wdata), .clk(f1230_clk), .rst(f1230_rst), .rdata(f1230_rdata));
  assign f1230_clk = clk;
  assign f1230_rst = rst;
  // Bindings to f1230

  // f1232
  logic [0:0] f1232_wen;
  logic [31:0] f1232_wdata;
  logic [0:0] f1232_clk;
  logic [0:0] f1232_rst;
  logic [31:0] f1232_rdata;
  sr_buffer_32_1 f1232(.wen(f1232_wen), .wdata(f1232_wdata), .clk(f1232_clk), .rst(f1232_rst), .rdata(f1232_rdata));
  assign f1232_clk = clk;
  assign f1232_rst = rst;
  // Bindings to f1232

  // f1234
  logic [0:0] f1234_wen;
  logic [31:0] f1234_wdata;
  logic [0:0] f1234_clk;
  logic [0:0] f1234_rst;
  logic [31:0] f1234_rdata;
  sr_buffer_32_1 f1234(.wen(f1234_wen), .wdata(f1234_wdata), .clk(f1234_clk), .rst(f1234_rst), .rdata(f1234_rdata));
  assign f1234_clk = clk;
  assign f1234_rst = rst;
  // Bindings to f1234

  // f1236
  logic [0:0] f1236_wen;
  logic [31:0] f1236_wdata;
  logic [0:0] f1236_clk;
  logic [0:0] f1236_rst;
  logic [31:0] f1236_rdata;
  sr_buffer_32_1 f1236(.wen(f1236_wen), .wdata(f1236_wdata), .clk(f1236_clk), .rst(f1236_rst), .rdata(f1236_rdata));
  assign f1236_clk = clk;
  assign f1236_rst = rst;
  // Bindings to f1236

  // f1238
  logic [0:0] f1238_wen;
  logic [31:0] f1238_wdata;
  logic [0:0] f1238_clk;
  logic [0:0] f1238_rst;
  logic [31:0] f1238_rdata;
  sr_buffer_32_1 f1238(.wen(f1238_wen), .wdata(f1238_wdata), .clk(f1238_clk), .rst(f1238_rst), .rdata(f1238_rdata));
  assign f1238_clk = clk;
  assign f1238_rst = rst;
  // Bindings to f1238

  // f1240
  logic [0:0] f1240_wen;
  logic [31:0] f1240_wdata;
  logic [0:0] f1240_clk;
  logic [0:0] f1240_rst;
  logic [31:0] f1240_rdata;
  sr_buffer_32_1 f1240(.wen(f1240_wen), .wdata(f1240_wdata), .clk(f1240_clk), .rst(f1240_rst), .rdata(f1240_rdata));
  assign f1240_clk = clk;
  assign f1240_rst = rst;
  // Bindings to f1240

  // f1242
  logic [0:0] f1242_wen;
  logic [31:0] f1242_wdata;
  logic [0:0] f1242_clk;
  logic [0:0] f1242_rst;
  logic [31:0] f1242_rdata;
  sr_buffer_32_1 f1242(.wen(f1242_wen), .wdata(f1242_wdata), .clk(f1242_clk), .rst(f1242_rst), .rdata(f1242_rdata));
  assign f1242_clk = clk;
  assign f1242_rst = rst;
  // Bindings to f1242

  // f1244
  logic [0:0] f1244_wen;
  logic [31:0] f1244_wdata;
  logic [0:0] f1244_clk;
  logic [0:0] f1244_rst;
  logic [31:0] f1244_rdata;
  sr_buffer_32_1 f1244(.wen(f1244_wen), .wdata(f1244_wdata), .clk(f1244_clk), .rst(f1244_rst), .rdata(f1244_rdata));
  assign f1244_clk = clk;
  assign f1244_rst = rst;
  // Bindings to f1244

  // f1246
  logic [0:0] f1246_wen;
  logic [31:0] f1246_wdata;
  logic [0:0] f1246_clk;
  logic [0:0] f1246_rst;
  logic [31:0] f1246_rdata;
  sr_buffer_32_1 f1246(.wen(f1246_wen), .wdata(f1246_wdata), .clk(f1246_clk), .rst(f1246_rst), .rdata(f1246_rdata));
  assign f1246_clk = clk;
  assign f1246_rst = rst;
  // Bindings to f1246

  // f1248
  logic [0:0] f1248_wen;
  logic [31:0] f1248_wdata;
  logic [0:0] f1248_clk;
  logic [0:0] f1248_rst;
  logic [31:0] f1248_rdata;
  sr_buffer_32_1 f1248(.wen(f1248_wen), .wdata(f1248_wdata), .clk(f1248_clk), .rst(f1248_rst), .rdata(f1248_rdata));
  assign f1248_clk = clk;
  assign f1248_rst = rst;
  // Bindings to f1248

  // f1250
  logic [0:0] f1250_wen;
  logic [31:0] f1250_wdata;
  logic [0:0] f1250_clk;
  logic [0:0] f1250_rst;
  logic [31:0] f1250_rdata;
  sr_buffer_32_1 f1250(.wen(f1250_wen), .wdata(f1250_wdata), .clk(f1250_clk), .rst(f1250_rst), .rdata(f1250_rdata));
  assign f1250_clk = clk;
  assign f1250_rst = rst;
  // Bindings to f1250

  // f1252
  logic [0:0] f1252_wen;
  logic [31:0] f1252_wdata;
  logic [0:0] f1252_clk;
  logic [0:0] f1252_rst;
  logic [31:0] f1252_rdata;
  sr_buffer_32_1 f1252(.wen(f1252_wen), .wdata(f1252_wdata), .clk(f1252_clk), .rst(f1252_rst), .rdata(f1252_rdata));
  assign f1252_clk = clk;
  assign f1252_rst = rst;
  // Bindings to f1252

  // f1254
  logic [0:0] f1254_wen;
  logic [31:0] f1254_wdata;
  logic [0:0] f1254_clk;
  logic [0:0] f1254_rst;
  logic [31:0] f1254_rdata;
  sr_buffer_32_1 f1254(.wen(f1254_wen), .wdata(f1254_wdata), .clk(f1254_clk), .rst(f1254_rst), .rdata(f1254_rdata));
  assign f1254_clk = clk;
  assign f1254_rst = rst;
  // Bindings to f1254

  // f1256
  logic [0:0] f1256_wen;
  logic [31:0] f1256_wdata;
  logic [0:0] f1256_clk;
  logic [0:0] f1256_rst;
  logic [31:0] f1256_rdata;
  sr_buffer_32_1 f1256(.wen(f1256_wen), .wdata(f1256_wdata), .clk(f1256_clk), .rst(f1256_rst), .rdata(f1256_rdata));
  assign f1256_clk = clk;
  assign f1256_rst = rst;
  // Bindings to f1256

  // f1258
  logic [0:0] f1258_wen;
  logic [31:0] f1258_wdata;
  logic [0:0] f1258_clk;
  logic [0:0] f1258_rst;
  logic [31:0] f1258_rdata;
  sr_buffer_32_1 f1258(.wen(f1258_wen), .wdata(f1258_wdata), .clk(f1258_clk), .rst(f1258_rst), .rdata(f1258_rdata));
  assign f1258_clk = clk;
  assign f1258_rst = rst;
  // Bindings to f1258

  // f1260
  logic [0:0] f1260_wen;
  logic [31:0] f1260_wdata;
  logic [0:0] f1260_clk;
  logic [0:0] f1260_rst;
  logic [31:0] f1260_rdata;
  sr_buffer_32_1 f1260(.wen(f1260_wen), .wdata(f1260_wdata), .clk(f1260_clk), .rst(f1260_rst), .rdata(f1260_rdata));
  assign f1260_clk = clk;
  assign f1260_rst = rst;
  // Bindings to f1260

  // f1262
  logic [0:0] f1262_wen;
  logic [31:0] f1262_wdata;
  logic [0:0] f1262_clk;
  logic [0:0] f1262_rst;
  logic [31:0] f1262_rdata;
  sr_buffer_32_1 f1262(.wen(f1262_wen), .wdata(f1262_wdata), .clk(f1262_clk), .rst(f1262_rst), .rdata(f1262_rdata));
  assign f1262_clk = clk;
  assign f1262_rst = rst;
  // Bindings to f1262

  // f1264
  logic [0:0] f1264_wen;
  logic [31:0] f1264_wdata;
  logic [0:0] f1264_clk;
  logic [0:0] f1264_rst;
  logic [31:0] f1264_rdata;
  sr_buffer_32_1 f1264(.wen(f1264_wen), .wdata(f1264_wdata), .clk(f1264_clk), .rst(f1264_rst), .rdata(f1264_rdata));
  assign f1264_clk = clk;
  assign f1264_rst = rst;
  // Bindings to f1264

  // f1266
  logic [0:0] f1266_wen;
  logic [31:0] f1266_wdata;
  logic [0:0] f1266_clk;
  logic [0:0] f1266_rst;
  logic [31:0] f1266_rdata;
  sr_buffer_32_1 f1266(.wen(f1266_wen), .wdata(f1266_wdata), .clk(f1266_clk), .rst(f1266_rst), .rdata(f1266_rdata));
  assign f1266_clk = clk;
  assign f1266_rst = rst;
  // Bindings to f1266

  // f1268
  logic [0:0] f1268_wen;
  logic [31:0] f1268_wdata;
  logic [0:0] f1268_clk;
  logic [0:0] f1268_rst;
  logic [31:0] f1268_rdata;
  sr_buffer_32_1 f1268(.wen(f1268_wen), .wdata(f1268_wdata), .clk(f1268_clk), .rst(f1268_rst), .rdata(f1268_rdata));
  assign f1268_clk = clk;
  assign f1268_rst = rst;
  // Bindings to f1268

  // f1270
  logic [0:0] f1270_wen;
  logic [31:0] f1270_wdata;
  logic [0:0] f1270_clk;
  logic [0:0] f1270_rst;
  logic [31:0] f1270_rdata;
  sr_buffer_32_1 f1270(.wen(f1270_wen), .wdata(f1270_wdata), .clk(f1270_clk), .rst(f1270_rst), .rdata(f1270_rdata));
  assign f1270_clk = clk;
  assign f1270_rst = rst;
  // Bindings to f1270

  // f1272
  logic [0:0] f1272_wen;
  logic [31:0] f1272_wdata;
  logic [0:0] f1272_clk;
  logic [0:0] f1272_rst;
  logic [31:0] f1272_rdata;
  sr_buffer_32_1 f1272(.wen(f1272_wen), .wdata(f1272_wdata), .clk(f1272_clk), .rst(f1272_rst), .rdata(f1272_rdata));
  assign f1272_clk = clk;
  assign f1272_rst = rst;
  // Bindings to f1272

  // f1274
  logic [0:0] f1274_wen;
  logic [31:0] f1274_wdata;
  logic [0:0] f1274_clk;
  logic [0:0] f1274_rst;
  logic [31:0] f1274_rdata;
  sr_buffer_32_1 f1274(.wen(f1274_wen), .wdata(f1274_wdata), .clk(f1274_clk), .rst(f1274_rst), .rdata(f1274_rdata));
  assign f1274_clk = clk;
  assign f1274_rst = rst;
  // Bindings to f1274

  // f1276
  logic [0:0] f1276_wen;
  logic [31:0] f1276_wdata;
  logic [0:0] f1276_clk;
  logic [0:0] f1276_rst;
  logic [31:0] f1276_rdata;
  sr_buffer_32_1 f1276(.wen(f1276_wen), .wdata(f1276_wdata), .clk(f1276_clk), .rst(f1276_rst), .rdata(f1276_rdata));
  assign f1276_clk = clk;
  assign f1276_rst = rst;
  // Bindings to f1276

  // f1278
  logic [0:0] f1278_wen;
  logic [31:0] f1278_wdata;
  logic [0:0] f1278_clk;
  logic [0:0] f1278_rst;
  logic [31:0] f1278_rdata;
  sr_buffer_32_1 f1278(.wen(f1278_wen), .wdata(f1278_wdata), .clk(f1278_clk), .rst(f1278_rst), .rdata(f1278_rdata));
  assign f1278_clk = clk;
  assign f1278_rst = rst;
  // Bindings to f1278

  // f1280
  logic [0:0] f1280_wen;
  logic [31:0] f1280_wdata;
  logic [0:0] f1280_clk;
  logic [0:0] f1280_rst;
  logic [31:0] f1280_rdata;
  sr_buffer_32_1 f1280(.wen(f1280_wen), .wdata(f1280_wdata), .clk(f1280_clk), .rst(f1280_rst), .rdata(f1280_rdata));
  assign f1280_clk = clk;
  assign f1280_rst = rst;
  // Bindings to f1280

  // f1282
  logic [0:0] f1282_wen;
  logic [31:0] f1282_wdata;
  logic [0:0] f1282_clk;
  logic [0:0] f1282_rst;
  logic [31:0] f1282_rdata;
  sr_buffer_32_1 f1282(.wen(f1282_wen), .wdata(f1282_wdata), .clk(f1282_clk), .rst(f1282_rst), .rdata(f1282_rdata));
  assign f1282_clk = clk;
  assign f1282_rst = rst;
  // Bindings to f1282

  // f1284
  logic [0:0] f1284_wen;
  logic [31:0] f1284_wdata;
  logic [0:0] f1284_clk;
  logic [0:0] f1284_rst;
  logic [31:0] f1284_rdata;
  sr_buffer_32_1 f1284(.wen(f1284_wen), .wdata(f1284_wdata), .clk(f1284_clk), .rst(f1284_rst), .rdata(f1284_rdata));
  assign f1284_clk = clk;
  assign f1284_rst = rst;
  // Bindings to f1284

  // f1286
  logic [0:0] f1286_wen;
  logic [31:0] f1286_wdata;
  logic [0:0] f1286_clk;
  logic [0:0] f1286_rst;
  logic [31:0] f1286_rdata;
  sr_buffer_32_1 f1286(.wen(f1286_wen), .wdata(f1286_wdata), .clk(f1286_clk), .rst(f1286_rst), .rdata(f1286_rdata));
  assign f1286_clk = clk;
  assign f1286_rst = rst;
  // Bindings to f1286

  // f1288
  logic [0:0] f1288_wen;
  logic [31:0] f1288_wdata;
  logic [0:0] f1288_clk;
  logic [0:0] f1288_rst;
  logic [31:0] f1288_rdata;
  sr_buffer_32_1 f1288(.wen(f1288_wen), .wdata(f1288_wdata), .clk(f1288_clk), .rst(f1288_rst), .rdata(f1288_rdata));
  assign f1288_clk = clk;
  assign f1288_rst = rst;
  // Bindings to f1288

  // f1290
  logic [0:0] f1290_wen;
  logic [31:0] f1290_wdata;
  logic [0:0] f1290_clk;
  logic [0:0] f1290_rst;
  logic [31:0] f1290_rdata;
  sr_buffer_32_1 f1290(.wen(f1290_wen), .wdata(f1290_wdata), .clk(f1290_clk), .rst(f1290_rst), .rdata(f1290_rdata));
  assign f1290_clk = clk;
  assign f1290_rst = rst;
  // Bindings to f1290

  // f1292
  logic [0:0] f1292_wen;
  logic [31:0] f1292_wdata;
  logic [0:0] f1292_clk;
  logic [0:0] f1292_rst;
  logic [31:0] f1292_rdata;
  sr_buffer_32_1 f1292(.wen(f1292_wen), .wdata(f1292_wdata), .clk(f1292_clk), .rst(f1292_rst), .rdata(f1292_rdata));
  assign f1292_clk = clk;
  assign f1292_rst = rst;
  // Bindings to f1292

  // f1294
  logic [0:0] f1294_wen;
  logic [31:0] f1294_wdata;
  logic [0:0] f1294_clk;
  logic [0:0] f1294_rst;
  logic [31:0] f1294_rdata;
  sr_buffer_32_1 f1294(.wen(f1294_wen), .wdata(f1294_wdata), .clk(f1294_clk), .rst(f1294_rst), .rdata(f1294_rdata));
  assign f1294_clk = clk;
  assign f1294_rst = rst;
  // Bindings to f1294

  // f1296
  logic [0:0] f1296_wen;
  logic [31:0] f1296_wdata;
  logic [0:0] f1296_clk;
  logic [0:0] f1296_rst;
  logic [31:0] f1296_rdata;
  sr_buffer_32_1 f1296(.wen(f1296_wen), .wdata(f1296_wdata), .clk(f1296_clk), .rst(f1296_rst), .rdata(f1296_rdata));
  assign f1296_clk = clk;
  assign f1296_rst = rst;
  // Bindings to f1296

  // f1298
  logic [0:0] f1298_wen;
  logic [31:0] f1298_wdata;
  logic [0:0] f1298_clk;
  logic [0:0] f1298_rst;
  logic [31:0] f1298_rdata;
  sr_buffer_32_1 f1298(.wen(f1298_wen), .wdata(f1298_wdata), .clk(f1298_clk), .rst(f1298_rst), .rdata(f1298_rdata));
  assign f1298_clk = clk;
  assign f1298_rst = rst;
  // Bindings to f1298

  // f1300
  logic [0:0] f1300_wen;
  logic [31:0] f1300_wdata;
  logic [0:0] f1300_clk;
  logic [0:0] f1300_rst;
  logic [31:0] f1300_rdata;
  sr_buffer_32_1 f1300(.wen(f1300_wen), .wdata(f1300_wdata), .clk(f1300_clk), .rst(f1300_rst), .rdata(f1300_rdata));
  assign f1300_clk = clk;
  assign f1300_rst = rst;
  // Bindings to f1300

  // f1302
  logic [0:0] f1302_wen;
  logic [31:0] f1302_wdata;
  logic [0:0] f1302_clk;
  logic [0:0] f1302_rst;
  logic [31:0] f1302_rdata;
  sr_buffer_32_1 f1302(.wen(f1302_wen), .wdata(f1302_wdata), .clk(f1302_clk), .rst(f1302_rst), .rdata(f1302_rdata));
  assign f1302_clk = clk;
  assign f1302_rst = rst;
  // Bindings to f1302

  // f1304
  logic [0:0] f1304_wen;
  logic [31:0] f1304_wdata;
  logic [0:0] f1304_clk;
  logic [0:0] f1304_rst;
  logic [31:0] f1304_rdata;
  sr_buffer_32_1 f1304(.wen(f1304_wen), .wdata(f1304_wdata), .clk(f1304_clk), .rst(f1304_rst), .rdata(f1304_rdata));
  assign f1304_clk = clk;
  assign f1304_rst = rst;
  // Bindings to f1304

  // f1306
  logic [0:0] f1306_wen;
  logic [31:0] f1306_wdata;
  logic [0:0] f1306_clk;
  logic [0:0] f1306_rst;
  logic [31:0] f1306_rdata;
  sr_buffer_32_1 f1306(.wen(f1306_wen), .wdata(f1306_wdata), .clk(f1306_clk), .rst(f1306_rst), .rdata(f1306_rdata));
  assign f1306_clk = clk;
  assign f1306_rst = rst;
  // Bindings to f1306

  // f1308
  logic [0:0] f1308_wen;
  logic [31:0] f1308_wdata;
  logic [0:0] f1308_clk;
  logic [0:0] f1308_rst;
  logic [31:0] f1308_rdata;
  sr_buffer_32_1 f1308(.wen(f1308_wen), .wdata(f1308_wdata), .clk(f1308_clk), .rst(f1308_rst), .rdata(f1308_rdata));
  assign f1308_clk = clk;
  assign f1308_rst = rst;
  // Bindings to f1308

  // f1310
  logic [0:0] f1310_wen;
  logic [31:0] f1310_wdata;
  logic [0:0] f1310_clk;
  logic [0:0] f1310_rst;
  logic [31:0] f1310_rdata;
  sr_buffer_32_1 f1310(.wen(f1310_wen), .wdata(f1310_wdata), .clk(f1310_clk), .rst(f1310_rst), .rdata(f1310_rdata));
  assign f1310_clk = clk;
  assign f1310_rst = rst;
  // Bindings to f1310

  // f1312
  logic [0:0] f1312_wen;
  logic [31:0] f1312_wdata;
  logic [0:0] f1312_clk;
  logic [0:0] f1312_rst;
  logic [31:0] f1312_rdata;
  sr_buffer_32_1 f1312(.wen(f1312_wen), .wdata(f1312_wdata), .clk(f1312_clk), .rst(f1312_rst), .rdata(f1312_rdata));
  assign f1312_clk = clk;
  assign f1312_rst = rst;
  // Bindings to f1312

  // f1314
  logic [0:0] f1314_wen;
  logic [31:0] f1314_wdata;
  logic [0:0] f1314_clk;
  logic [0:0] f1314_rst;
  logic [31:0] f1314_rdata;
  sr_buffer_32_1 f1314(.wen(f1314_wen), .wdata(f1314_wdata), .clk(f1314_clk), .rst(f1314_rst), .rdata(f1314_rdata));
  assign f1314_clk = clk;
  assign f1314_rst = rst;
  // Bindings to f1314

  // f1316
  logic [0:0] f1316_wen;
  logic [31:0] f1316_wdata;
  logic [0:0] f1316_clk;
  logic [0:0] f1316_rst;
  logic [31:0] f1316_rdata;
  sr_buffer_32_1 f1316(.wen(f1316_wen), .wdata(f1316_wdata), .clk(f1316_clk), .rst(f1316_rst), .rdata(f1316_rdata));
  assign f1316_clk = clk;
  assign f1316_rst = rst;
  // Bindings to f1316

  // f1318
  logic [0:0] f1318_wen;
  logic [31:0] f1318_wdata;
  logic [0:0] f1318_clk;
  logic [0:0] f1318_rst;
  logic [31:0] f1318_rdata;
  sr_buffer_32_1 f1318(.wen(f1318_wen), .wdata(f1318_wdata), .clk(f1318_clk), .rst(f1318_rst), .rdata(f1318_rdata));
  assign f1318_clk = clk;
  assign f1318_rst = rst;
  // Bindings to f1318

  // f1320
  logic [0:0] f1320_wen;
  logic [31:0] f1320_wdata;
  logic [0:0] f1320_clk;
  logic [0:0] f1320_rst;
  logic [31:0] f1320_rdata;
  sr_buffer_32_1 f1320(.wen(f1320_wen), .wdata(f1320_wdata), .clk(f1320_clk), .rst(f1320_rst), .rdata(f1320_rdata));
  assign f1320_clk = clk;
  assign f1320_rst = rst;
  // Bindings to f1320

  // f1322
  logic [0:0] f1322_wen;
  logic [31:0] f1322_wdata;
  logic [0:0] f1322_clk;
  logic [0:0] f1322_rst;
  logic [31:0] f1322_rdata;
  sr_buffer_32_1 f1322(.wen(f1322_wen), .wdata(f1322_wdata), .clk(f1322_clk), .rst(f1322_rst), .rdata(f1322_rdata));
  assign f1322_clk = clk;
  assign f1322_rst = rst;
  // Bindings to f1322

  // f1324
  logic [0:0] f1324_wen;
  logic [31:0] f1324_wdata;
  logic [0:0] f1324_clk;
  logic [0:0] f1324_rst;
  logic [31:0] f1324_rdata;
  sr_buffer_32_1 f1324(.wen(f1324_wen), .wdata(f1324_wdata), .clk(f1324_clk), .rst(f1324_rst), .rdata(f1324_rdata));
  assign f1324_clk = clk;
  assign f1324_rst = rst;
  // Bindings to f1324

  // f1326
  logic [0:0] f1326_wen;
  logic [31:0] f1326_wdata;
  logic [0:0] f1326_clk;
  logic [0:0] f1326_rst;
  logic [31:0] f1326_rdata;
  sr_buffer_32_1 f1326(.wen(f1326_wen), .wdata(f1326_wdata), .clk(f1326_clk), .rst(f1326_rst), .rdata(f1326_rdata));
  assign f1326_clk = clk;
  assign f1326_rst = rst;
  // Bindings to f1326

  // f1328
  logic [0:0] f1328_wen;
  logic [31:0] f1328_wdata;
  logic [0:0] f1328_clk;
  logic [0:0] f1328_rst;
  logic [31:0] f1328_rdata;
  sr_buffer_32_1 f1328(.wen(f1328_wen), .wdata(f1328_wdata), .clk(f1328_clk), .rst(f1328_rst), .rdata(f1328_rdata));
  assign f1328_clk = clk;
  assign f1328_rst = rst;
  // Bindings to f1328

  // f1330
  logic [0:0] f1330_wen;
  logic [31:0] f1330_wdata;
  logic [0:0] f1330_clk;
  logic [0:0] f1330_rst;
  logic [31:0] f1330_rdata;
  sr_buffer_32_1 f1330(.wen(f1330_wen), .wdata(f1330_wdata), .clk(f1330_clk), .rst(f1330_rst), .rdata(f1330_rdata));
  assign f1330_clk = clk;
  assign f1330_rst = rst;
  // Bindings to f1330

  // f1332
  logic [0:0] f1332_wen;
  logic [31:0] f1332_wdata;
  logic [0:0] f1332_clk;
  logic [0:0] f1332_rst;
  logic [31:0] f1332_rdata;
  sr_buffer_32_1 f1332(.wen(f1332_wen), .wdata(f1332_wdata), .clk(f1332_clk), .rst(f1332_rst), .rdata(f1332_rdata));
  assign f1332_clk = clk;
  assign f1332_rst = rst;
  // Bindings to f1332

  // f1334
  logic [0:0] f1334_wen;
  logic [31:0] f1334_wdata;
  logic [0:0] f1334_clk;
  logic [0:0] f1334_rst;
  logic [31:0] f1334_rdata;
  sr_buffer_32_1 f1334(.wen(f1334_wen), .wdata(f1334_wdata), .clk(f1334_clk), .rst(f1334_rst), .rdata(f1334_rdata));
  assign f1334_clk = clk;
  assign f1334_rst = rst;
  // Bindings to f1334

  // f1336
  logic [0:0] f1336_wen;
  logic [31:0] f1336_wdata;
  logic [0:0] f1336_clk;
  logic [0:0] f1336_rst;
  logic [31:0] f1336_rdata;
  sr_buffer_32_1 f1336(.wen(f1336_wen), .wdata(f1336_wdata), .clk(f1336_clk), .rst(f1336_rst), .rdata(f1336_rdata));
  assign f1336_clk = clk;
  assign f1336_rst = rst;
  // Bindings to f1336

  // f1338
  logic [0:0] f1338_wen;
  logic [31:0] f1338_wdata;
  logic [0:0] f1338_clk;
  logic [0:0] f1338_rst;
  logic [31:0] f1338_rdata;
  sr_buffer_32_1 f1338(.wen(f1338_wen), .wdata(f1338_wdata), .clk(f1338_clk), .rst(f1338_rst), .rdata(f1338_rdata));
  assign f1338_clk = clk;
  assign f1338_rst = rst;
  // Bindings to f1338

  // f1340
  logic [0:0] f1340_wen;
  logic [31:0] f1340_wdata;
  logic [0:0] f1340_clk;
  logic [0:0] f1340_rst;
  logic [31:0] f1340_rdata;
  sr_buffer_32_1 f1340(.wen(f1340_wen), .wdata(f1340_wdata), .clk(f1340_clk), .rst(f1340_rst), .rdata(f1340_rdata));
  assign f1340_clk = clk;
  assign f1340_rst = rst;
  // Bindings to f1340

  // f1342
  logic [0:0] f1342_wen;
  logic [31:0] f1342_wdata;
  logic [0:0] f1342_clk;
  logic [0:0] f1342_rst;
  logic [31:0] f1342_rdata;
  sr_buffer_32_1 f1342(.wen(f1342_wen), .wdata(f1342_wdata), .clk(f1342_clk), .rst(f1342_rst), .rdata(f1342_rdata));
  assign f1342_clk = clk;
  assign f1342_rst = rst;
  // Bindings to f1342

  // f1344
  logic [0:0] f1344_wen;
  logic [31:0] f1344_wdata;
  logic [0:0] f1344_clk;
  logic [0:0] f1344_rst;
  logic [31:0] f1344_rdata;
  sr_buffer_32_1 f1344(.wen(f1344_wen), .wdata(f1344_wdata), .clk(f1344_clk), .rst(f1344_rst), .rdata(f1344_rdata));
  assign f1344_clk = clk;
  assign f1344_rst = rst;
  // Bindings to f1344

  // f1346
  logic [0:0] f1346_wen;
  logic [31:0] f1346_wdata;
  logic [0:0] f1346_clk;
  logic [0:0] f1346_rst;
  logic [31:0] f1346_rdata;
  sr_buffer_32_1 f1346(.wen(f1346_wen), .wdata(f1346_wdata), .clk(f1346_clk), .rst(f1346_rst), .rdata(f1346_rdata));
  assign f1346_clk = clk;
  assign f1346_rst = rst;
  // Bindings to f1346

  // f1348
  logic [0:0] f1348_wen;
  logic [31:0] f1348_wdata;
  logic [0:0] f1348_clk;
  logic [0:0] f1348_rst;
  logic [31:0] f1348_rdata;
  sr_buffer_32_1 f1348(.wen(f1348_wen), .wdata(f1348_wdata), .clk(f1348_clk), .rst(f1348_rst), .rdata(f1348_rdata));
  assign f1348_clk = clk;
  assign f1348_rst = rst;
  // Bindings to f1348

  // f1350
  logic [0:0] f1350_wen;
  logic [31:0] f1350_wdata;
  logic [0:0] f1350_clk;
  logic [0:0] f1350_rst;
  logic [31:0] f1350_rdata;
  sr_buffer_32_1 f1350(.wen(f1350_wen), .wdata(f1350_wdata), .clk(f1350_clk), .rst(f1350_rst), .rdata(f1350_rdata));
  assign f1350_clk = clk;
  assign f1350_rst = rst;
  // Bindings to f1350

  // f1352
  logic [0:0] f1352_wen;
  logic [31:0] f1352_wdata;
  logic [0:0] f1352_clk;
  logic [0:0] f1352_rst;
  logic [31:0] f1352_rdata;
  sr_buffer_32_1 f1352(.wen(f1352_wen), .wdata(f1352_wdata), .clk(f1352_clk), .rst(f1352_rst), .rdata(f1352_rdata));
  assign f1352_clk = clk;
  assign f1352_rst = rst;
  // Bindings to f1352

  // f1354
  logic [0:0] f1354_wen;
  logic [31:0] f1354_wdata;
  logic [0:0] f1354_clk;
  logic [0:0] f1354_rst;
  logic [31:0] f1354_rdata;
  sr_buffer_32_1 f1354(.wen(f1354_wen), .wdata(f1354_wdata), .clk(f1354_clk), .rst(f1354_rst), .rdata(f1354_rdata));
  assign f1354_clk = clk;
  assign f1354_rst = rst;
  // Bindings to f1354

  // f1356
  logic [0:0] f1356_wen;
  logic [31:0] f1356_wdata;
  logic [0:0] f1356_clk;
  logic [0:0] f1356_rst;
  logic [31:0] f1356_rdata;
  sr_buffer_32_1 f1356(.wen(f1356_wen), .wdata(f1356_wdata), .clk(f1356_clk), .rst(f1356_rst), .rdata(f1356_rdata));
  assign f1356_clk = clk;
  assign f1356_rst = rst;
  // Bindings to f1356

  // f1358
  logic [0:0] f1358_wen;
  logic [31:0] f1358_wdata;
  logic [0:0] f1358_clk;
  logic [0:0] f1358_rst;
  logic [31:0] f1358_rdata;
  sr_buffer_32_1 f1358(.wen(f1358_wen), .wdata(f1358_wdata), .clk(f1358_clk), .rst(f1358_rst), .rdata(f1358_rdata));
  assign f1358_clk = clk;
  assign f1358_rst = rst;
  // Bindings to f1358

  // f1360
  logic [0:0] f1360_wen;
  logic [31:0] f1360_wdata;
  logic [0:0] f1360_clk;
  logic [0:0] f1360_rst;
  logic [31:0] f1360_rdata;
  sr_buffer_32_1 f1360(.wen(f1360_wen), .wdata(f1360_wdata), .clk(f1360_clk), .rst(f1360_rst), .rdata(f1360_rdata));
  assign f1360_clk = clk;
  assign f1360_rst = rst;
  // Bindings to f1360

  // f1362
  logic [0:0] f1362_wen;
  logic [31:0] f1362_wdata;
  logic [0:0] f1362_clk;
  logic [0:0] f1362_rst;
  logic [31:0] f1362_rdata;
  sr_buffer_32_1 f1362(.wen(f1362_wen), .wdata(f1362_wdata), .clk(f1362_clk), .rst(f1362_rst), .rdata(f1362_rdata));
  assign f1362_clk = clk;
  assign f1362_rst = rst;
  // Bindings to f1362

  // f1364
  logic [0:0] f1364_wen;
  logic [31:0] f1364_wdata;
  logic [0:0] f1364_clk;
  logic [0:0] f1364_rst;
  logic [31:0] f1364_rdata;
  sr_buffer_32_1 f1364(.wen(f1364_wen), .wdata(f1364_wdata), .clk(f1364_clk), .rst(f1364_rst), .rdata(f1364_rdata));
  assign f1364_clk = clk;
  assign f1364_rst = rst;
  // Bindings to f1364

  // f1366
  logic [0:0] f1366_wen;
  logic [31:0] f1366_wdata;
  logic [0:0] f1366_clk;
  logic [0:0] f1366_rst;
  logic [31:0] f1366_rdata;
  sr_buffer_32_1 f1366(.wen(f1366_wen), .wdata(f1366_wdata), .clk(f1366_clk), .rst(f1366_rst), .rdata(f1366_rdata));
  assign f1366_clk = clk;
  assign f1366_rst = rst;
  // Bindings to f1366

  // f1368
  logic [0:0] f1368_wen;
  logic [31:0] f1368_wdata;
  logic [0:0] f1368_clk;
  logic [0:0] f1368_rst;
  logic [31:0] f1368_rdata;
  sr_buffer_32_1 f1368(.wen(f1368_wen), .wdata(f1368_wdata), .clk(f1368_clk), .rst(f1368_rst), .rdata(f1368_rdata));
  assign f1368_clk = clk;
  assign f1368_rst = rst;
  // Bindings to f1368

  // f1370
  logic [0:0] f1370_wen;
  logic [31:0] f1370_wdata;
  logic [0:0] f1370_clk;
  logic [0:0] f1370_rst;
  logic [31:0] f1370_rdata;
  sr_buffer_32_1 f1370(.wen(f1370_wen), .wdata(f1370_wdata), .clk(f1370_clk), .rst(f1370_rst), .rdata(f1370_rdata));
  assign f1370_clk = clk;
  assign f1370_rst = rst;
  // Bindings to f1370

  // f1372
  logic [0:0] f1372_wen;
  logic [31:0] f1372_wdata;
  logic [0:0] f1372_clk;
  logic [0:0] f1372_rst;
  logic [31:0] f1372_rdata;
  sr_buffer_32_1 f1372(.wen(f1372_wen), .wdata(f1372_wdata), .clk(f1372_clk), .rst(f1372_rst), .rdata(f1372_rdata));
  assign f1372_clk = clk;
  assign f1372_rst = rst;
  // Bindings to f1372

  // f1374
  logic [0:0] f1374_wen;
  logic [31:0] f1374_wdata;
  logic [0:0] f1374_clk;
  logic [0:0] f1374_rst;
  logic [31:0] f1374_rdata;
  sr_buffer_32_1 f1374(.wen(f1374_wen), .wdata(f1374_wdata), .clk(f1374_clk), .rst(f1374_rst), .rdata(f1374_rdata));
  assign f1374_clk = clk;
  assign f1374_rst = rst;
  // Bindings to f1374

  // f1376
  logic [0:0] f1376_wen;
  logic [31:0] f1376_wdata;
  logic [0:0] f1376_clk;
  logic [0:0] f1376_rst;
  logic [31:0] f1376_rdata;
  sr_buffer_32_1 f1376(.wen(f1376_wen), .wdata(f1376_wdata), .clk(f1376_clk), .rst(f1376_rst), .rdata(f1376_rdata));
  assign f1376_clk = clk;
  assign f1376_rst = rst;
  // Bindings to f1376

  // f1378
  logic [0:0] f1378_wen;
  logic [31:0] f1378_wdata;
  logic [0:0] f1378_clk;
  logic [0:0] f1378_rst;
  logic [31:0] f1378_rdata;
  sr_buffer_32_1 f1378(.wen(f1378_wen), .wdata(f1378_wdata), .clk(f1378_clk), .rst(f1378_rst), .rdata(f1378_rdata));
  assign f1378_clk = clk;
  assign f1378_rst = rst;
  // Bindings to f1378

  // f1380
  logic [0:0] f1380_wen;
  logic [31:0] f1380_wdata;
  logic [0:0] f1380_clk;
  logic [0:0] f1380_rst;
  logic [31:0] f1380_rdata;
  sr_buffer_32_1 f1380(.wen(f1380_wen), .wdata(f1380_wdata), .clk(f1380_clk), .rst(f1380_rst), .rdata(f1380_rdata));
  assign f1380_clk = clk;
  assign f1380_rst = rst;
  // Bindings to f1380

  // f1382
  logic [0:0] f1382_wen;
  logic [31:0] f1382_wdata;
  logic [0:0] f1382_clk;
  logic [0:0] f1382_rst;
  logic [31:0] f1382_rdata;
  sr_buffer_32_1 f1382(.wen(f1382_wen), .wdata(f1382_wdata), .clk(f1382_clk), .rst(f1382_rst), .rdata(f1382_rdata));
  assign f1382_clk = clk;
  assign f1382_rst = rst;
  // Bindings to f1382

  // f1384
  logic [0:0] f1384_wen;
  logic [31:0] f1384_wdata;
  logic [0:0] f1384_clk;
  logic [0:0] f1384_rst;
  logic [31:0] f1384_rdata;
  sr_buffer_32_1 f1384(.wen(f1384_wen), .wdata(f1384_wdata), .clk(f1384_clk), .rst(f1384_rst), .rdata(f1384_rdata));
  assign f1384_clk = clk;
  assign f1384_rst = rst;
  // Bindings to f1384

  // f1386
  logic [0:0] f1386_wen;
  logic [31:0] f1386_wdata;
  logic [0:0] f1386_clk;
  logic [0:0] f1386_rst;
  logic [31:0] f1386_rdata;
  sr_buffer_32_1 f1386(.wen(f1386_wen), .wdata(f1386_wdata), .clk(f1386_clk), .rst(f1386_rst), .rdata(f1386_rdata));
  assign f1386_clk = clk;
  assign f1386_rst = rst;
  // Bindings to f1386

  // f1388
  logic [0:0] f1388_wen;
  logic [31:0] f1388_wdata;
  logic [0:0] f1388_clk;
  logic [0:0] f1388_rst;
  logic [31:0] f1388_rdata;
  sr_buffer_32_1 f1388(.wen(f1388_wen), .wdata(f1388_wdata), .clk(f1388_clk), .rst(f1388_rst), .rdata(f1388_rdata));
  assign f1388_clk = clk;
  assign f1388_rst = rst;
  // Bindings to f1388

  // f1390
  logic [0:0] f1390_wen;
  logic [31:0] f1390_wdata;
  logic [0:0] f1390_clk;
  logic [0:0] f1390_rst;
  logic [31:0] f1390_rdata;
  sr_buffer_32_1 f1390(.wen(f1390_wen), .wdata(f1390_wdata), .clk(f1390_clk), .rst(f1390_rst), .rdata(f1390_rdata));
  assign f1390_clk = clk;
  assign f1390_rst = rst;
  // Bindings to f1390

  // f1392
  logic [0:0] f1392_wen;
  logic [31:0] f1392_wdata;
  logic [0:0] f1392_clk;
  logic [0:0] f1392_rst;
  logic [31:0] f1392_rdata;
  sr_buffer_32_1 f1392(.wen(f1392_wen), .wdata(f1392_wdata), .clk(f1392_clk), .rst(f1392_rst), .rdata(f1392_rdata));
  assign f1392_clk = clk;
  assign f1392_rst = rst;
  // Bindings to f1392

  // f1394
  logic [0:0] f1394_wen;
  logic [31:0] f1394_wdata;
  logic [0:0] f1394_clk;
  logic [0:0] f1394_rst;
  logic [31:0] f1394_rdata;
  sr_buffer_32_1 f1394(.wen(f1394_wen), .wdata(f1394_wdata), .clk(f1394_clk), .rst(f1394_rst), .rdata(f1394_rdata));
  assign f1394_clk = clk;
  assign f1394_rst = rst;
  // Bindings to f1394

  // f1396
  logic [0:0] f1396_wen;
  logic [31:0] f1396_wdata;
  logic [0:0] f1396_clk;
  logic [0:0] f1396_rst;
  logic [31:0] f1396_rdata;
  sr_buffer_32_1 f1396(.wen(f1396_wen), .wdata(f1396_wdata), .clk(f1396_clk), .rst(f1396_rst), .rdata(f1396_rdata));
  assign f1396_clk = clk;
  assign f1396_rst = rst;
  // Bindings to f1396

  // f1398
  logic [0:0] f1398_wen;
  logic [31:0] f1398_wdata;
  logic [0:0] f1398_clk;
  logic [0:0] f1398_rst;
  logic [31:0] f1398_rdata;
  sr_buffer_32_1 f1398(.wen(f1398_wen), .wdata(f1398_wdata), .clk(f1398_clk), .rst(f1398_rst), .rdata(f1398_rdata));
  assign f1398_clk = clk;
  assign f1398_rst = rst;
  // Bindings to f1398

  // f1400
  logic [0:0] f1400_wen;
  logic [31:0] f1400_wdata;
  logic [0:0] f1400_clk;
  logic [0:0] f1400_rst;
  logic [31:0] f1400_rdata;
  sr_buffer_32_1 f1400(.wen(f1400_wen), .wdata(f1400_wdata), .clk(f1400_clk), .rst(f1400_rst), .rdata(f1400_rdata));
  assign f1400_clk = clk;
  assign f1400_rst = rst;
  // Bindings to f1400

  // f1402
  logic [0:0] f1402_wen;
  logic [31:0] f1402_wdata;
  logic [0:0] f1402_clk;
  logic [0:0] f1402_rst;
  logic [31:0] f1402_rdata;
  sr_buffer_32_1 f1402(.wen(f1402_wen), .wdata(f1402_wdata), .clk(f1402_clk), .rst(f1402_rst), .rdata(f1402_rdata));
  assign f1402_clk = clk;
  assign f1402_rst = rst;
  // Bindings to f1402

  // f1404
  logic [0:0] f1404_wen;
  logic [31:0] f1404_wdata;
  logic [0:0] f1404_clk;
  logic [0:0] f1404_rst;
  logic [31:0] f1404_rdata;
  sr_buffer_32_1 f1404(.wen(f1404_wen), .wdata(f1404_wdata), .clk(f1404_clk), .rst(f1404_rst), .rdata(f1404_rdata));
  assign f1404_clk = clk;
  assign f1404_rst = rst;
  // Bindings to f1404

  // f1406
  logic [0:0] f1406_wen;
  logic [31:0] f1406_wdata;
  logic [0:0] f1406_clk;
  logic [0:0] f1406_rst;
  logic [31:0] f1406_rdata;
  sr_buffer_32_1 f1406(.wen(f1406_wen), .wdata(f1406_wdata), .clk(f1406_clk), .rst(f1406_rst), .rdata(f1406_rdata));
  assign f1406_clk = clk;
  assign f1406_rst = rst;
  // Bindings to f1406

  // f1408
  logic [0:0] f1408_wen;
  logic [31:0] f1408_wdata;
  logic [0:0] f1408_clk;
  logic [0:0] f1408_rst;
  logic [31:0] f1408_rdata;
  sr_buffer_32_1 f1408(.wen(f1408_wen), .wdata(f1408_wdata), .clk(f1408_clk), .rst(f1408_rst), .rdata(f1408_rdata));
  assign f1408_clk = clk;
  assign f1408_rst = rst;
  // Bindings to f1408

  // f1410
  logic [0:0] f1410_wen;
  logic [31:0] f1410_wdata;
  logic [0:0] f1410_clk;
  logic [0:0] f1410_rst;
  logic [31:0] f1410_rdata;
  sr_buffer_32_1 f1410(.wen(f1410_wen), .wdata(f1410_wdata), .clk(f1410_clk), .rst(f1410_rst), .rdata(f1410_rdata));
  assign f1410_clk = clk;
  assign f1410_rst = rst;
  // Bindings to f1410

  // f1412
  logic [0:0] f1412_wen;
  logic [31:0] f1412_wdata;
  logic [0:0] f1412_clk;
  logic [0:0] f1412_rst;
  logic [31:0] f1412_rdata;
  sr_buffer_32_1 f1412(.wen(f1412_wen), .wdata(f1412_wdata), .clk(f1412_clk), .rst(f1412_rst), .rdata(f1412_rdata));
  assign f1412_clk = clk;
  assign f1412_rst = rst;
  // Bindings to f1412

  // f1414
  logic [0:0] f1414_wen;
  logic [31:0] f1414_wdata;
  logic [0:0] f1414_clk;
  logic [0:0] f1414_rst;
  logic [31:0] f1414_rdata;
  sr_buffer_32_1 f1414(.wen(f1414_wen), .wdata(f1414_wdata), .clk(f1414_clk), .rst(f1414_rst), .rdata(f1414_rdata));
  assign f1414_clk = clk;
  assign f1414_rst = rst;
  // Bindings to f1414

  // f1416
  logic [0:0] f1416_wen;
  logic [31:0] f1416_wdata;
  logic [0:0] f1416_clk;
  logic [0:0] f1416_rst;
  logic [31:0] f1416_rdata;
  sr_buffer_32_1 f1416(.wen(f1416_wen), .wdata(f1416_wdata), .clk(f1416_clk), .rst(f1416_rst), .rdata(f1416_rdata));
  assign f1416_clk = clk;
  assign f1416_rst = rst;
  // Bindings to f1416

  // f1418
  logic [0:0] f1418_wen;
  logic [31:0] f1418_wdata;
  logic [0:0] f1418_clk;
  logic [0:0] f1418_rst;
  logic [31:0] f1418_rdata;
  sr_buffer_32_1 f1418(.wen(f1418_wen), .wdata(f1418_wdata), .clk(f1418_clk), .rst(f1418_rst), .rdata(f1418_rdata));
  assign f1418_clk = clk;
  assign f1418_rst = rst;
  // Bindings to f1418

  // f1420
  logic [0:0] f1420_wen;
  logic [31:0] f1420_wdata;
  logic [0:0] f1420_clk;
  logic [0:0] f1420_rst;
  logic [31:0] f1420_rdata;
  sr_buffer_32_1 f1420(.wen(f1420_wen), .wdata(f1420_wdata), .clk(f1420_clk), .rst(f1420_rst), .rdata(f1420_rdata));
  assign f1420_clk = clk;
  assign f1420_rst = rst;
  // Bindings to f1420

  // f1422
  logic [0:0] f1422_wen;
  logic [31:0] f1422_wdata;
  logic [0:0] f1422_clk;
  logic [0:0] f1422_rst;
  logic [31:0] f1422_rdata;
  sr_buffer_32_1 f1422(.wen(f1422_wen), .wdata(f1422_wdata), .clk(f1422_clk), .rst(f1422_rst), .rdata(f1422_rdata));
  assign f1422_clk = clk;
  assign f1422_rst = rst;
  // Bindings to f1422

  // f1424
  logic [0:0] f1424_wen;
  logic [31:0] f1424_wdata;
  logic [0:0] f1424_clk;
  logic [0:0] f1424_rst;
  logic [31:0] f1424_rdata;
  sr_buffer_32_1 f1424(.wen(f1424_wen), .wdata(f1424_wdata), .clk(f1424_clk), .rst(f1424_rst), .rdata(f1424_rdata));
  assign f1424_clk = clk;
  assign f1424_rst = rst;
  // Bindings to f1424

  // f1426
  logic [0:0] f1426_wen;
  logic [31:0] f1426_wdata;
  logic [0:0] f1426_clk;
  logic [0:0] f1426_rst;
  logic [31:0] f1426_rdata;
  sr_buffer_32_1 f1426(.wen(f1426_wen), .wdata(f1426_wdata), .clk(f1426_clk), .rst(f1426_rst), .rdata(f1426_rdata));
  assign f1426_clk = clk;
  assign f1426_rst = rst;
  // Bindings to f1426

  // f1428
  logic [0:0] f1428_wen;
  logic [31:0] f1428_wdata;
  logic [0:0] f1428_clk;
  logic [0:0] f1428_rst;
  logic [31:0] f1428_rdata;
  sr_buffer_32_1 f1428(.wen(f1428_wen), .wdata(f1428_wdata), .clk(f1428_clk), .rst(f1428_rst), .rdata(f1428_rdata));
  assign f1428_clk = clk;
  assign f1428_rst = rst;
  // Bindings to f1428

  // f1430
  logic [0:0] f1430_wen;
  logic [31:0] f1430_wdata;
  logic [0:0] f1430_clk;
  logic [0:0] f1430_rst;
  logic [31:0] f1430_rdata;
  sr_buffer_32_1 f1430(.wen(f1430_wen), .wdata(f1430_wdata), .clk(f1430_clk), .rst(f1430_rst), .rdata(f1430_rdata));
  assign f1430_clk = clk;
  assign f1430_rst = rst;
  // Bindings to f1430

  // f1432
  logic [0:0] f1432_wen;
  logic [31:0] f1432_wdata;
  logic [0:0] f1432_clk;
  logic [0:0] f1432_rst;
  logic [31:0] f1432_rdata;
  sr_buffer_32_1 f1432(.wen(f1432_wen), .wdata(f1432_wdata), .clk(f1432_clk), .rst(f1432_rst), .rdata(f1432_rdata));
  assign f1432_clk = clk;
  assign f1432_rst = rst;
  // Bindings to f1432

  // f1434
  logic [0:0] f1434_wen;
  logic [31:0] f1434_wdata;
  logic [0:0] f1434_clk;
  logic [0:0] f1434_rst;
  logic [31:0] f1434_rdata;
  sr_buffer_32_1 f1434(.wen(f1434_wen), .wdata(f1434_wdata), .clk(f1434_clk), .rst(f1434_rst), .rdata(f1434_rdata));
  assign f1434_clk = clk;
  assign f1434_rst = rst;
  // Bindings to f1434

  // f1436
  logic [0:0] f1436_wen;
  logic [31:0] f1436_wdata;
  logic [0:0] f1436_clk;
  logic [0:0] f1436_rst;
  logic [31:0] f1436_rdata;
  sr_buffer_32_1 f1436(.wen(f1436_wen), .wdata(f1436_wdata), .clk(f1436_clk), .rst(f1436_rst), .rdata(f1436_rdata));
  assign f1436_clk = clk;
  assign f1436_rst = rst;
  // Bindings to f1436

  // f1438
  logic [0:0] f1438_wen;
  logic [31:0] f1438_wdata;
  logic [0:0] f1438_clk;
  logic [0:0] f1438_rst;
  logic [31:0] f1438_rdata;
  sr_buffer_32_1 f1438(.wen(f1438_wen), .wdata(f1438_wdata), .clk(f1438_clk), .rst(f1438_rst), .rdata(f1438_rdata));
  assign f1438_clk = clk;
  assign f1438_rst = rst;
  // Bindings to f1438

  // f1440
  logic [0:0] f1440_wen;
  logic [31:0] f1440_wdata;
  logic [0:0] f1440_clk;
  logic [0:0] f1440_rst;
  logic [31:0] f1440_rdata;
  sr_buffer_32_1 f1440(.wen(f1440_wen), .wdata(f1440_wdata), .clk(f1440_clk), .rst(f1440_rst), .rdata(f1440_rdata));
  assign f1440_clk = clk;
  assign f1440_rst = rst;
  // Bindings to f1440

  // f1442
  logic [0:0] f1442_wen;
  logic [31:0] f1442_wdata;
  logic [0:0] f1442_clk;
  logic [0:0] f1442_rst;
  logic [31:0] f1442_rdata;
  sr_buffer_32_1 f1442(.wen(f1442_wen), .wdata(f1442_wdata), .clk(f1442_clk), .rst(f1442_rst), .rdata(f1442_rdata));
  assign f1442_clk = clk;
  assign f1442_rst = rst;
  // Bindings to f1442

  // f1444
  logic [0:0] f1444_wen;
  logic [31:0] f1444_wdata;
  logic [0:0] f1444_clk;
  logic [0:0] f1444_rst;
  logic [31:0] f1444_rdata;
  sr_buffer_32_1 f1444(.wen(f1444_wen), .wdata(f1444_wdata), .clk(f1444_clk), .rst(f1444_rst), .rdata(f1444_rdata));
  assign f1444_clk = clk;
  assign f1444_rst = rst;
  // Bindings to f1444

  // f1446
  logic [0:0] f1446_wen;
  logic [31:0] f1446_wdata;
  logic [0:0] f1446_clk;
  logic [0:0] f1446_rst;
  logic [31:0] f1446_rdata;
  sr_buffer_32_1 f1446(.wen(f1446_wen), .wdata(f1446_wdata), .clk(f1446_clk), .rst(f1446_rst), .rdata(f1446_rdata));
  assign f1446_clk = clk;
  assign f1446_rst = rst;
  // Bindings to f1446

  // f1448
  logic [0:0] f1448_wen;
  logic [31:0] f1448_wdata;
  logic [0:0] f1448_clk;
  logic [0:0] f1448_rst;
  logic [31:0] f1448_rdata;
  sr_buffer_32_1 f1448(.wen(f1448_wen), .wdata(f1448_wdata), .clk(f1448_clk), .rst(f1448_rst), .rdata(f1448_rdata));
  assign f1448_clk = clk;
  assign f1448_rst = rst;
  // Bindings to f1448

  // f1450
  logic [0:0] f1450_wen;
  logic [31:0] f1450_wdata;
  logic [0:0] f1450_clk;
  logic [0:0] f1450_rst;
  logic [31:0] f1450_rdata;
  sr_buffer_32_1 f1450(.wen(f1450_wen), .wdata(f1450_wdata), .clk(f1450_clk), .rst(f1450_rst), .rdata(f1450_rdata));
  assign f1450_clk = clk;
  assign f1450_rst = rst;
  // Bindings to f1450

  // f1452
  logic [0:0] f1452_wen;
  logic [31:0] f1452_wdata;
  logic [0:0] f1452_clk;
  logic [0:0] f1452_rst;
  logic [31:0] f1452_rdata;
  sr_buffer_32_1 f1452(.wen(f1452_wen), .wdata(f1452_wdata), .clk(f1452_clk), .rst(f1452_rst), .rdata(f1452_rdata));
  assign f1452_clk = clk;
  assign f1452_rst = rst;
  // Bindings to f1452

  // f1454
  logic [0:0] f1454_wen;
  logic [31:0] f1454_wdata;
  logic [0:0] f1454_clk;
  logic [0:0] f1454_rst;
  logic [31:0] f1454_rdata;
  sr_buffer_32_1 f1454(.wen(f1454_wen), .wdata(f1454_wdata), .clk(f1454_clk), .rst(f1454_rst), .rdata(f1454_rdata));
  assign f1454_clk = clk;
  assign f1454_rst = rst;
  // Bindings to f1454

  // f1456
  logic [0:0] f1456_wen;
  logic [31:0] f1456_wdata;
  logic [0:0] f1456_clk;
  logic [0:0] f1456_rst;
  logic [31:0] f1456_rdata;
  sr_buffer_32_1 f1456(.wen(f1456_wen), .wdata(f1456_wdata), .clk(f1456_clk), .rst(f1456_rst), .rdata(f1456_rdata));
  assign f1456_clk = clk;
  assign f1456_rst = rst;
  // Bindings to f1456

  // f1458
  logic [0:0] f1458_wen;
  logic [31:0] f1458_wdata;
  logic [0:0] f1458_clk;
  logic [0:0] f1458_rst;
  logic [31:0] f1458_rdata;
  sr_buffer_32_1 f1458(.wen(f1458_wen), .wdata(f1458_wdata), .clk(f1458_clk), .rst(f1458_rst), .rdata(f1458_rdata));
  assign f1458_clk = clk;
  assign f1458_rst = rst;
  // Bindings to f1458

  // f1460
  logic [0:0] f1460_wen;
  logic [31:0] f1460_wdata;
  logic [0:0] f1460_clk;
  logic [0:0] f1460_rst;
  logic [31:0] f1460_rdata;
  sr_buffer_32_1 f1460(.wen(f1460_wen), .wdata(f1460_wdata), .clk(f1460_clk), .rst(f1460_rst), .rdata(f1460_rdata));
  assign f1460_clk = clk;
  assign f1460_rst = rst;
  // Bindings to f1460

  // f1462
  logic [0:0] f1462_wen;
  logic [31:0] f1462_wdata;
  logic [0:0] f1462_clk;
  logic [0:0] f1462_rst;
  logic [31:0] f1462_rdata;
  sr_buffer_32_1 f1462(.wen(f1462_wen), .wdata(f1462_wdata), .clk(f1462_clk), .rst(f1462_rst), .rdata(f1462_rdata));
  assign f1462_clk = clk;
  assign f1462_rst = rst;
  // Bindings to f1462

  // f1464
  logic [0:0] f1464_wen;
  logic [31:0] f1464_wdata;
  logic [0:0] f1464_clk;
  logic [0:0] f1464_rst;
  logic [31:0] f1464_rdata;
  sr_buffer_32_1 f1464(.wen(f1464_wen), .wdata(f1464_wdata), .clk(f1464_clk), .rst(f1464_rst), .rdata(f1464_rdata));
  assign f1464_clk = clk;
  assign f1464_rst = rst;
  // Bindings to f1464

  // f1466
  logic [0:0] f1466_wen;
  logic [31:0] f1466_wdata;
  logic [0:0] f1466_clk;
  logic [0:0] f1466_rst;
  logic [31:0] f1466_rdata;
  sr_buffer_32_1 f1466(.wen(f1466_wen), .wdata(f1466_wdata), .clk(f1466_clk), .rst(f1466_rst), .rdata(f1466_rdata));
  assign f1466_clk = clk;
  assign f1466_rst = rst;
  // Bindings to f1466

  // f1468
  logic [0:0] f1468_wen;
  logic [31:0] f1468_wdata;
  logic [0:0] f1468_clk;
  logic [0:0] f1468_rst;
  logic [31:0] f1468_rdata;
  sr_buffer_32_1 f1468(.wen(f1468_wen), .wdata(f1468_wdata), .clk(f1468_clk), .rst(f1468_rst), .rdata(f1468_rdata));
  assign f1468_clk = clk;
  assign f1468_rst = rst;
  // Bindings to f1468

  // f1470
  logic [0:0] f1470_wen;
  logic [31:0] f1470_wdata;
  logic [0:0] f1470_clk;
  logic [0:0] f1470_rst;
  logic [31:0] f1470_rdata;
  sr_buffer_32_1 f1470(.wen(f1470_wen), .wdata(f1470_wdata), .clk(f1470_clk), .rst(f1470_rst), .rdata(f1470_rdata));
  assign f1470_clk = clk;
  assign f1470_rst = rst;
  // Bindings to f1470

  // f1472
  logic [0:0] f1472_wen;
  logic [31:0] f1472_wdata;
  logic [0:0] f1472_clk;
  logic [0:0] f1472_rst;
  logic [31:0] f1472_rdata;
  sr_buffer_32_1 f1472(.wen(f1472_wen), .wdata(f1472_wdata), .clk(f1472_clk), .rst(f1472_rst), .rdata(f1472_rdata));
  assign f1472_clk = clk;
  assign f1472_rst = rst;
  // Bindings to f1472

  // f1474
  logic [0:0] f1474_wen;
  logic [31:0] f1474_wdata;
  logic [0:0] f1474_clk;
  logic [0:0] f1474_rst;
  logic [31:0] f1474_rdata;
  sr_buffer_32_1 f1474(.wen(f1474_wen), .wdata(f1474_wdata), .clk(f1474_clk), .rst(f1474_rst), .rdata(f1474_rdata));
  assign f1474_clk = clk;
  assign f1474_rst = rst;
  // Bindings to f1474

  // f1476
  logic [0:0] f1476_wen;
  logic [31:0] f1476_wdata;
  logic [0:0] f1476_clk;
  logic [0:0] f1476_rst;
  logic [31:0] f1476_rdata;
  sr_buffer_32_1 f1476(.wen(f1476_wen), .wdata(f1476_wdata), .clk(f1476_clk), .rst(f1476_rst), .rdata(f1476_rdata));
  assign f1476_clk = clk;
  assign f1476_rst = rst;
  // Bindings to f1476

  // f1478
  logic [0:0] f1478_wen;
  logic [31:0] f1478_wdata;
  logic [0:0] f1478_clk;
  logic [0:0] f1478_rst;
  logic [31:0] f1478_rdata;
  sr_buffer_32_1 f1478(.wen(f1478_wen), .wdata(f1478_wdata), .clk(f1478_clk), .rst(f1478_rst), .rdata(f1478_rdata));
  assign f1478_clk = clk;
  assign f1478_rst = rst;
  // Bindings to f1478

  // f1480
  logic [0:0] f1480_wen;
  logic [31:0] f1480_wdata;
  logic [0:0] f1480_clk;
  logic [0:0] f1480_rst;
  logic [31:0] f1480_rdata;
  sr_buffer_32_1 f1480(.wen(f1480_wen), .wdata(f1480_wdata), .clk(f1480_clk), .rst(f1480_rst), .rdata(f1480_rdata));
  assign f1480_clk = clk;
  assign f1480_rst = rst;
  // Bindings to f1480

  // f1482
  logic [0:0] f1482_wen;
  logic [31:0] f1482_wdata;
  logic [0:0] f1482_clk;
  logic [0:0] f1482_rst;
  logic [31:0] f1482_rdata;
  sr_buffer_32_1 f1482(.wen(f1482_wen), .wdata(f1482_wdata), .clk(f1482_clk), .rst(f1482_rst), .rdata(f1482_rdata));
  assign f1482_clk = clk;
  assign f1482_rst = rst;
  // Bindings to f1482

  // f1484
  logic [0:0] f1484_wen;
  logic [31:0] f1484_wdata;
  logic [0:0] f1484_clk;
  logic [0:0] f1484_rst;
  logic [31:0] f1484_rdata;
  sr_buffer_32_1 f1484(.wen(f1484_wen), .wdata(f1484_wdata), .clk(f1484_clk), .rst(f1484_rst), .rdata(f1484_rdata));
  assign f1484_clk = clk;
  assign f1484_rst = rst;
  // Bindings to f1484

  // f1486
  logic [0:0] f1486_wen;
  logic [31:0] f1486_wdata;
  logic [0:0] f1486_clk;
  logic [0:0] f1486_rst;
  logic [31:0] f1486_rdata;
  sr_buffer_32_1 f1486(.wen(f1486_wen), .wdata(f1486_wdata), .clk(f1486_clk), .rst(f1486_rst), .rdata(f1486_rdata));
  assign f1486_clk = clk;
  assign f1486_rst = rst;
  // Bindings to f1486

  // f1488
  logic [0:0] f1488_wen;
  logic [31:0] f1488_wdata;
  logic [0:0] f1488_clk;
  logic [0:0] f1488_rst;
  logic [31:0] f1488_rdata;
  sr_buffer_32_1 f1488(.wen(f1488_wen), .wdata(f1488_wdata), .clk(f1488_clk), .rst(f1488_rst), .rdata(f1488_rdata));
  assign f1488_clk = clk;
  assign f1488_rst = rst;
  // Bindings to f1488

  // f1490
  logic [0:0] f1490_wen;
  logic [31:0] f1490_wdata;
  logic [0:0] f1490_clk;
  logic [0:0] f1490_rst;
  logic [31:0] f1490_rdata;
  sr_buffer_32_1 f1490(.wen(f1490_wen), .wdata(f1490_wdata), .clk(f1490_clk), .rst(f1490_rst), .rdata(f1490_rdata));
  assign f1490_clk = clk;
  assign f1490_rst = rst;
  // Bindings to f1490

  // f1492
  logic [0:0] f1492_wen;
  logic [31:0] f1492_wdata;
  logic [0:0] f1492_clk;
  logic [0:0] f1492_rst;
  logic [31:0] f1492_rdata;
  sr_buffer_32_1 f1492(.wen(f1492_wen), .wdata(f1492_wdata), .clk(f1492_clk), .rst(f1492_rst), .rdata(f1492_rdata));
  assign f1492_clk = clk;
  assign f1492_rst = rst;
  // Bindings to f1492

  // f1494
  logic [0:0] f1494_wen;
  logic [31:0] f1494_wdata;
  logic [0:0] f1494_clk;
  logic [0:0] f1494_rst;
  logic [31:0] f1494_rdata;
  sr_buffer_32_1 f1494(.wen(f1494_wen), .wdata(f1494_wdata), .clk(f1494_clk), .rst(f1494_rst), .rdata(f1494_rdata));
  assign f1494_clk = clk;
  assign f1494_rst = rst;
  // Bindings to f1494

  // f1496
  logic [0:0] f1496_wen;
  logic [31:0] f1496_wdata;
  logic [0:0] f1496_clk;
  logic [0:0] f1496_rst;
  logic [31:0] f1496_rdata;
  sr_buffer_32_1 f1496(.wen(f1496_wen), .wdata(f1496_wdata), .clk(f1496_clk), .rst(f1496_rst), .rdata(f1496_rdata));
  assign f1496_clk = clk;
  assign f1496_rst = rst;
  // Bindings to f1496

  // f1498
  logic [0:0] f1498_wen;
  logic [31:0] f1498_wdata;
  logic [0:0] f1498_clk;
  logic [0:0] f1498_rst;
  logic [31:0] f1498_rdata;
  sr_buffer_32_1 f1498(.wen(f1498_wen), .wdata(f1498_wdata), .clk(f1498_clk), .rst(f1498_rst), .rdata(f1498_rdata));
  assign f1498_clk = clk;
  assign f1498_rst = rst;
  // Bindings to f1498

  // f1500
  logic [0:0] f1500_wen;
  logic [31:0] f1500_wdata;
  logic [0:0] f1500_clk;
  logic [0:0] f1500_rst;
  logic [31:0] f1500_rdata;
  sr_buffer_32_1 f1500(.wen(f1500_wen), .wdata(f1500_wdata), .clk(f1500_clk), .rst(f1500_rst), .rdata(f1500_rdata));
  assign f1500_clk = clk;
  assign f1500_rst = rst;
  // Bindings to f1500

  // f1502
  logic [0:0] f1502_wen;
  logic [31:0] f1502_wdata;
  logic [0:0] f1502_clk;
  logic [0:0] f1502_rst;
  logic [31:0] f1502_rdata;
  sr_buffer_32_1 f1502(.wen(f1502_wen), .wdata(f1502_wdata), .clk(f1502_clk), .rst(f1502_rst), .rdata(f1502_rdata));
  assign f1502_clk = clk;
  assign f1502_rst = rst;
  // Bindings to f1502

  // f1504
  logic [0:0] f1504_wen;
  logic [31:0] f1504_wdata;
  logic [0:0] f1504_clk;
  logic [0:0] f1504_rst;
  logic [31:0] f1504_rdata;
  sr_buffer_32_1 f1504(.wen(f1504_wen), .wdata(f1504_wdata), .clk(f1504_clk), .rst(f1504_rst), .rdata(f1504_rdata));
  assign f1504_clk = clk;
  assign f1504_rst = rst;
  // Bindings to f1504

  // f1506
  logic [0:0] f1506_wen;
  logic [31:0] f1506_wdata;
  logic [0:0] f1506_clk;
  logic [0:0] f1506_rst;
  logic [31:0] f1506_rdata;
  sr_buffer_32_1 f1506(.wen(f1506_wen), .wdata(f1506_wdata), .clk(f1506_clk), .rst(f1506_rst), .rdata(f1506_rdata));
  assign f1506_clk = clk;
  assign f1506_rst = rst;
  // Bindings to f1506

  // f1508
  logic [0:0] f1508_wen;
  logic [31:0] f1508_wdata;
  logic [0:0] f1508_clk;
  logic [0:0] f1508_rst;
  logic [31:0] f1508_rdata;
  sr_buffer_32_1 f1508(.wen(f1508_wen), .wdata(f1508_wdata), .clk(f1508_clk), .rst(f1508_rst), .rdata(f1508_rdata));
  assign f1508_clk = clk;
  assign f1508_rst = rst;
  // Bindings to f1508

  // f1510
  logic [0:0] f1510_wen;
  logic [31:0] f1510_wdata;
  logic [0:0] f1510_clk;
  logic [0:0] f1510_rst;
  logic [31:0] f1510_rdata;
  sr_buffer_32_1 f1510(.wen(f1510_wen), .wdata(f1510_wdata), .clk(f1510_clk), .rst(f1510_rst), .rdata(f1510_rdata));
  assign f1510_clk = clk;
  assign f1510_rst = rst;
  // Bindings to f1510

  // f1512
  logic [0:0] f1512_wen;
  logic [31:0] f1512_wdata;
  logic [0:0] f1512_clk;
  logic [0:0] f1512_rst;
  logic [31:0] f1512_rdata;
  sr_buffer_32_1 f1512(.wen(f1512_wen), .wdata(f1512_wdata), .clk(f1512_clk), .rst(f1512_rst), .rdata(f1512_rdata));
  assign f1512_clk = clk;
  assign f1512_rst = rst;
  // Bindings to f1512

  // f1514
  logic [0:0] f1514_wen;
  logic [31:0] f1514_wdata;
  logic [0:0] f1514_clk;
  logic [0:0] f1514_rst;
  logic [31:0] f1514_rdata;
  sr_buffer_32_1 f1514(.wen(f1514_wen), .wdata(f1514_wdata), .clk(f1514_clk), .rst(f1514_rst), .rdata(f1514_rdata));
  assign f1514_clk = clk;
  assign f1514_rst = rst;
  // Bindings to f1514

  // f1516
  logic [0:0] f1516_wen;
  logic [31:0] f1516_wdata;
  logic [0:0] f1516_clk;
  logic [0:0] f1516_rst;
  logic [31:0] f1516_rdata;
  sr_buffer_32_1 f1516(.wen(f1516_wen), .wdata(f1516_wdata), .clk(f1516_clk), .rst(f1516_rst), .rdata(f1516_rdata));
  assign f1516_clk = clk;
  assign f1516_rst = rst;
  // Bindings to f1516

  // f1518
  logic [0:0] f1518_wen;
  logic [31:0] f1518_wdata;
  logic [0:0] f1518_clk;
  logic [0:0] f1518_rst;
  logic [31:0] f1518_rdata;
  sr_buffer_32_1 f1518(.wen(f1518_wen), .wdata(f1518_wdata), .clk(f1518_clk), .rst(f1518_rst), .rdata(f1518_rdata));
  assign f1518_clk = clk;
  assign f1518_rst = rst;
  // Bindings to f1518

  // f1520
  logic [0:0] f1520_wen;
  logic [31:0] f1520_wdata;
  logic [0:0] f1520_clk;
  logic [0:0] f1520_rst;
  logic [31:0] f1520_rdata;
  sr_buffer_32_1 f1520(.wen(f1520_wen), .wdata(f1520_wdata), .clk(f1520_clk), .rst(f1520_rst), .rdata(f1520_rdata));
  assign f1520_clk = clk;
  assign f1520_rst = rst;
  // Bindings to f1520

  // f1522
  logic [0:0] f1522_wen;
  logic [31:0] f1522_wdata;
  logic [0:0] f1522_clk;
  logic [0:0] f1522_rst;
  logic [31:0] f1522_rdata;
  sr_buffer_32_1 f1522(.wen(f1522_wen), .wdata(f1522_wdata), .clk(f1522_clk), .rst(f1522_rst), .rdata(f1522_rdata));
  assign f1522_clk = clk;
  assign f1522_rst = rst;
  // Bindings to f1522

  // f1524
  logic [0:0] f1524_wen;
  logic [31:0] f1524_wdata;
  logic [0:0] f1524_clk;
  logic [0:0] f1524_rst;
  logic [31:0] f1524_rdata;
  sr_buffer_32_1 f1524(.wen(f1524_wen), .wdata(f1524_wdata), .clk(f1524_clk), .rst(f1524_rst), .rdata(f1524_rdata));
  assign f1524_clk = clk;
  assign f1524_rst = rst;
  // Bindings to f1524

  // f1526
  logic [0:0] f1526_wen;
  logic [31:0] f1526_wdata;
  logic [0:0] f1526_clk;
  logic [0:0] f1526_rst;
  logic [31:0] f1526_rdata;
  sr_buffer_32_1 f1526(.wen(f1526_wen), .wdata(f1526_wdata), .clk(f1526_clk), .rst(f1526_rst), .rdata(f1526_rdata));
  assign f1526_clk = clk;
  assign f1526_rst = rst;
  // Bindings to f1526

  // f1528
  logic [0:0] f1528_wen;
  logic [31:0] f1528_wdata;
  logic [0:0] f1528_clk;
  logic [0:0] f1528_rst;
  logic [31:0] f1528_rdata;
  sr_buffer_32_1 f1528(.wen(f1528_wen), .wdata(f1528_wdata), .clk(f1528_clk), .rst(f1528_rst), .rdata(f1528_rdata));
  assign f1528_clk = clk;
  assign f1528_rst = rst;
  // Bindings to f1528

  // f1530
  logic [0:0] f1530_wen;
  logic [31:0] f1530_wdata;
  logic [0:0] f1530_clk;
  logic [0:0] f1530_rst;
  logic [31:0] f1530_rdata;
  sr_buffer_32_1 f1530(.wen(f1530_wen), .wdata(f1530_wdata), .clk(f1530_clk), .rst(f1530_rst), .rdata(f1530_rdata));
  assign f1530_clk = clk;
  assign f1530_rst = rst;
  // Bindings to f1530

  // f1532
  logic [0:0] f1532_wen;
  logic [31:0] f1532_wdata;
  logic [0:0] f1532_clk;
  logic [0:0] f1532_rst;
  logic [31:0] f1532_rdata;
  sr_buffer_32_1 f1532(.wen(f1532_wen), .wdata(f1532_wdata), .clk(f1532_clk), .rst(f1532_rst), .rdata(f1532_rdata));
  assign f1532_clk = clk;
  assign f1532_rst = rst;
  // Bindings to f1532

  // f1534
  logic [0:0] f1534_wen;
  logic [31:0] f1534_wdata;
  logic [0:0] f1534_clk;
  logic [0:0] f1534_rst;
  logic [31:0] f1534_rdata;
  sr_buffer_32_1 f1534(.wen(f1534_wen), .wdata(f1534_wdata), .clk(f1534_clk), .rst(f1534_rst), .rdata(f1534_rdata));
  assign f1534_clk = clk;
  assign f1534_rst = rst;
  // Bindings to f1534

  // f1536
  logic [0:0] f1536_wen;
  logic [31:0] f1536_wdata;
  logic [0:0] f1536_clk;
  logic [0:0] f1536_rst;
  logic [31:0] f1536_rdata;
  sr_buffer_32_1 f1536(.wen(f1536_wen), .wdata(f1536_wdata), .clk(f1536_clk), .rst(f1536_rst), .rdata(f1536_rdata));
  assign f1536_clk = clk;
  assign f1536_rst = rst;
  // Bindings to f1536

  // f1538
  logic [0:0] f1538_wen;
  logic [31:0] f1538_wdata;
  logic [0:0] f1538_clk;
  logic [0:0] f1538_rst;
  logic [31:0] f1538_rdata;
  sr_buffer_32_1 f1538(.wen(f1538_wen), .wdata(f1538_wdata), .clk(f1538_clk), .rst(f1538_rst), .rdata(f1538_rdata));
  assign f1538_clk = clk;
  assign f1538_rst = rst;
  // Bindings to f1538

  // f1540
  logic [0:0] f1540_wen;
  logic [31:0] f1540_wdata;
  logic [0:0] f1540_clk;
  logic [0:0] f1540_rst;
  logic [31:0] f1540_rdata;
  sr_buffer_32_1 f1540(.wen(f1540_wen), .wdata(f1540_wdata), .clk(f1540_clk), .rst(f1540_rst), .rdata(f1540_rdata));
  assign f1540_clk = clk;
  assign f1540_rst = rst;
  // Bindings to f1540

  // f1542
  logic [0:0] f1542_wen;
  logic [31:0] f1542_wdata;
  logic [0:0] f1542_clk;
  logic [0:0] f1542_rst;
  logic [31:0] f1542_rdata;
  sr_buffer_32_1 f1542(.wen(f1542_wen), .wdata(f1542_wdata), .clk(f1542_clk), .rst(f1542_rst), .rdata(f1542_rdata));
  assign f1542_clk = clk;
  assign f1542_rst = rst;
  // Bindings to f1542

  // f1544
  logic [0:0] f1544_wen;
  logic [31:0] f1544_wdata;
  logic [0:0] f1544_clk;
  logic [0:0] f1544_rst;
  logic [31:0] f1544_rdata;
  sr_buffer_32_1 f1544(.wen(f1544_wen), .wdata(f1544_wdata), .clk(f1544_clk), .rst(f1544_rst), .rdata(f1544_rdata));
  assign f1544_clk = clk;
  assign f1544_rst = rst;
  // Bindings to f1544

  // f1546
  logic [0:0] f1546_wen;
  logic [31:0] f1546_wdata;
  logic [0:0] f1546_clk;
  logic [0:0] f1546_rst;
  logic [31:0] f1546_rdata;
  sr_buffer_32_1 f1546(.wen(f1546_wen), .wdata(f1546_wdata), .clk(f1546_clk), .rst(f1546_rst), .rdata(f1546_rdata));
  assign f1546_clk = clk;
  assign f1546_rst = rst;
  // Bindings to f1546

  // f1548
  logic [0:0] f1548_wen;
  logic [31:0] f1548_wdata;
  logic [0:0] f1548_clk;
  logic [0:0] f1548_rst;
  logic [31:0] f1548_rdata;
  sr_buffer_32_1 f1548(.wen(f1548_wen), .wdata(f1548_wdata), .clk(f1548_clk), .rst(f1548_rst), .rdata(f1548_rdata));
  assign f1548_clk = clk;
  assign f1548_rst = rst;
  // Bindings to f1548

  // f1550
  logic [0:0] f1550_wen;
  logic [31:0] f1550_wdata;
  logic [0:0] f1550_clk;
  logic [0:0] f1550_rst;
  logic [31:0] f1550_rdata;
  sr_buffer_32_1 f1550(.wen(f1550_wen), .wdata(f1550_wdata), .clk(f1550_clk), .rst(f1550_rst), .rdata(f1550_rdata));
  assign f1550_clk = clk;
  assign f1550_rst = rst;
  // Bindings to f1550

  // f1552
  logic [0:0] f1552_wen;
  logic [31:0] f1552_wdata;
  logic [0:0] f1552_clk;
  logic [0:0] f1552_rst;
  logic [31:0] f1552_rdata;
  sr_buffer_32_1 f1552(.wen(f1552_wen), .wdata(f1552_wdata), .clk(f1552_clk), .rst(f1552_rst), .rdata(f1552_rdata));
  assign f1552_clk = clk;
  assign f1552_rst = rst;
  // Bindings to f1552

  // f1554
  logic [0:0] f1554_wen;
  logic [31:0] f1554_wdata;
  logic [0:0] f1554_clk;
  logic [0:0] f1554_rst;
  logic [31:0] f1554_rdata;
  sr_buffer_32_1 f1554(.wen(f1554_wen), .wdata(f1554_wdata), .clk(f1554_clk), .rst(f1554_rst), .rdata(f1554_rdata));
  assign f1554_clk = clk;
  assign f1554_rst = rst;
  // Bindings to f1554

  // f1556
  logic [0:0] f1556_wen;
  logic [31:0] f1556_wdata;
  logic [0:0] f1556_clk;
  logic [0:0] f1556_rst;
  logic [31:0] f1556_rdata;
  sr_buffer_32_1 f1556(.wen(f1556_wen), .wdata(f1556_wdata), .clk(f1556_clk), .rst(f1556_rst), .rdata(f1556_rdata));
  assign f1556_clk = clk;
  assign f1556_rst = rst;
  // Bindings to f1556

  // f1558
  logic [0:0] f1558_wen;
  logic [31:0] f1558_wdata;
  logic [0:0] f1558_clk;
  logic [0:0] f1558_rst;
  logic [31:0] f1558_rdata;
  sr_buffer_32_1 f1558(.wen(f1558_wen), .wdata(f1558_wdata), .clk(f1558_clk), .rst(f1558_rst), .rdata(f1558_rdata));
  assign f1558_clk = clk;
  assign f1558_rst = rst;
  // Bindings to f1558

  // f1560
  logic [0:0] f1560_wen;
  logic [31:0] f1560_wdata;
  logic [0:0] f1560_clk;
  logic [0:0] f1560_rst;
  logic [31:0] f1560_rdata;
  sr_buffer_32_1 f1560(.wen(f1560_wen), .wdata(f1560_wdata), .clk(f1560_clk), .rst(f1560_rst), .rdata(f1560_rdata));
  assign f1560_clk = clk;
  assign f1560_rst = rst;
  // Bindings to f1560

  // f1562
  logic [0:0] f1562_wen;
  logic [31:0] f1562_wdata;
  logic [0:0] f1562_clk;
  logic [0:0] f1562_rst;
  logic [31:0] f1562_rdata;
  sr_buffer_32_1 f1562(.wen(f1562_wen), .wdata(f1562_wdata), .clk(f1562_clk), .rst(f1562_rst), .rdata(f1562_rdata));
  assign f1562_clk = clk;
  assign f1562_rst = rst;
  // Bindings to f1562

  // f1564
  logic [0:0] f1564_wen;
  logic [31:0] f1564_wdata;
  logic [0:0] f1564_clk;
  logic [0:0] f1564_rst;
  logic [31:0] f1564_rdata;
  sr_buffer_32_1 f1564(.wen(f1564_wen), .wdata(f1564_wdata), .clk(f1564_clk), .rst(f1564_rst), .rdata(f1564_rdata));
  assign f1564_clk = clk;
  assign f1564_rst = rst;
  // Bindings to f1564

  // f1566
  logic [0:0] f1566_wen;
  logic [31:0] f1566_wdata;
  logic [0:0] f1566_clk;
  logic [0:0] f1566_rst;
  logic [31:0] f1566_rdata;
  sr_buffer_32_1 f1566(.wen(f1566_wen), .wdata(f1566_wdata), .clk(f1566_clk), .rst(f1566_rst), .rdata(f1566_rdata));
  assign f1566_clk = clk;
  assign f1566_rst = rst;
  // Bindings to f1566

  // f1568
  logic [0:0] f1568_wen;
  logic [31:0] f1568_wdata;
  logic [0:0] f1568_clk;
  logic [0:0] f1568_rst;
  logic [31:0] f1568_rdata;
  sr_buffer_32_1 f1568(.wen(f1568_wen), .wdata(f1568_wdata), .clk(f1568_clk), .rst(f1568_rst), .rdata(f1568_rdata));
  assign f1568_clk = clk;
  assign f1568_rst = rst;
  // Bindings to f1568

  // f1570
  logic [0:0] f1570_wen;
  logic [31:0] f1570_wdata;
  logic [0:0] f1570_clk;
  logic [0:0] f1570_rst;
  logic [31:0] f1570_rdata;
  sr_buffer_32_1 f1570(.wen(f1570_wen), .wdata(f1570_wdata), .clk(f1570_clk), .rst(f1570_rst), .rdata(f1570_rdata));
  assign f1570_clk = clk;
  assign f1570_rst = rst;
  // Bindings to f1570

  // f1572
  logic [0:0] f1572_wen;
  logic [31:0] f1572_wdata;
  logic [0:0] f1572_clk;
  logic [0:0] f1572_rst;
  logic [31:0] f1572_rdata;
  sr_buffer_32_1 f1572(.wen(f1572_wen), .wdata(f1572_wdata), .clk(f1572_clk), .rst(f1572_rst), .rdata(f1572_rdata));
  assign f1572_clk = clk;
  assign f1572_rst = rst;
  // Bindings to f1572

  // f1574
  logic [0:0] f1574_wen;
  logic [31:0] f1574_wdata;
  logic [0:0] f1574_clk;
  logic [0:0] f1574_rst;
  logic [31:0] f1574_rdata;
  sr_buffer_32_1 f1574(.wen(f1574_wen), .wdata(f1574_wdata), .clk(f1574_clk), .rst(f1574_rst), .rdata(f1574_rdata));
  assign f1574_clk = clk;
  assign f1574_rst = rst;
  // Bindings to f1574

  // f1576
  logic [0:0] f1576_wen;
  logic [31:0] f1576_wdata;
  logic [0:0] f1576_clk;
  logic [0:0] f1576_rst;
  logic [31:0] f1576_rdata;
  sr_buffer_32_1 f1576(.wen(f1576_wen), .wdata(f1576_wdata), .clk(f1576_clk), .rst(f1576_rst), .rdata(f1576_rdata));
  assign f1576_clk = clk;
  assign f1576_rst = rst;
  // Bindings to f1576

  // f1578
  logic [0:0] f1578_wen;
  logic [31:0] f1578_wdata;
  logic [0:0] f1578_clk;
  logic [0:0] f1578_rst;
  logic [31:0] f1578_rdata;
  sr_buffer_32_1 f1578(.wen(f1578_wen), .wdata(f1578_wdata), .clk(f1578_clk), .rst(f1578_rst), .rdata(f1578_rdata));
  assign f1578_clk = clk;
  assign f1578_rst = rst;
  // Bindings to f1578

  // f1580
  logic [0:0] f1580_wen;
  logic [31:0] f1580_wdata;
  logic [0:0] f1580_clk;
  logic [0:0] f1580_rst;
  logic [31:0] f1580_rdata;
  sr_buffer_32_1 f1580(.wen(f1580_wen), .wdata(f1580_wdata), .clk(f1580_clk), .rst(f1580_rst), .rdata(f1580_rdata));
  assign f1580_clk = clk;
  assign f1580_rst = rst;
  // Bindings to f1580

  // f1582
  logic [0:0] f1582_wen;
  logic [31:0] f1582_wdata;
  logic [0:0] f1582_clk;
  logic [0:0] f1582_rst;
  logic [31:0] f1582_rdata;
  sr_buffer_32_1 f1582(.wen(f1582_wen), .wdata(f1582_wdata), .clk(f1582_clk), .rst(f1582_rst), .rdata(f1582_rdata));
  assign f1582_clk = clk;
  assign f1582_rst = rst;
  // Bindings to f1582

  // f1584
  logic [0:0] f1584_wen;
  logic [31:0] f1584_wdata;
  logic [0:0] f1584_clk;
  logic [0:0] f1584_rst;
  logic [31:0] f1584_rdata;
  sr_buffer_32_1 f1584(.wen(f1584_wen), .wdata(f1584_wdata), .clk(f1584_clk), .rst(f1584_rst), .rdata(f1584_rdata));
  assign f1584_clk = clk;
  assign f1584_rst = rst;
  // Bindings to f1584

  // f1586
  logic [0:0] f1586_wen;
  logic [31:0] f1586_wdata;
  logic [0:0] f1586_clk;
  logic [0:0] f1586_rst;
  logic [31:0] f1586_rdata;
  sr_buffer_32_1 f1586(.wen(f1586_wen), .wdata(f1586_wdata), .clk(f1586_clk), .rst(f1586_rst), .rdata(f1586_rdata));
  assign f1586_clk = clk;
  assign f1586_rst = rst;
  // Bindings to f1586

  // f1588
  logic [0:0] f1588_wen;
  logic [31:0] f1588_wdata;
  logic [0:0] f1588_clk;
  logic [0:0] f1588_rst;
  logic [31:0] f1588_rdata;
  sr_buffer_32_1 f1588(.wen(f1588_wen), .wdata(f1588_wdata), .clk(f1588_clk), .rst(f1588_rst), .rdata(f1588_rdata));
  assign f1588_clk = clk;
  assign f1588_rst = rst;
  // Bindings to f1588

  // f1590
  logic [0:0] f1590_wen;
  logic [31:0] f1590_wdata;
  logic [0:0] f1590_clk;
  logic [0:0] f1590_rst;
  logic [31:0] f1590_rdata;
  sr_buffer_32_1 f1590(.wen(f1590_wen), .wdata(f1590_wdata), .clk(f1590_clk), .rst(f1590_rst), .rdata(f1590_rdata));
  assign f1590_clk = clk;
  assign f1590_rst = rst;
  // Bindings to f1590

  // f1592
  logic [0:0] f1592_wen;
  logic [31:0] f1592_wdata;
  logic [0:0] f1592_clk;
  logic [0:0] f1592_rst;
  logic [31:0] f1592_rdata;
  sr_buffer_32_1 f1592(.wen(f1592_wen), .wdata(f1592_wdata), .clk(f1592_clk), .rst(f1592_rst), .rdata(f1592_rdata));
  assign f1592_clk = clk;
  assign f1592_rst = rst;
  // Bindings to f1592

  // f1594
  logic [0:0] f1594_wen;
  logic [31:0] f1594_wdata;
  logic [0:0] f1594_clk;
  logic [0:0] f1594_rst;
  logic [31:0] f1594_rdata;
  sr_buffer_32_1 f1594(.wen(f1594_wen), .wdata(f1594_wdata), .clk(f1594_clk), .rst(f1594_rst), .rdata(f1594_rdata));
  assign f1594_clk = clk;
  assign f1594_rst = rst;
  // Bindings to f1594

  // f1596
  logic [0:0] f1596_wen;
  logic [31:0] f1596_wdata;
  logic [0:0] f1596_clk;
  logic [0:0] f1596_rst;
  logic [31:0] f1596_rdata;
  sr_buffer_32_1 f1596(.wen(f1596_wen), .wdata(f1596_wdata), .clk(f1596_clk), .rst(f1596_rst), .rdata(f1596_rdata));
  assign f1596_clk = clk;
  assign f1596_rst = rst;
  // Bindings to f1596

  // f1598
  logic [0:0] f1598_wen;
  logic [31:0] f1598_wdata;
  logic [0:0] f1598_clk;
  logic [0:0] f1598_rst;
  logic [31:0] f1598_rdata;
  sr_buffer_32_1 f1598(.wen(f1598_wen), .wdata(f1598_wdata), .clk(f1598_clk), .rst(f1598_rst), .rdata(f1598_rdata));
  assign f1598_clk = clk;
  assign f1598_rst = rst;
  // Bindings to f1598

  // f1600
  logic [0:0] f1600_wen;
  logic [31:0] f1600_wdata;
  logic [0:0] f1600_clk;
  logic [0:0] f1600_rst;
  logic [31:0] f1600_rdata;
  sr_buffer_32_1 f1600(.wen(f1600_wen), .wdata(f1600_wdata), .clk(f1600_clk), .rst(f1600_rst), .rdata(f1600_rdata));
  assign f1600_clk = clk;
  assign f1600_rst = rst;
  // Bindings to f1600

  // f1602
  logic [0:0] f1602_wen;
  logic [31:0] f1602_wdata;
  logic [0:0] f1602_clk;
  logic [0:0] f1602_rst;
  logic [31:0] f1602_rdata;
  sr_buffer_32_1 f1602(.wen(f1602_wen), .wdata(f1602_wdata), .clk(f1602_clk), .rst(f1602_rst), .rdata(f1602_rdata));
  assign f1602_clk = clk;
  assign f1602_rst = rst;
  // Bindings to f1602

  // f1604
  logic [0:0] f1604_wen;
  logic [31:0] f1604_wdata;
  logic [0:0] f1604_clk;
  logic [0:0] f1604_rst;
  logic [31:0] f1604_rdata;
  sr_buffer_32_1 f1604(.wen(f1604_wen), .wdata(f1604_wdata), .clk(f1604_clk), .rst(f1604_rst), .rdata(f1604_rdata));
  assign f1604_clk = clk;
  assign f1604_rst = rst;
  // Bindings to f1604

  // f1606
  logic [0:0] f1606_wen;
  logic [31:0] f1606_wdata;
  logic [0:0] f1606_clk;
  logic [0:0] f1606_rst;
  logic [31:0] f1606_rdata;
  sr_buffer_32_1 f1606(.wen(f1606_wen), .wdata(f1606_wdata), .clk(f1606_clk), .rst(f1606_rst), .rdata(f1606_rdata));
  assign f1606_clk = clk;
  assign f1606_rst = rst;
  // Bindings to f1606

  // f1608
  logic [0:0] f1608_wen;
  logic [31:0] f1608_wdata;
  logic [0:0] f1608_clk;
  logic [0:0] f1608_rst;
  logic [31:0] f1608_rdata;
  sr_buffer_32_1 f1608(.wen(f1608_wen), .wdata(f1608_wdata), .clk(f1608_clk), .rst(f1608_rst), .rdata(f1608_rdata));
  assign f1608_clk = clk;
  assign f1608_rst = rst;
  // Bindings to f1608

  // f1610
  logic [0:0] f1610_wen;
  logic [31:0] f1610_wdata;
  logic [0:0] f1610_clk;
  logic [0:0] f1610_rst;
  logic [31:0] f1610_rdata;
  sr_buffer_32_1 f1610(.wen(f1610_wen), .wdata(f1610_wdata), .clk(f1610_clk), .rst(f1610_rst), .rdata(f1610_rdata));
  assign f1610_clk = clk;
  assign f1610_rst = rst;
  // Bindings to f1610

  // f1612
  logic [0:0] f1612_wen;
  logic [31:0] f1612_wdata;
  logic [0:0] f1612_clk;
  logic [0:0] f1612_rst;
  logic [31:0] f1612_rdata;
  sr_buffer_32_1 f1612(.wen(f1612_wen), .wdata(f1612_wdata), .clk(f1612_clk), .rst(f1612_rst), .rdata(f1612_rdata));
  assign f1612_clk = clk;
  assign f1612_rst = rst;
  // Bindings to f1612

  // f1614
  logic [0:0] f1614_wen;
  logic [31:0] f1614_wdata;
  logic [0:0] f1614_clk;
  logic [0:0] f1614_rst;
  logic [31:0] f1614_rdata;
  sr_buffer_32_1 f1614(.wen(f1614_wen), .wdata(f1614_wdata), .clk(f1614_clk), .rst(f1614_rst), .rdata(f1614_rdata));
  assign f1614_clk = clk;
  assign f1614_rst = rst;
  // Bindings to f1614

  // f1616
  logic [0:0] f1616_wen;
  logic [31:0] f1616_wdata;
  logic [0:0] f1616_clk;
  logic [0:0] f1616_rst;
  logic [31:0] f1616_rdata;
  sr_buffer_32_1 f1616(.wen(f1616_wen), .wdata(f1616_wdata), .clk(f1616_clk), .rst(f1616_rst), .rdata(f1616_rdata));
  assign f1616_clk = clk;
  assign f1616_rst = rst;
  // Bindings to f1616

  // f1618
  logic [0:0] f1618_wen;
  logic [31:0] f1618_wdata;
  logic [0:0] f1618_clk;
  logic [0:0] f1618_rst;
  logic [31:0] f1618_rdata;
  sr_buffer_32_1 f1618(.wen(f1618_wen), .wdata(f1618_wdata), .clk(f1618_clk), .rst(f1618_rst), .rdata(f1618_rdata));
  assign f1618_clk = clk;
  assign f1618_rst = rst;
  // Bindings to f1618

  // f1620
  logic [0:0] f1620_wen;
  logic [31:0] f1620_wdata;
  logic [0:0] f1620_clk;
  logic [0:0] f1620_rst;
  logic [31:0] f1620_rdata;
  sr_buffer_32_1 f1620(.wen(f1620_wen), .wdata(f1620_wdata), .clk(f1620_clk), .rst(f1620_rst), .rdata(f1620_rdata));
  assign f1620_clk = clk;
  assign f1620_rst = rst;
  // Bindings to f1620

  // f1622
  logic [0:0] f1622_wen;
  logic [31:0] f1622_wdata;
  logic [0:0] f1622_clk;
  logic [0:0] f1622_rst;
  logic [31:0] f1622_rdata;
  sr_buffer_32_1 f1622(.wen(f1622_wen), .wdata(f1622_wdata), .clk(f1622_clk), .rst(f1622_rst), .rdata(f1622_rdata));
  assign f1622_clk = clk;
  assign f1622_rst = rst;
  // Bindings to f1622

  // f1624
  logic [0:0] f1624_wen;
  logic [31:0] f1624_wdata;
  logic [0:0] f1624_clk;
  logic [0:0] f1624_rst;
  logic [31:0] f1624_rdata;
  sr_buffer_32_1 f1624(.wen(f1624_wen), .wdata(f1624_wdata), .clk(f1624_clk), .rst(f1624_rst), .rdata(f1624_rdata));
  assign f1624_clk = clk;
  assign f1624_rst = rst;
  // Bindings to f1624

  // f1626
  logic [0:0] f1626_wen;
  logic [31:0] f1626_wdata;
  logic [0:0] f1626_clk;
  logic [0:0] f1626_rst;
  logic [31:0] f1626_rdata;
  sr_buffer_32_1 f1626(.wen(f1626_wen), .wdata(f1626_wdata), .clk(f1626_clk), .rst(f1626_rst), .rdata(f1626_rdata));
  assign f1626_clk = clk;
  assign f1626_rst = rst;
  // Bindings to f1626

  // f1628
  logic [0:0] f1628_wen;
  logic [31:0] f1628_wdata;
  logic [0:0] f1628_clk;
  logic [0:0] f1628_rst;
  logic [31:0] f1628_rdata;
  sr_buffer_32_1 f1628(.wen(f1628_wen), .wdata(f1628_wdata), .clk(f1628_clk), .rst(f1628_rst), .rdata(f1628_rdata));
  assign f1628_clk = clk;
  assign f1628_rst = rst;
  // Bindings to f1628

  // f1630
  logic [0:0] f1630_wen;
  logic [31:0] f1630_wdata;
  logic [0:0] f1630_clk;
  logic [0:0] f1630_rst;
  logic [31:0] f1630_rdata;
  sr_buffer_32_1 f1630(.wen(f1630_wen), .wdata(f1630_wdata), .clk(f1630_clk), .rst(f1630_rst), .rdata(f1630_rdata));
  assign f1630_clk = clk;
  assign f1630_rst = rst;
  // Bindings to f1630

  // f1632
  logic [0:0] f1632_wen;
  logic [31:0] f1632_wdata;
  logic [0:0] f1632_clk;
  logic [0:0] f1632_rst;
  logic [31:0] f1632_rdata;
  sr_buffer_32_1 f1632(.wen(f1632_wen), .wdata(f1632_wdata), .clk(f1632_clk), .rst(f1632_rst), .rdata(f1632_rdata));
  assign f1632_clk = clk;
  assign f1632_rst = rst;
  // Bindings to f1632

  // f1634
  logic [0:0] f1634_wen;
  logic [31:0] f1634_wdata;
  logic [0:0] f1634_clk;
  logic [0:0] f1634_rst;
  logic [31:0] f1634_rdata;
  sr_buffer_32_1 f1634(.wen(f1634_wen), .wdata(f1634_wdata), .clk(f1634_clk), .rst(f1634_rst), .rdata(f1634_rdata));
  assign f1634_clk = clk;
  assign f1634_rst = rst;
  // Bindings to f1634

  // f1636
  logic [0:0] f1636_wen;
  logic [31:0] f1636_wdata;
  logic [0:0] f1636_clk;
  logic [0:0] f1636_rst;
  logic [31:0] f1636_rdata;
  sr_buffer_32_1 f1636(.wen(f1636_wen), .wdata(f1636_wdata), .clk(f1636_clk), .rst(f1636_rst), .rdata(f1636_rdata));
  assign f1636_clk = clk;
  assign f1636_rst = rst;
  // Bindings to f1636

  // f1638
  logic [0:0] f1638_wen;
  logic [31:0] f1638_wdata;
  logic [0:0] f1638_clk;
  logic [0:0] f1638_rst;
  logic [31:0] f1638_rdata;
  sr_buffer_32_1 f1638(.wen(f1638_wen), .wdata(f1638_wdata), .clk(f1638_clk), .rst(f1638_rst), .rdata(f1638_rdata));
  assign f1638_clk = clk;
  assign f1638_rst = rst;
  // Bindings to f1638

  // f1640
  logic [0:0] f1640_wen;
  logic [31:0] f1640_wdata;
  logic [0:0] f1640_clk;
  logic [0:0] f1640_rst;
  logic [31:0] f1640_rdata;
  sr_buffer_32_1 f1640(.wen(f1640_wen), .wdata(f1640_wdata), .clk(f1640_clk), .rst(f1640_rst), .rdata(f1640_rdata));
  assign f1640_clk = clk;
  assign f1640_rst = rst;
  // Bindings to f1640

  // f1642
  logic [0:0] f1642_wen;
  logic [31:0] f1642_wdata;
  logic [0:0] f1642_clk;
  logic [0:0] f1642_rst;
  logic [31:0] f1642_rdata;
  sr_buffer_32_1 f1642(.wen(f1642_wen), .wdata(f1642_wdata), .clk(f1642_clk), .rst(f1642_rst), .rdata(f1642_rdata));
  assign f1642_clk = clk;
  assign f1642_rst = rst;
  // Bindings to f1642

  // f1644
  logic [0:0] f1644_wen;
  logic [31:0] f1644_wdata;
  logic [0:0] f1644_clk;
  logic [0:0] f1644_rst;
  logic [31:0] f1644_rdata;
  sr_buffer_32_1 f1644(.wen(f1644_wen), .wdata(f1644_wdata), .clk(f1644_clk), .rst(f1644_rst), .rdata(f1644_rdata));
  assign f1644_clk = clk;
  assign f1644_rst = rst;
  // Bindings to f1644

  // f1646
  logic [0:0] f1646_wen;
  logic [31:0] f1646_wdata;
  logic [0:0] f1646_clk;
  logic [0:0] f1646_rst;
  logic [31:0] f1646_rdata;
  sr_buffer_32_1 f1646(.wen(f1646_wen), .wdata(f1646_wdata), .clk(f1646_clk), .rst(f1646_rst), .rdata(f1646_rdata));
  assign f1646_clk = clk;
  assign f1646_rst = rst;
  // Bindings to f1646

  // f1648
  logic [0:0] f1648_wen;
  logic [31:0] f1648_wdata;
  logic [0:0] f1648_clk;
  logic [0:0] f1648_rst;
  logic [31:0] f1648_rdata;
  sr_buffer_32_1 f1648(.wen(f1648_wen), .wdata(f1648_wdata), .clk(f1648_clk), .rst(f1648_rst), .rdata(f1648_rdata));
  assign f1648_clk = clk;
  assign f1648_rst = rst;
  // Bindings to f1648

  // f1650
  logic [0:0] f1650_wen;
  logic [31:0] f1650_wdata;
  logic [0:0] f1650_clk;
  logic [0:0] f1650_rst;
  logic [31:0] f1650_rdata;
  sr_buffer_32_1 f1650(.wen(f1650_wen), .wdata(f1650_wdata), .clk(f1650_clk), .rst(f1650_rst), .rdata(f1650_rdata));
  assign f1650_clk = clk;
  assign f1650_rst = rst;
  // Bindings to f1650

  // f1652
  logic [0:0] f1652_wen;
  logic [31:0] f1652_wdata;
  logic [0:0] f1652_clk;
  logic [0:0] f1652_rst;
  logic [31:0] f1652_rdata;
  sr_buffer_32_1 f1652(.wen(f1652_wen), .wdata(f1652_wdata), .clk(f1652_clk), .rst(f1652_rst), .rdata(f1652_rdata));
  assign f1652_clk = clk;
  assign f1652_rst = rst;
  // Bindings to f1652

  // f1654
  logic [0:0] f1654_wen;
  logic [31:0] f1654_wdata;
  logic [0:0] f1654_clk;
  logic [0:0] f1654_rst;
  logic [31:0] f1654_rdata;
  sr_buffer_32_1 f1654(.wen(f1654_wen), .wdata(f1654_wdata), .clk(f1654_clk), .rst(f1654_rst), .rdata(f1654_rdata));
  assign f1654_clk = clk;
  assign f1654_rst = rst;
  // Bindings to f1654

  // f1656
  logic [0:0] f1656_wen;
  logic [31:0] f1656_wdata;
  logic [0:0] f1656_clk;
  logic [0:0] f1656_rst;
  logic [31:0] f1656_rdata;
  sr_buffer_32_1 f1656(.wen(f1656_wen), .wdata(f1656_wdata), .clk(f1656_clk), .rst(f1656_rst), .rdata(f1656_rdata));
  assign f1656_clk = clk;
  assign f1656_rst = rst;
  // Bindings to f1656

  // f1658
  logic [0:0] f1658_wen;
  logic [31:0] f1658_wdata;
  logic [0:0] f1658_clk;
  logic [0:0] f1658_rst;
  logic [31:0] f1658_rdata;
  sr_buffer_32_1 f1658(.wen(f1658_wen), .wdata(f1658_wdata), .clk(f1658_clk), .rst(f1658_rst), .rdata(f1658_rdata));
  assign f1658_clk = clk;
  assign f1658_rst = rst;
  // Bindings to f1658

  // f1660
  logic [0:0] f1660_wen;
  logic [31:0] f1660_wdata;
  logic [0:0] f1660_clk;
  logic [0:0] f1660_rst;
  logic [31:0] f1660_rdata;
  sr_buffer_32_1 f1660(.wen(f1660_wen), .wdata(f1660_wdata), .clk(f1660_clk), .rst(f1660_rst), .rdata(f1660_rdata));
  assign f1660_clk = clk;
  assign f1660_rst = rst;
  // Bindings to f1660

  // f1662
  logic [0:0] f1662_wen;
  logic [31:0] f1662_wdata;
  logic [0:0] f1662_clk;
  logic [0:0] f1662_rst;
  logic [31:0] f1662_rdata;
  sr_buffer_32_1 f1662(.wen(f1662_wen), .wdata(f1662_wdata), .clk(f1662_clk), .rst(f1662_rst), .rdata(f1662_rdata));
  assign f1662_clk = clk;
  assign f1662_rst = rst;
  // Bindings to f1662

  // f1664
  logic [0:0] f1664_wen;
  logic [31:0] f1664_wdata;
  logic [0:0] f1664_clk;
  logic [0:0] f1664_rst;
  logic [31:0] f1664_rdata;
  sr_buffer_32_1 f1664(.wen(f1664_wen), .wdata(f1664_wdata), .clk(f1664_clk), .rst(f1664_rst), .rdata(f1664_rdata));
  assign f1664_clk = clk;
  assign f1664_rst = rst;
  // Bindings to f1664

  // f1666
  logic [0:0] f1666_wen;
  logic [31:0] f1666_wdata;
  logic [0:0] f1666_clk;
  logic [0:0] f1666_rst;
  logic [31:0] f1666_rdata;
  sr_buffer_32_1 f1666(.wen(f1666_wen), .wdata(f1666_wdata), .clk(f1666_clk), .rst(f1666_rst), .rdata(f1666_rdata));
  assign f1666_clk = clk;
  assign f1666_rst = rst;
  // Bindings to f1666

  // f1668
  logic [0:0] f1668_wen;
  logic [31:0] f1668_wdata;
  logic [0:0] f1668_clk;
  logic [0:0] f1668_rst;
  logic [31:0] f1668_rdata;
  sr_buffer_32_1 f1668(.wen(f1668_wen), .wdata(f1668_wdata), .clk(f1668_clk), .rst(f1668_rst), .rdata(f1668_rdata));
  assign f1668_clk = clk;
  assign f1668_rst = rst;
  // Bindings to f1668

  // f1670
  logic [0:0] f1670_wen;
  logic [31:0] f1670_wdata;
  logic [0:0] f1670_clk;
  logic [0:0] f1670_rst;
  logic [31:0] f1670_rdata;
  sr_buffer_32_1 f1670(.wen(f1670_wen), .wdata(f1670_wdata), .clk(f1670_clk), .rst(f1670_rst), .rdata(f1670_rdata));
  assign f1670_clk = clk;
  assign f1670_rst = rst;
  // Bindings to f1670

  // f1672
  logic [0:0] f1672_wen;
  logic [31:0] f1672_wdata;
  logic [0:0] f1672_clk;
  logic [0:0] f1672_rst;
  logic [31:0] f1672_rdata;
  sr_buffer_32_1 f1672(.wen(f1672_wen), .wdata(f1672_wdata), .clk(f1672_clk), .rst(f1672_rst), .rdata(f1672_rdata));
  assign f1672_clk = clk;
  assign f1672_rst = rst;
  // Bindings to f1672

  // f1674
  logic [0:0] f1674_wen;
  logic [31:0] f1674_wdata;
  logic [0:0] f1674_clk;
  logic [0:0] f1674_rst;
  logic [31:0] f1674_rdata;
  sr_buffer_32_1 f1674(.wen(f1674_wen), .wdata(f1674_wdata), .clk(f1674_clk), .rst(f1674_rst), .rdata(f1674_rdata));
  assign f1674_clk = clk;
  assign f1674_rst = rst;
  // Bindings to f1674

  // f1676
  logic [0:0] f1676_wen;
  logic [31:0] f1676_wdata;
  logic [0:0] f1676_clk;
  logic [0:0] f1676_rst;
  logic [31:0] f1676_rdata;
  sr_buffer_32_1 f1676(.wen(f1676_wen), .wdata(f1676_wdata), .clk(f1676_clk), .rst(f1676_rst), .rdata(f1676_rdata));
  assign f1676_clk = clk;
  assign f1676_rst = rst;
  // Bindings to f1676

  // f1678
  logic [0:0] f1678_wen;
  logic [31:0] f1678_wdata;
  logic [0:0] f1678_clk;
  logic [0:0] f1678_rst;
  logic [31:0] f1678_rdata;
  sr_buffer_32_1 f1678(.wen(f1678_wen), .wdata(f1678_wdata), .clk(f1678_clk), .rst(f1678_rst), .rdata(f1678_rdata));
  assign f1678_clk = clk;
  assign f1678_rst = rst;
  // Bindings to f1678

  // f1680
  logic [0:0] f1680_wen;
  logic [31:0] f1680_wdata;
  logic [0:0] f1680_clk;
  logic [0:0] f1680_rst;
  logic [31:0] f1680_rdata;
  sr_buffer_32_1 f1680(.wen(f1680_wen), .wdata(f1680_wdata), .clk(f1680_clk), .rst(f1680_rst), .rdata(f1680_rdata));
  assign f1680_clk = clk;
  assign f1680_rst = rst;
  // Bindings to f1680

  // f1682
  logic [0:0] f1682_wen;
  logic [31:0] f1682_wdata;
  logic [0:0] f1682_clk;
  logic [0:0] f1682_rst;
  logic [31:0] f1682_rdata;
  sr_buffer_32_1 f1682(.wen(f1682_wen), .wdata(f1682_wdata), .clk(f1682_clk), .rst(f1682_rst), .rdata(f1682_rdata));
  assign f1682_clk = clk;
  assign f1682_rst = rst;
  // Bindings to f1682

  // f1684
  logic [0:0] f1684_wen;
  logic [31:0] f1684_wdata;
  logic [0:0] f1684_clk;
  logic [0:0] f1684_rst;
  logic [31:0] f1684_rdata;
  sr_buffer_32_1 f1684(.wen(f1684_wen), .wdata(f1684_wdata), .clk(f1684_clk), .rst(f1684_rst), .rdata(f1684_rdata));
  assign f1684_clk = clk;
  assign f1684_rst = rst;
  // Bindings to f1684

  // f1686
  logic [0:0] f1686_wen;
  logic [31:0] f1686_wdata;
  logic [0:0] f1686_clk;
  logic [0:0] f1686_rst;
  logic [31:0] f1686_rdata;
  sr_buffer_32_1 f1686(.wen(f1686_wen), .wdata(f1686_wdata), .clk(f1686_clk), .rst(f1686_rst), .rdata(f1686_rdata));
  assign f1686_clk = clk;
  assign f1686_rst = rst;
  // Bindings to f1686

  // f1688
  logic [0:0] f1688_wen;
  logic [31:0] f1688_wdata;
  logic [0:0] f1688_clk;
  logic [0:0] f1688_rst;
  logic [31:0] f1688_rdata;
  sr_buffer_32_1 f1688(.wen(f1688_wen), .wdata(f1688_wdata), .clk(f1688_clk), .rst(f1688_rst), .rdata(f1688_rdata));
  assign f1688_clk = clk;
  assign f1688_rst = rst;
  // Bindings to f1688

  // f1690
  logic [0:0] f1690_wen;
  logic [31:0] f1690_wdata;
  logic [0:0] f1690_clk;
  logic [0:0] f1690_rst;
  logic [31:0] f1690_rdata;
  sr_buffer_32_1 f1690(.wen(f1690_wen), .wdata(f1690_wdata), .clk(f1690_clk), .rst(f1690_rst), .rdata(f1690_rdata));
  assign f1690_clk = clk;
  assign f1690_rst = rst;
  // Bindings to f1690

  // f1692
  logic [0:0] f1692_wen;
  logic [31:0] f1692_wdata;
  logic [0:0] f1692_clk;
  logic [0:0] f1692_rst;
  logic [31:0] f1692_rdata;
  sr_buffer_32_1 f1692(.wen(f1692_wen), .wdata(f1692_wdata), .clk(f1692_clk), .rst(f1692_rst), .rdata(f1692_rdata));
  assign f1692_clk = clk;
  assign f1692_rst = rst;
  // Bindings to f1692

  // f1694
  logic [0:0] f1694_wen;
  logic [31:0] f1694_wdata;
  logic [0:0] f1694_clk;
  logic [0:0] f1694_rst;
  logic [31:0] f1694_rdata;
  sr_buffer_32_1 f1694(.wen(f1694_wen), .wdata(f1694_wdata), .clk(f1694_clk), .rst(f1694_rst), .rdata(f1694_rdata));
  assign f1694_clk = clk;
  assign f1694_rst = rst;
  // Bindings to f1694

  // f1696
  logic [0:0] f1696_wen;
  logic [31:0] f1696_wdata;
  logic [0:0] f1696_clk;
  logic [0:0] f1696_rst;
  logic [31:0] f1696_rdata;
  sr_buffer_32_1 f1696(.wen(f1696_wen), .wdata(f1696_wdata), .clk(f1696_clk), .rst(f1696_rst), .rdata(f1696_rdata));
  assign f1696_clk = clk;
  assign f1696_rst = rst;
  // Bindings to f1696

  // f1698
  logic [0:0] f1698_wen;
  logic [31:0] f1698_wdata;
  logic [0:0] f1698_clk;
  logic [0:0] f1698_rst;
  logic [31:0] f1698_rdata;
  sr_buffer_32_1 f1698(.wen(f1698_wen), .wdata(f1698_wdata), .clk(f1698_clk), .rst(f1698_rst), .rdata(f1698_rdata));
  assign f1698_clk = clk;
  assign f1698_rst = rst;
  // Bindings to f1698

  // f1700
  logic [0:0] f1700_wen;
  logic [31:0] f1700_wdata;
  logic [0:0] f1700_clk;
  logic [0:0] f1700_rst;
  logic [31:0] f1700_rdata;
  sr_buffer_32_1 f1700(.wen(f1700_wen), .wdata(f1700_wdata), .clk(f1700_clk), .rst(f1700_rst), .rdata(f1700_rdata));
  assign f1700_clk = clk;
  assign f1700_rst = rst;
  // Bindings to f1700

  // f1702
  logic [0:0] f1702_wen;
  logic [31:0] f1702_wdata;
  logic [0:0] f1702_clk;
  logic [0:0] f1702_rst;
  logic [31:0] f1702_rdata;
  sr_buffer_32_1 f1702(.wen(f1702_wen), .wdata(f1702_wdata), .clk(f1702_clk), .rst(f1702_rst), .rdata(f1702_rdata));
  assign f1702_clk = clk;
  assign f1702_rst = rst;
  // Bindings to f1702

  // f1704
  logic [0:0] f1704_wen;
  logic [31:0] f1704_wdata;
  logic [0:0] f1704_clk;
  logic [0:0] f1704_rst;
  logic [31:0] f1704_rdata;
  sr_buffer_32_1 f1704(.wen(f1704_wen), .wdata(f1704_wdata), .clk(f1704_clk), .rst(f1704_rst), .rdata(f1704_rdata));
  assign f1704_clk = clk;
  assign f1704_rst = rst;
  // Bindings to f1704

  // f1706
  logic [0:0] f1706_wen;
  logic [31:0] f1706_wdata;
  logic [0:0] f1706_clk;
  logic [0:0] f1706_rst;
  logic [31:0] f1706_rdata;
  sr_buffer_32_1 f1706(.wen(f1706_wen), .wdata(f1706_wdata), .clk(f1706_clk), .rst(f1706_rst), .rdata(f1706_rdata));
  assign f1706_clk = clk;
  assign f1706_rst = rst;
  // Bindings to f1706

  // f1708
  logic [0:0] f1708_wen;
  logic [31:0] f1708_wdata;
  logic [0:0] f1708_clk;
  logic [0:0] f1708_rst;
  logic [31:0] f1708_rdata;
  sr_buffer_32_1 f1708(.wen(f1708_wen), .wdata(f1708_wdata), .clk(f1708_clk), .rst(f1708_rst), .rdata(f1708_rdata));
  assign f1708_clk = clk;
  assign f1708_rst = rst;
  // Bindings to f1708

  // f1710
  logic [0:0] f1710_wen;
  logic [31:0] f1710_wdata;
  logic [0:0] f1710_clk;
  logic [0:0] f1710_rst;
  logic [31:0] f1710_rdata;
  sr_buffer_32_1 f1710(.wen(f1710_wen), .wdata(f1710_wdata), .clk(f1710_clk), .rst(f1710_rst), .rdata(f1710_rdata));
  assign f1710_clk = clk;
  assign f1710_rst = rst;
  // Bindings to f1710

  // f1712
  logic [0:0] f1712_wen;
  logic [31:0] f1712_wdata;
  logic [0:0] f1712_clk;
  logic [0:0] f1712_rst;
  logic [31:0] f1712_rdata;
  sr_buffer_32_1 f1712(.wen(f1712_wen), .wdata(f1712_wdata), .clk(f1712_clk), .rst(f1712_rst), .rdata(f1712_rdata));
  assign f1712_clk = clk;
  assign f1712_rst = rst;
  // Bindings to f1712

  // f1714
  logic [0:0] f1714_wen;
  logic [31:0] f1714_wdata;
  logic [0:0] f1714_clk;
  logic [0:0] f1714_rst;
  logic [31:0] f1714_rdata;
  sr_buffer_32_1 f1714(.wen(f1714_wen), .wdata(f1714_wdata), .clk(f1714_clk), .rst(f1714_rst), .rdata(f1714_rdata));
  assign f1714_clk = clk;
  assign f1714_rst = rst;
  // Bindings to f1714

  // f1770
  logic [0:0] f1770_wen;
  logic [31:0] f1770_wdata;
  logic [0:0] f1770_clk;
  logic [0:0] f1770_rst;
  logic [31:0] f1770_rdata;
  sr_buffer_32_1 f1770(.wen(f1770_wen), .wdata(f1770_wdata), .clk(f1770_clk), .rst(f1770_rst), .rdata(f1770_rdata));
  assign f1770_clk = clk;
  assign f1770_rst = rst;
  // Bindings to f1770

  // f1772
  logic [0:0] f1772_wen;
  logic [31:0] f1772_wdata;
  logic [0:0] f1772_clk;
  logic [0:0] f1772_rst;
  logic [31:0] f1772_rdata;
  sr_buffer_32_1 f1772(.wen(f1772_wen), .wdata(f1772_wdata), .clk(f1772_clk), .rst(f1772_rst), .rdata(f1772_rdata));
  assign f1772_clk = clk;
  assign f1772_rst = rst;
  // Bindings to f1772

  // f1718
  logic [0:0] f1718_wen;
  logic [31:0] f1718_wdata;
  logic [0:0] f1718_clk;
  logic [0:0] f1718_rst;
  logic [31:0] f1718_rdata;
  sr_buffer_32_1 f1718(.wen(f1718_wen), .wdata(f1718_wdata), .clk(f1718_clk), .rst(f1718_rst), .rdata(f1718_rdata));
  assign f1718_clk = clk;
  assign f1718_rst = rst;
  // Bindings to f1718

  // f1720
  logic [0:0] f1720_wen;
  logic [31:0] f1720_wdata;
  logic [0:0] f1720_clk;
  logic [0:0] f1720_rst;
  logic [31:0] f1720_rdata;
  sr_buffer_32_1 f1720(.wen(f1720_wen), .wdata(f1720_wdata), .clk(f1720_clk), .rst(f1720_rst), .rdata(f1720_rdata));
  assign f1720_clk = clk;
  assign f1720_rst = rst;
  // Bindings to f1720

  // f1716
  logic [0:0] f1716_wen;
  logic [31:0] f1716_wdata;
  logic [0:0] f1716_clk;
  logic [0:0] f1716_rst;
  logic [31:0] f1716_rdata;
  sr_buffer_32_1 f1716(.wen(f1716_wen), .wdata(f1716_wdata), .clk(f1716_clk), .rst(f1716_rst), .rdata(f1716_rdata));
  assign f1716_clk = clk;
  assign f1716_rst = rst;
  // Bindings to f1716

  // f1722
  logic [0:0] f1722_wen;
  logic [31:0] f1722_wdata;
  logic [0:0] f1722_clk;
  logic [0:0] f1722_rst;
  logic [31:0] f1722_rdata;
  sr_buffer_32_1 f1722(.wen(f1722_wen), .wdata(f1722_wdata), .clk(f1722_clk), .rst(f1722_rst), .rdata(f1722_rdata));
  assign f1722_clk = clk;
  assign f1722_rst = rst;
  // Bindings to f1722

  // f1730
  logic [0:0] f1730_wen;
  logic [31:0] f1730_wdata;
  logic [0:0] f1730_clk;
  logic [0:0] f1730_rst;
  logic [31:0] f1730_rdata;
  sr_buffer_32_1 f1730(.wen(f1730_wen), .wdata(f1730_wdata), .clk(f1730_clk), .rst(f1730_rst), .rdata(f1730_rdata));
  assign f1730_clk = clk;
  assign f1730_rst = rst;
  // Bindings to f1730

  // f1732
  logic [0:0] f1732_wen;
  logic [31:0] f1732_wdata;
  logic [0:0] f1732_clk;
  logic [0:0] f1732_rst;
  logic [31:0] f1732_rdata;
  sr_buffer_32_1 f1732(.wen(f1732_wen), .wdata(f1732_wdata), .clk(f1732_clk), .rst(f1732_rst), .rdata(f1732_rdata));
  assign f1732_clk = clk;
  assign f1732_rst = rst;
  // Bindings to f1732

  // f1728
  logic [0:0] f1728_wen;
  logic [31:0] f1728_wdata;
  logic [0:0] f1728_clk;
  logic [0:0] f1728_rst;
  logic [31:0] f1728_rdata;
  sr_buffer_32_1 f1728(.wen(f1728_wen), .wdata(f1728_wdata), .clk(f1728_clk), .rst(f1728_rst), .rdata(f1728_rdata));
  assign f1728_clk = clk;
  assign f1728_rst = rst;
  // Bindings to f1728

  // f1740
  logic [0:0] f1740_wen;
  logic [31:0] f1740_wdata;
  logic [0:0] f1740_clk;
  logic [0:0] f1740_rst;
  logic [31:0] f1740_rdata;
  sr_buffer_32_1 f1740(.wen(f1740_wen), .wdata(f1740_wdata), .clk(f1740_clk), .rst(f1740_rst), .rdata(f1740_rdata));
  assign f1740_clk = clk;
  assign f1740_rst = rst;
  // Bindings to f1740

  // f1734
  logic [0:0] f1734_wen;
  logic [31:0] f1734_wdata;
  logic [0:0] f1734_clk;
  logic [0:0] f1734_rst;
  logic [31:0] f1734_rdata;
  sr_buffer_32_1 f1734(.wen(f1734_wen), .wdata(f1734_wdata), .clk(f1734_clk), .rst(f1734_rst), .rdata(f1734_rdata));
  assign f1734_clk = clk;
  assign f1734_rst = rst;
  // Bindings to f1734

  // f1736
  logic [0:0] f1736_wen;
  logic [31:0] f1736_wdata;
  logic [0:0] f1736_clk;
  logic [0:0] f1736_rst;
  logic [31:0] f1736_rdata;
  sr_buffer_32_1 f1736(.wen(f1736_wen), .wdata(f1736_wdata), .clk(f1736_clk), .rst(f1736_rst), .rdata(f1736_rdata));
  assign f1736_clk = clk;
  assign f1736_rst = rst;
  // Bindings to f1736

  // f1750
  logic [0:0] f1750_wen;
  logic [31:0] f1750_wdata;
  logic [0:0] f1750_clk;
  logic [0:0] f1750_rst;
  logic [31:0] f1750_rdata;
  sr_buffer_32_1 f1750(.wen(f1750_wen), .wdata(f1750_wdata), .clk(f1750_clk), .rst(f1750_rst), .rdata(f1750_rdata));
  assign f1750_clk = clk;
  assign f1750_rst = rst;
  // Bindings to f1750

  // f1738
  logic [0:0] f1738_wen;
  logic [31:0] f1738_wdata;
  logic [0:0] f1738_clk;
  logic [0:0] f1738_rst;
  logic [31:0] f1738_rdata;
  sr_buffer_32_1 f1738(.wen(f1738_wen), .wdata(f1738_wdata), .clk(f1738_clk), .rst(f1738_rst), .rdata(f1738_rdata));
  assign f1738_clk = clk;
  assign f1738_rst = rst;
  // Bindings to f1738

  // f1742
  logic [0:0] f1742_wen;
  logic [31:0] f1742_wdata;
  logic [0:0] f1742_clk;
  logic [0:0] f1742_rst;
  logic [31:0] f1742_rdata;
  sr_buffer_32_1 f1742(.wen(f1742_wen), .wdata(f1742_wdata), .clk(f1742_clk), .rst(f1742_rst), .rdata(f1742_rdata));
  assign f1742_clk = clk;
  assign f1742_rst = rst;
  // Bindings to f1742

  // f1744
  logic [0:0] f1744_wen;
  logic [31:0] f1744_wdata;
  logic [0:0] f1744_clk;
  logic [0:0] f1744_rst;
  logic [31:0] f1744_rdata;
  sr_buffer_32_1 f1744(.wen(f1744_wen), .wdata(f1744_wdata), .clk(f1744_clk), .rst(f1744_rst), .rdata(f1744_rdata));
  assign f1744_clk = clk;
  assign f1744_rst = rst;
  // Bindings to f1744

  // f1726
  logic [0:0] f1726_wen;
  logic [31:0] f1726_wdata;
  logic [0:0] f1726_clk;
  logic [0:0] f1726_rst;
  logic [31:0] f1726_rdata;
  sr_buffer_32_1 f1726(.wen(f1726_wen), .wdata(f1726_wdata), .clk(f1726_clk), .rst(f1726_rst), .rdata(f1726_rdata));
  assign f1726_clk = clk;
  assign f1726_rst = rst;
  // Bindings to f1726

  // f1746
  logic [0:0] f1746_wen;
  logic [31:0] f1746_wdata;
  logic [0:0] f1746_clk;
  logic [0:0] f1746_rst;
  logic [31:0] f1746_rdata;
  sr_buffer_32_1 f1746(.wen(f1746_wen), .wdata(f1746_wdata), .clk(f1746_clk), .rst(f1746_rst), .rdata(f1746_rdata));
  assign f1746_clk = clk;
  assign f1746_rst = rst;
  // Bindings to f1746

  // f1766
  logic [0:0] f1766_wen;
  logic [31:0] f1766_wdata;
  logic [0:0] f1766_clk;
  logic [0:0] f1766_rst;
  logic [31:0] f1766_rdata;
  sr_buffer_32_1 f1766(.wen(f1766_wen), .wdata(f1766_wdata), .clk(f1766_clk), .rst(f1766_rst), .rdata(f1766_rdata));
  assign f1766_clk = clk;
  assign f1766_rst = rst;
  // Bindings to f1766

  // f1748
  logic [0:0] f1748_wen;
  logic [31:0] f1748_wdata;
  logic [0:0] f1748_clk;
  logic [0:0] f1748_rst;
  logic [31:0] f1748_rdata;
  sr_buffer_32_1 f1748(.wen(f1748_wen), .wdata(f1748_wdata), .clk(f1748_clk), .rst(f1748_rst), .rdata(f1748_rdata));
  assign f1748_clk = clk;
  assign f1748_rst = rst;
  // Bindings to f1748

  // f1764
  logic [0:0] f1764_wen;
  logic [31:0] f1764_wdata;
  logic [0:0] f1764_clk;
  logic [0:0] f1764_rst;
  logic [31:0] f1764_rdata;
  sr_buffer_32_1 f1764(.wen(f1764_wen), .wdata(f1764_wdata), .clk(f1764_clk), .rst(f1764_rst), .rdata(f1764_rdata));
  assign f1764_clk = clk;
  assign f1764_rst = rst;
  // Bindings to f1764

  // f1724
  logic [0:0] f1724_wen;
  logic [31:0] f1724_wdata;
  logic [0:0] f1724_clk;
  logic [0:0] f1724_rst;
  logic [31:0] f1724_rdata;
  sr_buffer_32_1 f1724(.wen(f1724_wen), .wdata(f1724_wdata), .clk(f1724_clk), .rst(f1724_rst), .rdata(f1724_rdata));
  assign f1724_clk = clk;
  assign f1724_rst = rst;
  // Bindings to f1724

  // f1762
  logic [0:0] f1762_wen;
  logic [31:0] f1762_wdata;
  logic [0:0] f1762_clk;
  logic [0:0] f1762_rst;
  logic [31:0] f1762_rdata;
  sr_buffer_32_1 f1762(.wen(f1762_wen), .wdata(f1762_wdata), .clk(f1762_clk), .rst(f1762_rst), .rdata(f1762_rdata));
  assign f1762_clk = clk;
  assign f1762_rst = rst;
  // Bindings to f1762

  // f1774
  logic [0:0] f1774_wen;
  logic [31:0] f1774_wdata;
  logic [0:0] f1774_clk;
  logic [0:0] f1774_rst;
  logic [31:0] f1774_rdata;
  sr_buffer_32_1 f1774(.wen(f1774_wen), .wdata(f1774_wdata), .clk(f1774_clk), .rst(f1774_rst), .rdata(f1774_rdata));
  assign f1774_clk = clk;
  assign f1774_rst = rst;
  // Bindings to f1774

  // f1756
  logic [0:0] f1756_wen;
  logic [31:0] f1756_wdata;
  logic [0:0] f1756_clk;
  logic [0:0] f1756_rst;
  logic [31:0] f1756_rdata;
  sr_buffer_32_1 f1756(.wen(f1756_wen), .wdata(f1756_wdata), .clk(f1756_clk), .rst(f1756_rst), .rdata(f1756_rdata));
  assign f1756_clk = clk;
  assign f1756_rst = rst;
  // Bindings to f1756

  // f1754
  logic [0:0] f1754_wen;
  logic [31:0] f1754_wdata;
  logic [0:0] f1754_clk;
  logic [0:0] f1754_rst;
  logic [31:0] f1754_rdata;
  sr_buffer_32_1 f1754(.wen(f1754_wen), .wdata(f1754_wdata), .clk(f1754_clk), .rst(f1754_rst), .rdata(f1754_rdata));
  assign f1754_clk = clk;
  assign f1754_rst = rst;
  // Bindings to f1754

  // f1760
  logic [0:0] f1760_wen;
  logic [31:0] f1760_wdata;
  logic [0:0] f1760_clk;
  logic [0:0] f1760_rst;
  logic [31:0] f1760_rdata;
  sr_buffer_32_1 f1760(.wen(f1760_wen), .wdata(f1760_wdata), .clk(f1760_clk), .rst(f1760_rst), .rdata(f1760_rdata));
  assign f1760_clk = clk;
  assign f1760_rst = rst;
  // Bindings to f1760

  // f1752
  logic [0:0] f1752_wen;
  logic [31:0] f1752_wdata;
  logic [0:0] f1752_clk;
  logic [0:0] f1752_rst;
  logic [31:0] f1752_rdata;
  sr_buffer_32_1 f1752(.wen(f1752_wen), .wdata(f1752_wdata), .clk(f1752_clk), .rst(f1752_rst), .rdata(f1752_rdata));
  assign f1752_clk = clk;
  assign f1752_rst = rst;
  // Bindings to f1752

  // f1768
  logic [0:0] f1768_wen;
  logic [31:0] f1768_wdata;
  logic [0:0] f1768_clk;
  logic [0:0] f1768_rst;
  logic [31:0] f1768_rdata;
  sr_buffer_32_1 f1768(.wen(f1768_wen), .wdata(f1768_wdata), .clk(f1768_clk), .rst(f1768_rst), .rdata(f1768_rdata));
  assign f1768_clk = clk;
  assign f1768_rst = rst;
  // Bindings to f1768

  // f1758
  logic [0:0] f1758_wen;
  logic [31:0] f1758_wdata;
  logic [0:0] f1758_clk;
  logic [0:0] f1758_rst;
  logic [31:0] f1758_rdata;
  sr_buffer_32_1 f1758(.wen(f1758_wen), .wdata(f1758_wdata), .clk(f1758_clk), .rst(f1758_rst), .rdata(f1758_rdata));
  assign f1758_clk = clk;
  assign f1758_rst = rst;
  // Bindings to f1758

  // f1776
  logic [0:0] f1776_wen;
  logic [31:0] f1776_wdata;
  logic [0:0] f1776_clk;
  logic [0:0] f1776_rst;
  logic [31:0] f1776_rdata;
  sr_buffer_32_1 f1776(.wen(f1776_wen), .wdata(f1776_wdata), .clk(f1776_clk), .rst(f1776_rst), .rdata(f1776_rdata));
  assign f1776_clk = clk;
  assign f1776_rst = rst;
  // Bindings to f1776

  // f1778
  logic [0:0] f1778_wen;
  logic [31:0] f1778_wdata;
  logic [0:0] f1778_clk;
  logic [0:0] f1778_rst;
  logic [31:0] f1778_rdata;
  sr_buffer_32_1 f1778(.wen(f1778_wen), .wdata(f1778_wdata), .clk(f1778_clk), .rst(f1778_rst), .rdata(f1778_rdata));
  assign f1778_clk = clk;
  assign f1778_rst = rst;
  // Bindings to f1778

  // f1780
  logic [0:0] f1780_wen;
  logic [31:0] f1780_wdata;
  logic [0:0] f1780_clk;
  logic [0:0] f1780_rst;
  logic [31:0] f1780_rdata;
  sr_buffer_32_1 f1780(.wen(f1780_wen), .wdata(f1780_wdata), .clk(f1780_clk), .rst(f1780_rst), .rdata(f1780_rdata));
  assign f1780_clk = clk;
  assign f1780_rst = rst;
  // Bindings to f1780

  // f1782
  logic [0:0] f1782_wen;
  logic [31:0] f1782_wdata;
  logic [0:0] f1782_clk;
  logic [0:0] f1782_rst;
  logic [31:0] f1782_rdata;
  sr_buffer_32_1 f1782(.wen(f1782_wen), .wdata(f1782_wdata), .clk(f1782_clk), .rst(f1782_rst), .rdata(f1782_rdata));
  assign f1782_clk = clk;
  assign f1782_rst = rst;
  // Bindings to f1782

  // f1784
  logic [0:0] f1784_wen;
  logic [31:0] f1784_wdata;
  logic [0:0] f1784_clk;
  logic [0:0] f1784_rst;
  logic [31:0] f1784_rdata;
  sr_buffer_32_1 f1784(.wen(f1784_wen), .wdata(f1784_wdata), .clk(f1784_clk), .rst(f1784_rst), .rdata(f1784_rdata));
  assign f1784_clk = clk;
  assign f1784_rst = rst;
  // Bindings to f1784

  // f1786
  logic [0:0] f1786_wen;
  logic [31:0] f1786_wdata;
  logic [0:0] f1786_clk;
  logic [0:0] f1786_rst;
  logic [31:0] f1786_rdata;
  sr_buffer_32_1 f1786(.wen(f1786_wen), .wdata(f1786_wdata), .clk(f1786_clk), .rst(f1786_rst), .rdata(f1786_rdata));
  assign f1786_clk = clk;
  assign f1786_rst = rst;
  // Bindings to f1786

  // f1788
  logic [0:0] f1788_wen;
  logic [31:0] f1788_wdata;
  logic [0:0] f1788_clk;
  logic [0:0] f1788_rst;
  logic [31:0] f1788_rdata;
  sr_buffer_32_1 f1788(.wen(f1788_wen), .wdata(f1788_wdata), .clk(f1788_clk), .rst(f1788_rst), .rdata(f1788_rdata));
  assign f1788_clk = clk;
  assign f1788_rst = rst;
  // Bindings to f1788

  // f1790
  logic [0:0] f1790_wen;
  logic [31:0] f1790_wdata;
  logic [0:0] f1790_clk;
  logic [0:0] f1790_rst;
  logic [31:0] f1790_rdata;
  sr_buffer_32_1 f1790(.wen(f1790_wen), .wdata(f1790_wdata), .clk(f1790_clk), .rst(f1790_rst), .rdata(f1790_rdata));
  assign f1790_clk = clk;
  assign f1790_rst = rst;
  // Bindings to f1790

  // f1792
  logic [0:0] f1792_wen;
  logic [31:0] f1792_wdata;
  logic [0:0] f1792_clk;
  logic [0:0] f1792_rst;
  logic [31:0] f1792_rdata;
  sr_buffer_32_1 f1792(.wen(f1792_wen), .wdata(f1792_wdata), .clk(f1792_clk), .rst(f1792_rst), .rdata(f1792_rdata));
  assign f1792_clk = clk;
  assign f1792_rst = rst;
  // Bindings to f1792

  // f1794
  logic [0:0] f1794_wen;
  logic [31:0] f1794_wdata;
  logic [0:0] f1794_clk;
  logic [0:0] f1794_rst;
  logic [31:0] f1794_rdata;
  sr_buffer_32_1 f1794(.wen(f1794_wen), .wdata(f1794_wdata), .clk(f1794_clk), .rst(f1794_rst), .rdata(f1794_rdata));
  assign f1794_clk = clk;
  assign f1794_rst = rst;
  // Bindings to f1794

  // f1796
  logic [0:0] f1796_wen;
  logic [31:0] f1796_wdata;
  logic [0:0] f1796_clk;
  logic [0:0] f1796_rst;
  logic [31:0] f1796_rdata;
  sr_buffer_32_1 f1796(.wen(f1796_wen), .wdata(f1796_wdata), .clk(f1796_clk), .rst(f1796_rst), .rdata(f1796_rdata));
  assign f1796_clk = clk;
  assign f1796_rst = rst;
  // Bindings to f1796

  // f1798
  logic [0:0] f1798_wen;
  logic [31:0] f1798_wdata;
  logic [0:0] f1798_clk;
  logic [0:0] f1798_rst;
  logic [31:0] f1798_rdata;
  sr_buffer_32_1 f1798(.wen(f1798_wen), .wdata(f1798_wdata), .clk(f1798_clk), .rst(f1798_rst), .rdata(f1798_rdata));
  assign f1798_clk = clk;
  assign f1798_rst = rst;
  // Bindings to f1798

  // f1800
  logic [0:0] f1800_wen;
  logic [31:0] f1800_wdata;
  logic [0:0] f1800_clk;
  logic [0:0] f1800_rst;
  logic [31:0] f1800_rdata;
  sr_buffer_32_1 f1800(.wen(f1800_wen), .wdata(f1800_wdata), .clk(f1800_clk), .rst(f1800_rst), .rdata(f1800_rdata));
  assign f1800_clk = clk;
  assign f1800_rst = rst;
  // Bindings to f1800

  // f1802
  logic [0:0] f1802_wen;
  logic [31:0] f1802_wdata;
  logic [0:0] f1802_clk;
  logic [0:0] f1802_rst;
  logic [31:0] f1802_rdata;
  sr_buffer_32_1 f1802(.wen(f1802_wen), .wdata(f1802_wdata), .clk(f1802_clk), .rst(f1802_rst), .rdata(f1802_rdata));
  assign f1802_clk = clk;
  assign f1802_rst = rst;
  // Bindings to f1802

  // f1804
  logic [0:0] f1804_wen;
  logic [31:0] f1804_wdata;
  logic [0:0] f1804_clk;
  logic [0:0] f1804_rst;
  logic [31:0] f1804_rdata;
  sr_buffer_32_1 f1804(.wen(f1804_wen), .wdata(f1804_wdata), .clk(f1804_clk), .rst(f1804_rst), .rdata(f1804_rdata));
  assign f1804_clk = clk;
  assign f1804_rst = rst;
  // Bindings to f1804

  // f1806
  logic [0:0] f1806_wen;
  logic [31:0] f1806_wdata;
  logic [0:0] f1806_clk;
  logic [0:0] f1806_rst;
  logic [31:0] f1806_rdata;
  sr_buffer_32_1 f1806(.wen(f1806_wen), .wdata(f1806_wdata), .clk(f1806_clk), .rst(f1806_rst), .rdata(f1806_rdata));
  assign f1806_clk = clk;
  assign f1806_rst = rst;
  // Bindings to f1806

  // f1808
  logic [0:0] f1808_wen;
  logic [31:0] f1808_wdata;
  logic [0:0] f1808_clk;
  logic [0:0] f1808_rst;
  logic [31:0] f1808_rdata;
  sr_buffer_32_1 f1808(.wen(f1808_wen), .wdata(f1808_wdata), .clk(f1808_clk), .rst(f1808_rst), .rdata(f1808_rdata));
  assign f1808_clk = clk;
  assign f1808_rst = rst;
  // Bindings to f1808

  // f1810
  logic [0:0] f1810_wen;
  logic [31:0] f1810_wdata;
  logic [0:0] f1810_clk;
  logic [0:0] f1810_rst;
  logic [31:0] f1810_rdata;
  sr_buffer_32_1 f1810(.wen(f1810_wen), .wdata(f1810_wdata), .clk(f1810_clk), .rst(f1810_rst), .rdata(f1810_rdata));
  assign f1810_clk = clk;
  assign f1810_rst = rst;
  // Bindings to f1810

  // f1812
  logic [0:0] f1812_wen;
  logic [31:0] f1812_wdata;
  logic [0:0] f1812_clk;
  logic [0:0] f1812_rst;
  logic [31:0] f1812_rdata;
  sr_buffer_32_1 f1812(.wen(f1812_wen), .wdata(f1812_wdata), .clk(f1812_clk), .rst(f1812_rst), .rdata(f1812_rdata));
  assign f1812_clk = clk;
  assign f1812_rst = rst;
  // Bindings to f1812

  // f1814
  logic [0:0] f1814_wen;
  logic [31:0] f1814_wdata;
  logic [0:0] f1814_clk;
  logic [0:0] f1814_rst;
  logic [31:0] f1814_rdata;
  sr_buffer_32_1 f1814(.wen(f1814_wen), .wdata(f1814_wdata), .clk(f1814_clk), .rst(f1814_rst), .rdata(f1814_rdata));
  assign f1814_clk = clk;
  assign f1814_rst = rst;
  // Bindings to f1814

  // f1816
  logic [0:0] f1816_wen;
  logic [31:0] f1816_wdata;
  logic [0:0] f1816_clk;
  logic [0:0] f1816_rst;
  logic [31:0] f1816_rdata;
  sr_buffer_32_1 f1816(.wen(f1816_wen), .wdata(f1816_wdata), .clk(f1816_clk), .rst(f1816_rst), .rdata(f1816_rdata));
  assign f1816_clk = clk;
  assign f1816_rst = rst;
  // Bindings to f1816

  // f1818
  logic [0:0] f1818_wen;
  logic [31:0] f1818_wdata;
  logic [0:0] f1818_clk;
  logic [0:0] f1818_rst;
  logic [31:0] f1818_rdata;
  sr_buffer_32_1 f1818(.wen(f1818_wen), .wdata(f1818_wdata), .clk(f1818_clk), .rst(f1818_rst), .rdata(f1818_rdata));
  assign f1818_clk = clk;
  assign f1818_rst = rst;
  // Bindings to f1818

  // f1820
  logic [0:0] f1820_wen;
  logic [31:0] f1820_wdata;
  logic [0:0] f1820_clk;
  logic [0:0] f1820_rst;
  logic [31:0] f1820_rdata;
  sr_buffer_32_1 f1820(.wen(f1820_wen), .wdata(f1820_wdata), .clk(f1820_clk), .rst(f1820_rst), .rdata(f1820_rdata));
  assign f1820_clk = clk;
  assign f1820_rst = rst;
  // Bindings to f1820

  // f1822
  logic [0:0] f1822_wen;
  logic [31:0] f1822_wdata;
  logic [0:0] f1822_clk;
  logic [0:0] f1822_rst;
  logic [31:0] f1822_rdata;
  sr_buffer_32_1 f1822(.wen(f1822_wen), .wdata(f1822_wdata), .clk(f1822_clk), .rst(f1822_rst), .rdata(f1822_rdata));
  assign f1822_clk = clk;
  assign f1822_rst = rst;
  // Bindings to f1822

  // f1824
  logic [0:0] f1824_wen;
  logic [31:0] f1824_wdata;
  logic [0:0] f1824_clk;
  logic [0:0] f1824_rst;
  logic [31:0] f1824_rdata;
  sr_buffer_32_1 f1824(.wen(f1824_wen), .wdata(f1824_wdata), .clk(f1824_clk), .rst(f1824_rst), .rdata(f1824_rdata));
  assign f1824_clk = clk;
  assign f1824_rst = rst;
  // Bindings to f1824

  // f1826
  logic [0:0] f1826_wen;
  logic [31:0] f1826_wdata;
  logic [0:0] f1826_clk;
  logic [0:0] f1826_rst;
  logic [31:0] f1826_rdata;
  sr_buffer_32_1 f1826(.wen(f1826_wen), .wdata(f1826_wdata), .clk(f1826_clk), .rst(f1826_rst), .rdata(f1826_rdata));
  assign f1826_clk = clk;
  assign f1826_rst = rst;
  // Bindings to f1826

  // f1828
  logic [0:0] f1828_wen;
  logic [31:0] f1828_wdata;
  logic [0:0] f1828_clk;
  logic [0:0] f1828_rst;
  logic [31:0] f1828_rdata;
  sr_buffer_32_1 f1828(.wen(f1828_wen), .wdata(f1828_wdata), .clk(f1828_clk), .rst(f1828_rst), .rdata(f1828_rdata));
  assign f1828_clk = clk;
  assign f1828_rst = rst;
  // Bindings to f1828

  // f1830
  logic [0:0] f1830_wen;
  logic [31:0] f1830_wdata;
  logic [0:0] f1830_clk;
  logic [0:0] f1830_rst;
  logic [31:0] f1830_rdata;
  sr_buffer_32_1 f1830(.wen(f1830_wen), .wdata(f1830_wdata), .clk(f1830_clk), .rst(f1830_rst), .rdata(f1830_rdata));
  assign f1830_clk = clk;
  assign f1830_rst = rst;
  // Bindings to f1830

  // f1832
  logic [0:0] f1832_wen;
  logic [31:0] f1832_wdata;
  logic [0:0] f1832_clk;
  logic [0:0] f1832_rst;
  logic [31:0] f1832_rdata;
  sr_buffer_32_1 f1832(.wen(f1832_wen), .wdata(f1832_wdata), .clk(f1832_clk), .rst(f1832_rst), .rdata(f1832_rdata));
  assign f1832_clk = clk;
  assign f1832_rst = rst;
  // Bindings to f1832

  // f1834
  logic [0:0] f1834_wen;
  logic [31:0] f1834_wdata;
  logic [0:0] f1834_clk;
  logic [0:0] f1834_rst;
  logic [31:0] f1834_rdata;
  sr_buffer_32_1 f1834(.wen(f1834_wen), .wdata(f1834_wdata), .clk(f1834_clk), .rst(f1834_rst), .rdata(f1834_rdata));
  assign f1834_clk = clk;
  assign f1834_rst = rst;
  // Bindings to f1834

  // f1836
  logic [0:0] f1836_wen;
  logic [31:0] f1836_wdata;
  logic [0:0] f1836_clk;
  logic [0:0] f1836_rst;
  logic [31:0] f1836_rdata;
  sr_buffer_32_1 f1836(.wen(f1836_wen), .wdata(f1836_wdata), .clk(f1836_clk), .rst(f1836_rst), .rdata(f1836_rdata));
  assign f1836_clk = clk;
  assign f1836_rst = rst;
  // Bindings to f1836

  // f1838
  logic [0:0] f1838_wen;
  logic [31:0] f1838_wdata;
  logic [0:0] f1838_clk;
  logic [0:0] f1838_rst;
  logic [31:0] f1838_rdata;
  sr_buffer_32_1 f1838(.wen(f1838_wen), .wdata(f1838_wdata), .clk(f1838_clk), .rst(f1838_rst), .rdata(f1838_rdata));
  assign f1838_clk = clk;
  assign f1838_rst = rst;
  // Bindings to f1838

  // f1840
  logic [0:0] f1840_wen;
  logic [31:0] f1840_wdata;
  logic [0:0] f1840_clk;
  logic [0:0] f1840_rst;
  logic [31:0] f1840_rdata;
  sr_buffer_32_1 f1840(.wen(f1840_wen), .wdata(f1840_wdata), .clk(f1840_clk), .rst(f1840_rst), .rdata(f1840_rdata));
  assign f1840_clk = clk;
  assign f1840_rst = rst;
  // Bindings to f1840

  // f1842
  logic [0:0] f1842_wen;
  logic [31:0] f1842_wdata;
  logic [0:0] f1842_clk;
  logic [0:0] f1842_rst;
  logic [31:0] f1842_rdata;
  sr_buffer_32_1 f1842(.wen(f1842_wen), .wdata(f1842_wdata), .clk(f1842_clk), .rst(f1842_rst), .rdata(f1842_rdata));
  assign f1842_clk = clk;
  assign f1842_rst = rst;
  // Bindings to f1842

  // f1844
  logic [0:0] f1844_wen;
  logic [31:0] f1844_wdata;
  logic [0:0] f1844_clk;
  logic [0:0] f1844_rst;
  logic [31:0] f1844_rdata;
  sr_buffer_32_1 f1844(.wen(f1844_wen), .wdata(f1844_wdata), .clk(f1844_clk), .rst(f1844_rst), .rdata(f1844_rdata));
  assign f1844_clk = clk;
  assign f1844_rst = rst;
  // Bindings to f1844

  // f1846
  logic [0:0] f1846_wen;
  logic [31:0] f1846_wdata;
  logic [0:0] f1846_clk;
  logic [0:0] f1846_rst;
  logic [31:0] f1846_rdata;
  sr_buffer_32_1 f1846(.wen(f1846_wen), .wdata(f1846_wdata), .clk(f1846_clk), .rst(f1846_rst), .rdata(f1846_rdata));
  assign f1846_clk = clk;
  assign f1846_rst = rst;
  // Bindings to f1846

  // f1848
  logic [0:0] f1848_wen;
  logic [31:0] f1848_wdata;
  logic [0:0] f1848_clk;
  logic [0:0] f1848_rst;
  logic [31:0] f1848_rdata;
  sr_buffer_32_1 f1848(.wen(f1848_wen), .wdata(f1848_wdata), .clk(f1848_clk), .rst(f1848_rst), .rdata(f1848_rdata));
  assign f1848_clk = clk;
  assign f1848_rst = rst;
  // Bindings to f1848

  // f1850
  logic [0:0] f1850_wen;
  logic [31:0] f1850_wdata;
  logic [0:0] f1850_clk;
  logic [0:0] f1850_rst;
  logic [31:0] f1850_rdata;
  sr_buffer_32_1 f1850(.wen(f1850_wen), .wdata(f1850_wdata), .clk(f1850_clk), .rst(f1850_rst), .rdata(f1850_rdata));
  assign f1850_clk = clk;
  assign f1850_rst = rst;
  // Bindings to f1850

  // f1852
  logic [0:0] f1852_wen;
  logic [31:0] f1852_wdata;
  logic [0:0] f1852_clk;
  logic [0:0] f1852_rst;
  logic [31:0] f1852_rdata;
  sr_buffer_32_1 f1852(.wen(f1852_wen), .wdata(f1852_wdata), .clk(f1852_clk), .rst(f1852_rst), .rdata(f1852_rdata));
  assign f1852_clk = clk;
  assign f1852_rst = rst;
  // Bindings to f1852

  // f1854
  logic [0:0] f1854_wen;
  logic [31:0] f1854_wdata;
  logic [0:0] f1854_clk;
  logic [0:0] f1854_rst;
  logic [31:0] f1854_rdata;
  sr_buffer_32_1 f1854(.wen(f1854_wen), .wdata(f1854_wdata), .clk(f1854_clk), .rst(f1854_rst), .rdata(f1854_rdata));
  assign f1854_clk = clk;
  assign f1854_rst = rst;
  // Bindings to f1854

  // f1856
  logic [0:0] f1856_wen;
  logic [31:0] f1856_wdata;
  logic [0:0] f1856_clk;
  logic [0:0] f1856_rst;
  logic [31:0] f1856_rdata;
  sr_buffer_32_1 f1856(.wen(f1856_wen), .wdata(f1856_wdata), .clk(f1856_clk), .rst(f1856_rst), .rdata(f1856_rdata));
  assign f1856_clk = clk;
  assign f1856_rst = rst;
  // Bindings to f1856

  // f1858
  logic [0:0] f1858_wen;
  logic [31:0] f1858_wdata;
  logic [0:0] f1858_clk;
  logic [0:0] f1858_rst;
  logic [31:0] f1858_rdata;
  sr_buffer_32_1 f1858(.wen(f1858_wen), .wdata(f1858_wdata), .clk(f1858_clk), .rst(f1858_rst), .rdata(f1858_rdata));
  assign f1858_clk = clk;
  assign f1858_rst = rst;
  // Bindings to f1858

  // f1860
  logic [0:0] f1860_wen;
  logic [31:0] f1860_wdata;
  logic [0:0] f1860_clk;
  logic [0:0] f1860_rst;
  logic [31:0] f1860_rdata;
  sr_buffer_32_1 f1860(.wen(f1860_wen), .wdata(f1860_wdata), .clk(f1860_clk), .rst(f1860_rst), .rdata(f1860_rdata));
  assign f1860_clk = clk;
  assign f1860_rst = rst;
  // Bindings to f1860

  // f1862
  logic [0:0] f1862_wen;
  logic [31:0] f1862_wdata;
  logic [0:0] f1862_clk;
  logic [0:0] f1862_rst;
  logic [31:0] f1862_rdata;
  sr_buffer_32_1 f1862(.wen(f1862_wen), .wdata(f1862_wdata), .clk(f1862_clk), .rst(f1862_rst), .rdata(f1862_rdata));
  assign f1862_clk = clk;
  assign f1862_rst = rst;
  // Bindings to f1862

  // f1864
  logic [0:0] f1864_wen;
  logic [31:0] f1864_wdata;
  logic [0:0] f1864_clk;
  logic [0:0] f1864_rst;
  logic [31:0] f1864_rdata;
  sr_buffer_32_1 f1864(.wen(f1864_wen), .wdata(f1864_wdata), .clk(f1864_clk), .rst(f1864_rst), .rdata(f1864_rdata));
  assign f1864_clk = clk;
  assign f1864_rst = rst;
  // Bindings to f1864

  // f1866
  logic [0:0] f1866_wen;
  logic [31:0] f1866_wdata;
  logic [0:0] f1866_clk;
  logic [0:0] f1866_rst;
  logic [31:0] f1866_rdata;
  sr_buffer_32_1 f1866(.wen(f1866_wen), .wdata(f1866_wdata), .clk(f1866_clk), .rst(f1866_rst), .rdata(f1866_rdata));
  assign f1866_clk = clk;
  assign f1866_rst = rst;
  // Bindings to f1866

  // f1868
  logic [0:0] f1868_wen;
  logic [31:0] f1868_wdata;
  logic [0:0] f1868_clk;
  logic [0:0] f1868_rst;
  logic [31:0] f1868_rdata;
  sr_buffer_32_1 f1868(.wen(f1868_wen), .wdata(f1868_wdata), .clk(f1868_clk), .rst(f1868_rst), .rdata(f1868_rdata));
  assign f1868_clk = clk;
  assign f1868_rst = rst;
  // Bindings to f1868

  // f1870
  logic [0:0] f1870_wen;
  logic [31:0] f1870_wdata;
  logic [0:0] f1870_clk;
  logic [0:0] f1870_rst;
  logic [31:0] f1870_rdata;
  sr_buffer_32_1 f1870(.wen(f1870_wen), .wdata(f1870_wdata), .clk(f1870_clk), .rst(f1870_rst), .rdata(f1870_rdata));
  assign f1870_clk = clk;
  assign f1870_rst = rst;
  // Bindings to f1870

  // f1872
  logic [0:0] f1872_wen;
  logic [31:0] f1872_wdata;
  logic [0:0] f1872_clk;
  logic [0:0] f1872_rst;
  logic [31:0] f1872_rdata;
  sr_buffer_32_1 f1872(.wen(f1872_wen), .wdata(f1872_wdata), .clk(f1872_clk), .rst(f1872_rst), .rdata(f1872_rdata));
  assign f1872_clk = clk;
  assign f1872_rst = rst;
  // Bindings to f1872

  // f1874
  logic [0:0] f1874_wen;
  logic [31:0] f1874_wdata;
  logic [0:0] f1874_clk;
  logic [0:0] f1874_rst;
  logic [31:0] f1874_rdata;
  sr_buffer_32_1 f1874(.wen(f1874_wen), .wdata(f1874_wdata), .clk(f1874_clk), .rst(f1874_rst), .rdata(f1874_rdata));
  assign f1874_clk = clk;
  assign f1874_rst = rst;
  // Bindings to f1874

  // f1876
  logic [0:0] f1876_wen;
  logic [31:0] f1876_wdata;
  logic [0:0] f1876_clk;
  logic [0:0] f1876_rst;
  logic [31:0] f1876_rdata;
  sr_buffer_32_1 f1876(.wen(f1876_wen), .wdata(f1876_wdata), .clk(f1876_clk), .rst(f1876_rst), .rdata(f1876_rdata));
  assign f1876_clk = clk;
  assign f1876_rst = rst;
  // Bindings to f1876

  // f1878
  logic [0:0] f1878_wen;
  logic [31:0] f1878_wdata;
  logic [0:0] f1878_clk;
  logic [0:0] f1878_rst;
  logic [31:0] f1878_rdata;
  sr_buffer_32_1 f1878(.wen(f1878_wen), .wdata(f1878_wdata), .clk(f1878_clk), .rst(f1878_rst), .rdata(f1878_rdata));
  assign f1878_clk = clk;
  assign f1878_rst = rst;
  // Bindings to f1878

  // f1880
  logic [0:0] f1880_wen;
  logic [31:0] f1880_wdata;
  logic [0:0] f1880_clk;
  logic [0:0] f1880_rst;
  logic [31:0] f1880_rdata;
  sr_buffer_32_1 f1880(.wen(f1880_wen), .wdata(f1880_wdata), .clk(f1880_clk), .rst(f1880_rst), .rdata(f1880_rdata));
  assign f1880_clk = clk;
  assign f1880_rst = rst;
  // Bindings to f1880

  // f1882
  logic [0:0] f1882_wen;
  logic [31:0] f1882_wdata;
  logic [0:0] f1882_clk;
  logic [0:0] f1882_rst;
  logic [31:0] f1882_rdata;
  sr_buffer_32_1 f1882(.wen(f1882_wen), .wdata(f1882_wdata), .clk(f1882_clk), .rst(f1882_rst), .rdata(f1882_rdata));
  assign f1882_clk = clk;
  assign f1882_rst = rst;
  // Bindings to f1882

  // f1884
  logic [0:0] f1884_wen;
  logic [31:0] f1884_wdata;
  logic [0:0] f1884_clk;
  logic [0:0] f1884_rst;
  logic [31:0] f1884_rdata;
  sr_buffer_32_1 f1884(.wen(f1884_wen), .wdata(f1884_wdata), .clk(f1884_clk), .rst(f1884_rst), .rdata(f1884_rdata));
  assign f1884_clk = clk;
  assign f1884_rst = rst;
  // Bindings to f1884

  // f1886
  logic [0:0] f1886_wen;
  logic [31:0] f1886_wdata;
  logic [0:0] f1886_clk;
  logic [0:0] f1886_rst;
  logic [31:0] f1886_rdata;
  sr_buffer_32_1 f1886(.wen(f1886_wen), .wdata(f1886_wdata), .clk(f1886_clk), .rst(f1886_rst), .rdata(f1886_rdata));
  assign f1886_clk = clk;
  assign f1886_rst = rst;
  // Bindings to f1886

  // f1888
  logic [0:0] f1888_wen;
  logic [31:0] f1888_wdata;
  logic [0:0] f1888_clk;
  logic [0:0] f1888_rst;
  logic [31:0] f1888_rdata;
  sr_buffer_32_1 f1888(.wen(f1888_wen), .wdata(f1888_wdata), .clk(f1888_clk), .rst(f1888_rst), .rdata(f1888_rdata));
  assign f1888_clk = clk;
  assign f1888_rst = rst;
  // Bindings to f1888

  // f1890
  logic [0:0] f1890_wen;
  logic [31:0] f1890_wdata;
  logic [0:0] f1890_clk;
  logic [0:0] f1890_rst;
  logic [31:0] f1890_rdata;
  sr_buffer_32_1 f1890(.wen(f1890_wen), .wdata(f1890_wdata), .clk(f1890_clk), .rst(f1890_rst), .rdata(f1890_rdata));
  assign f1890_clk = clk;
  assign f1890_rst = rst;
  // Bindings to f1890

  // f1892
  logic [0:0] f1892_wen;
  logic [31:0] f1892_wdata;
  logic [0:0] f1892_clk;
  logic [0:0] f1892_rst;
  logic [31:0] f1892_rdata;
  sr_buffer_32_1 f1892(.wen(f1892_wen), .wdata(f1892_wdata), .clk(f1892_clk), .rst(f1892_rst), .rdata(f1892_rdata));
  assign f1892_clk = clk;
  assign f1892_rst = rst;
  // Bindings to f1892

  // f1894
  logic [0:0] f1894_wen;
  logic [31:0] f1894_wdata;
  logic [0:0] f1894_clk;
  logic [0:0] f1894_rst;
  logic [31:0] f1894_rdata;
  sr_buffer_32_1 f1894(.wen(f1894_wen), .wdata(f1894_wdata), .clk(f1894_clk), .rst(f1894_rst), .rdata(f1894_rdata));
  assign f1894_clk = clk;
  assign f1894_rst = rst;
  // Bindings to f1894

  // f1896
  logic [0:0] f1896_wen;
  logic [31:0] f1896_wdata;
  logic [0:0] f1896_clk;
  logic [0:0] f1896_rst;
  logic [31:0] f1896_rdata;
  sr_buffer_32_1 f1896(.wen(f1896_wen), .wdata(f1896_wdata), .clk(f1896_clk), .rst(f1896_rst), .rdata(f1896_rdata));
  assign f1896_clk = clk;
  assign f1896_rst = rst;
  // Bindings to f1896

  // f1898
  logic [0:0] f1898_wen;
  logic [31:0] f1898_wdata;
  logic [0:0] f1898_clk;
  logic [0:0] f1898_rst;
  logic [31:0] f1898_rdata;
  sr_buffer_32_1 f1898(.wen(f1898_wen), .wdata(f1898_wdata), .clk(f1898_clk), .rst(f1898_rst), .rdata(f1898_rdata));
  assign f1898_clk = clk;
  assign f1898_rst = rst;
  // Bindings to f1898

  // f1900
  logic [0:0] f1900_wen;
  logic [31:0] f1900_wdata;
  logic [0:0] f1900_clk;
  logic [0:0] f1900_rst;
  logic [31:0] f1900_rdata;
  sr_buffer_32_1 f1900(.wen(f1900_wen), .wdata(f1900_wdata), .clk(f1900_clk), .rst(f1900_rst), .rdata(f1900_rdata));
  assign f1900_clk = clk;
  assign f1900_rst = rst;
  // Bindings to f1900

  // f1902
  logic [0:0] f1902_wen;
  logic [31:0] f1902_wdata;
  logic [0:0] f1902_clk;
  logic [0:0] f1902_rst;
  logic [31:0] f1902_rdata;
  sr_buffer_32_1 f1902(.wen(f1902_wen), .wdata(f1902_wdata), .clk(f1902_clk), .rst(f1902_rst), .rdata(f1902_rdata));
  assign f1902_clk = clk;
  assign f1902_rst = rst;
  // Bindings to f1902

  // f1904
  logic [0:0] f1904_wen;
  logic [31:0] f1904_wdata;
  logic [0:0] f1904_clk;
  logic [0:0] f1904_rst;
  logic [31:0] f1904_rdata;
  sr_buffer_32_1 f1904(.wen(f1904_wen), .wdata(f1904_wdata), .clk(f1904_clk), .rst(f1904_rst), .rdata(f1904_rdata));
  assign f1904_clk = clk;
  assign f1904_rst = rst;
  // Bindings to f1904

  // f1906
  logic [0:0] f1906_wen;
  logic [31:0] f1906_wdata;
  logic [0:0] f1906_clk;
  logic [0:0] f1906_rst;
  logic [31:0] f1906_rdata;
  sr_buffer_32_1 f1906(.wen(f1906_wen), .wdata(f1906_wdata), .clk(f1906_clk), .rst(f1906_rst), .rdata(f1906_rdata));
  assign f1906_clk = clk;
  assign f1906_rst = rst;
  // Bindings to f1906

  // f1908
  logic [0:0] f1908_wen;
  logic [31:0] f1908_wdata;
  logic [0:0] f1908_clk;
  logic [0:0] f1908_rst;
  logic [31:0] f1908_rdata;
  sr_buffer_32_1 f1908(.wen(f1908_wen), .wdata(f1908_wdata), .clk(f1908_clk), .rst(f1908_rst), .rdata(f1908_rdata));
  assign f1908_clk = clk;
  assign f1908_rst = rst;
  // Bindings to f1908

  // f1910
  logic [0:0] f1910_wen;
  logic [31:0] f1910_wdata;
  logic [0:0] f1910_clk;
  logic [0:0] f1910_rst;
  logic [31:0] f1910_rdata;
  sr_buffer_32_1 f1910(.wen(f1910_wen), .wdata(f1910_wdata), .clk(f1910_clk), .rst(f1910_rst), .rdata(f1910_rdata));
  assign f1910_clk = clk;
  assign f1910_rst = rst;
  // Bindings to f1910

  // f1912
  logic [0:0] f1912_wen;
  logic [31:0] f1912_wdata;
  logic [0:0] f1912_clk;
  logic [0:0] f1912_rst;
  logic [31:0] f1912_rdata;
  sr_buffer_32_1 f1912(.wen(f1912_wen), .wdata(f1912_wdata), .clk(f1912_clk), .rst(f1912_rst), .rdata(f1912_rdata));
  assign f1912_clk = clk;
  assign f1912_rst = rst;
  // Bindings to f1912

  // f1914
  logic [0:0] f1914_wen;
  logic [31:0] f1914_wdata;
  logic [0:0] f1914_clk;
  logic [0:0] f1914_rst;
  logic [31:0] f1914_rdata;
  sr_buffer_32_1 f1914(.wen(f1914_wen), .wdata(f1914_wdata), .clk(f1914_clk), .rst(f1914_rst), .rdata(f1914_rdata));
  assign f1914_clk = clk;
  assign f1914_rst = rst;
  // Bindings to f1914

  // f1916
  logic [0:0] f1916_wen;
  logic [31:0] f1916_wdata;
  logic [0:0] f1916_clk;
  logic [0:0] f1916_rst;
  logic [31:0] f1916_rdata;
  sr_buffer_32_1 f1916(.wen(f1916_wen), .wdata(f1916_wdata), .clk(f1916_clk), .rst(f1916_rst), .rdata(f1916_rdata));
  assign f1916_clk = clk;
  assign f1916_rst = rst;
  // Bindings to f1916

  // f1918
  logic [0:0] f1918_wen;
  logic [31:0] f1918_wdata;
  logic [0:0] f1918_clk;
  logic [0:0] f1918_rst;
  logic [31:0] f1918_rdata;
  sr_buffer_32_1 f1918(.wen(f1918_wen), .wdata(f1918_wdata), .clk(f1918_clk), .rst(f1918_rst), .rdata(f1918_rdata));
  assign f1918_clk = clk;
  assign f1918_rst = rst;
  // Bindings to f1918

  // f1920
  logic [0:0] f1920_wen;
  logic [31:0] f1920_wdata;
  logic [0:0] f1920_clk;
  logic [0:0] f1920_rst;
  logic [31:0] f1920_rdata;
  sr_buffer_32_1 f1920(.wen(f1920_wen), .wdata(f1920_wdata), .clk(f1920_clk), .rst(f1920_rst), .rdata(f1920_rdata));
  assign f1920_clk = clk;
  assign f1920_rst = rst;
  // Bindings to f1920

  // f1922
  logic [0:0] f1922_wen;
  logic [31:0] f1922_wdata;
  logic [0:0] f1922_clk;
  logic [0:0] f1922_rst;
  logic [31:0] f1922_rdata;
  sr_buffer_32_1 f1922(.wen(f1922_wen), .wdata(f1922_wdata), .clk(f1922_clk), .rst(f1922_rst), .rdata(f1922_rdata));
  assign f1922_clk = clk;
  assign f1922_rst = rst;
  // Bindings to f1922

  // f1924
  logic [0:0] f1924_wen;
  logic [31:0] f1924_wdata;
  logic [0:0] f1924_clk;
  logic [0:0] f1924_rst;
  logic [31:0] f1924_rdata;
  sr_buffer_32_1 f1924(.wen(f1924_wen), .wdata(f1924_wdata), .clk(f1924_clk), .rst(f1924_rst), .rdata(f1924_rdata));
  assign f1924_clk = clk;
  assign f1924_rst = rst;
  // Bindings to f1924

  // f1926
  logic [0:0] f1926_wen;
  logic [31:0] f1926_wdata;
  logic [0:0] f1926_clk;
  logic [0:0] f1926_rst;
  logic [31:0] f1926_rdata;
  sr_buffer_32_1 f1926(.wen(f1926_wen), .wdata(f1926_wdata), .clk(f1926_clk), .rst(f1926_rst), .rdata(f1926_rdata));
  assign f1926_clk = clk;
  assign f1926_rst = rst;
  // Bindings to f1926

  // f1928
  logic [0:0] f1928_wen;
  logic [31:0] f1928_wdata;
  logic [0:0] f1928_clk;
  logic [0:0] f1928_rst;
  logic [31:0] f1928_rdata;
  sr_buffer_32_1 f1928(.wen(f1928_wen), .wdata(f1928_wdata), .clk(f1928_clk), .rst(f1928_rst), .rdata(f1928_rdata));
  assign f1928_clk = clk;
  assign f1928_rst = rst;
  // Bindings to f1928

  // f1930
  logic [0:0] f1930_wen;
  logic [31:0] f1930_wdata;
  logic [0:0] f1930_clk;
  logic [0:0] f1930_rst;
  logic [31:0] f1930_rdata;
  sr_buffer_32_1 f1930(.wen(f1930_wen), .wdata(f1930_wdata), .clk(f1930_clk), .rst(f1930_rst), .rdata(f1930_rdata));
  assign f1930_clk = clk;
  assign f1930_rst = rst;
  // Bindings to f1930

  // f1932
  logic [0:0] f1932_wen;
  logic [31:0] f1932_wdata;
  logic [0:0] f1932_clk;
  logic [0:0] f1932_rst;
  logic [31:0] f1932_rdata;
  sr_buffer_32_1 f1932(.wen(f1932_wen), .wdata(f1932_wdata), .clk(f1932_clk), .rst(f1932_rst), .rdata(f1932_rdata));
  assign f1932_clk = clk;
  assign f1932_rst = rst;
  // Bindings to f1932

  // f1934
  logic [0:0] f1934_wen;
  logic [31:0] f1934_wdata;
  logic [0:0] f1934_clk;
  logic [0:0] f1934_rst;
  logic [31:0] f1934_rdata;
  sr_buffer_32_1 f1934(.wen(f1934_wen), .wdata(f1934_wdata), .clk(f1934_clk), .rst(f1934_rst), .rdata(f1934_rdata));
  assign f1934_clk = clk;
  assign f1934_rst = rst;
  // Bindings to f1934

  // f1936
  logic [0:0] f1936_wen;
  logic [31:0] f1936_wdata;
  logic [0:0] f1936_clk;
  logic [0:0] f1936_rst;
  logic [31:0] f1936_rdata;
  sr_buffer_32_1 f1936(.wen(f1936_wen), .wdata(f1936_wdata), .clk(f1936_clk), .rst(f1936_rst), .rdata(f1936_rdata));
  assign f1936_clk = clk;
  assign f1936_rst = rst;
  // Bindings to f1936

  // f1938
  logic [0:0] f1938_wen;
  logic [31:0] f1938_wdata;
  logic [0:0] f1938_clk;
  logic [0:0] f1938_rst;
  logic [31:0] f1938_rdata;
  sr_buffer_32_1 f1938(.wen(f1938_wen), .wdata(f1938_wdata), .clk(f1938_clk), .rst(f1938_rst), .rdata(f1938_rdata));
  assign f1938_clk = clk;
  assign f1938_rst = rst;
  // Bindings to f1938

  // f1940
  logic [0:0] f1940_wen;
  logic [31:0] f1940_wdata;
  logic [0:0] f1940_clk;
  logic [0:0] f1940_rst;
  logic [31:0] f1940_rdata;
  sr_buffer_32_1 f1940(.wen(f1940_wen), .wdata(f1940_wdata), .clk(f1940_clk), .rst(f1940_rst), .rdata(f1940_rdata));
  assign f1940_clk = clk;
  assign f1940_rst = rst;
  // Bindings to f1940

  // f1942
  logic [0:0] f1942_wen;
  logic [31:0] f1942_wdata;
  logic [0:0] f1942_clk;
  logic [0:0] f1942_rst;
  logic [31:0] f1942_rdata;
  sr_buffer_32_1 f1942(.wen(f1942_wen), .wdata(f1942_wdata), .clk(f1942_clk), .rst(f1942_rst), .rdata(f1942_rdata));
  assign f1942_clk = clk;
  assign f1942_rst = rst;
  // Bindings to f1942

  // f1944
  logic [0:0] f1944_wen;
  logic [31:0] f1944_wdata;
  logic [0:0] f1944_clk;
  logic [0:0] f1944_rst;
  logic [31:0] f1944_rdata;
  sr_buffer_32_1 f1944(.wen(f1944_wen), .wdata(f1944_wdata), .clk(f1944_clk), .rst(f1944_rst), .rdata(f1944_rdata));
  assign f1944_clk = clk;
  assign f1944_rst = rst;
  // Bindings to f1944

  // f1946
  logic [0:0] f1946_wen;
  logic [31:0] f1946_wdata;
  logic [0:0] f1946_clk;
  logic [0:0] f1946_rst;
  logic [31:0] f1946_rdata;
  sr_buffer_32_1 f1946(.wen(f1946_wen), .wdata(f1946_wdata), .clk(f1946_clk), .rst(f1946_rst), .rdata(f1946_rdata));
  assign f1946_clk = clk;
  assign f1946_rst = rst;
  // Bindings to f1946

  // f1948
  logic [0:0] f1948_wen;
  logic [31:0] f1948_wdata;
  logic [0:0] f1948_clk;
  logic [0:0] f1948_rst;
  logic [31:0] f1948_rdata;
  sr_buffer_32_1 f1948(.wen(f1948_wen), .wdata(f1948_wdata), .clk(f1948_clk), .rst(f1948_rst), .rdata(f1948_rdata));
  assign f1948_clk = clk;
  assign f1948_rst = rst;
  // Bindings to f1948

  // f1950
  logic [0:0] f1950_wen;
  logic [31:0] f1950_wdata;
  logic [0:0] f1950_clk;
  logic [0:0] f1950_rst;
  logic [31:0] f1950_rdata;
  sr_buffer_32_1 f1950(.wen(f1950_wen), .wdata(f1950_wdata), .clk(f1950_clk), .rst(f1950_rst), .rdata(f1950_rdata));
  assign f1950_clk = clk;
  assign f1950_rst = rst;
  // Bindings to f1950

  // f1952
  logic [0:0] f1952_wen;
  logic [31:0] f1952_wdata;
  logic [0:0] f1952_clk;
  logic [0:0] f1952_rst;
  logic [31:0] f1952_rdata;
  sr_buffer_32_1 f1952(.wen(f1952_wen), .wdata(f1952_wdata), .clk(f1952_clk), .rst(f1952_rst), .rdata(f1952_rdata));
  assign f1952_clk = clk;
  assign f1952_rst = rst;
  // Bindings to f1952

  // f1954
  logic [0:0] f1954_wen;
  logic [31:0] f1954_wdata;
  logic [0:0] f1954_clk;
  logic [0:0] f1954_rst;
  logic [31:0] f1954_rdata;
  sr_buffer_32_1 f1954(.wen(f1954_wen), .wdata(f1954_wdata), .clk(f1954_clk), .rst(f1954_rst), .rdata(f1954_rdata));
  assign f1954_clk = clk;
  assign f1954_rst = rst;
  // Bindings to f1954

  // f1956
  logic [0:0] f1956_wen;
  logic [31:0] f1956_wdata;
  logic [0:0] f1956_clk;
  logic [0:0] f1956_rst;
  logic [31:0] f1956_rdata;
  sr_buffer_32_1 f1956(.wen(f1956_wen), .wdata(f1956_wdata), .clk(f1956_clk), .rst(f1956_rst), .rdata(f1956_rdata));
  assign f1956_clk = clk;
  assign f1956_rst = rst;
  // Bindings to f1956

  // f1958
  logic [0:0] f1958_wen;
  logic [31:0] f1958_wdata;
  logic [0:0] f1958_clk;
  logic [0:0] f1958_rst;
  logic [31:0] f1958_rdata;
  sr_buffer_32_1 f1958(.wen(f1958_wen), .wdata(f1958_wdata), .clk(f1958_clk), .rst(f1958_rst), .rdata(f1958_rdata));
  assign f1958_clk = clk;
  assign f1958_rst = rst;
  // Bindings to f1958

  // f1960
  logic [0:0] f1960_wen;
  logic [31:0] f1960_wdata;
  logic [0:0] f1960_clk;
  logic [0:0] f1960_rst;
  logic [31:0] f1960_rdata;
  sr_buffer_32_1 f1960(.wen(f1960_wen), .wdata(f1960_wdata), .clk(f1960_clk), .rst(f1960_rst), .rdata(f1960_rdata));
  assign f1960_clk = clk;
  assign f1960_rst = rst;
  // Bindings to f1960

  // f1962
  logic [0:0] f1962_wen;
  logic [31:0] f1962_wdata;
  logic [0:0] f1962_clk;
  logic [0:0] f1962_rst;
  logic [31:0] f1962_rdata;
  sr_buffer_32_1 f1962(.wen(f1962_wen), .wdata(f1962_wdata), .clk(f1962_clk), .rst(f1962_rst), .rdata(f1962_rdata));
  assign f1962_clk = clk;
  assign f1962_rst = rst;
  // Bindings to f1962

  // f1964
  logic [0:0] f1964_wen;
  logic [31:0] f1964_wdata;
  logic [0:0] f1964_clk;
  logic [0:0] f1964_rst;
  logic [31:0] f1964_rdata;
  sr_buffer_32_1 f1964(.wen(f1964_wen), .wdata(f1964_wdata), .clk(f1964_clk), .rst(f1964_rst), .rdata(f1964_rdata));
  assign f1964_clk = clk;
  assign f1964_rst = rst;
  // Bindings to f1964

  // f1966
  logic [0:0] f1966_wen;
  logic [31:0] f1966_wdata;
  logic [0:0] f1966_clk;
  logic [0:0] f1966_rst;
  logic [31:0] f1966_rdata;
  sr_buffer_32_1 f1966(.wen(f1966_wen), .wdata(f1966_wdata), .clk(f1966_clk), .rst(f1966_rst), .rdata(f1966_rdata));
  assign f1966_clk = clk;
  assign f1966_rst = rst;
  // Bindings to f1966

  // f1968
  logic [0:0] f1968_wen;
  logic [31:0] f1968_wdata;
  logic [0:0] f1968_clk;
  logic [0:0] f1968_rst;
  logic [31:0] f1968_rdata;
  sr_buffer_32_1 f1968(.wen(f1968_wen), .wdata(f1968_wdata), .clk(f1968_clk), .rst(f1968_rst), .rdata(f1968_rdata));
  assign f1968_clk = clk;
  assign f1968_rst = rst;
  // Bindings to f1968

  // f1970
  logic [0:0] f1970_wen;
  logic [31:0] f1970_wdata;
  logic [0:0] f1970_clk;
  logic [0:0] f1970_rst;
  logic [31:0] f1970_rdata;
  sr_buffer_32_1 f1970(.wen(f1970_wen), .wdata(f1970_wdata), .clk(f1970_clk), .rst(f1970_rst), .rdata(f1970_rdata));
  assign f1970_clk = clk;
  assign f1970_rst = rst;
  // Bindings to f1970

  // f1972
  logic [0:0] f1972_wen;
  logic [31:0] f1972_wdata;
  logic [0:0] f1972_clk;
  logic [0:0] f1972_rst;
  logic [31:0] f1972_rdata;
  sr_buffer_32_1 f1972(.wen(f1972_wen), .wdata(f1972_wdata), .clk(f1972_clk), .rst(f1972_rst), .rdata(f1972_rdata));
  assign f1972_clk = clk;
  assign f1972_rst = rst;
  // Bindings to f1972

  // f1974
  logic [0:0] f1974_wen;
  logic [31:0] f1974_wdata;
  logic [0:0] f1974_clk;
  logic [0:0] f1974_rst;
  logic [31:0] f1974_rdata;
  sr_buffer_32_1 f1974(.wen(f1974_wen), .wdata(f1974_wdata), .clk(f1974_clk), .rst(f1974_rst), .rdata(f1974_rdata));
  assign f1974_clk = clk;
  assign f1974_rst = rst;
  // Bindings to f1974

  // f1976
  logic [0:0] f1976_wen;
  logic [31:0] f1976_wdata;
  logic [0:0] f1976_clk;
  logic [0:0] f1976_rst;
  logic [31:0] f1976_rdata;
  sr_buffer_32_1 f1976(.wen(f1976_wen), .wdata(f1976_wdata), .clk(f1976_clk), .rst(f1976_rst), .rdata(f1976_rdata));
  assign f1976_clk = clk;
  assign f1976_rst = rst;
  // Bindings to f1976

  // f1978
  logic [0:0] f1978_wen;
  logic [31:0] f1978_wdata;
  logic [0:0] f1978_clk;
  logic [0:0] f1978_rst;
  logic [31:0] f1978_rdata;
  sr_buffer_32_1 f1978(.wen(f1978_wen), .wdata(f1978_wdata), .clk(f1978_clk), .rst(f1978_rst), .rdata(f1978_rdata));
  assign f1978_clk = clk;
  assign f1978_rst = rst;
  // Bindings to f1978

  // f1980
  logic [0:0] f1980_wen;
  logic [31:0] f1980_wdata;
  logic [0:0] f1980_clk;
  logic [0:0] f1980_rst;
  logic [31:0] f1980_rdata;
  sr_buffer_32_1 f1980(.wen(f1980_wen), .wdata(f1980_wdata), .clk(f1980_clk), .rst(f1980_rst), .rdata(f1980_rdata));
  assign f1980_clk = clk;
  assign f1980_rst = rst;
  // Bindings to f1980

  // f1982
  logic [0:0] f1982_wen;
  logic [31:0] f1982_wdata;
  logic [0:0] f1982_clk;
  logic [0:0] f1982_rst;
  logic [31:0] f1982_rdata;
  sr_buffer_32_1 f1982(.wen(f1982_wen), .wdata(f1982_wdata), .clk(f1982_clk), .rst(f1982_rst), .rdata(f1982_rdata));
  assign f1982_clk = clk;
  assign f1982_rst = rst;
  // Bindings to f1982

  // f1984
  logic [0:0] f1984_wen;
  logic [31:0] f1984_wdata;
  logic [0:0] f1984_clk;
  logic [0:0] f1984_rst;
  logic [31:0] f1984_rdata;
  sr_buffer_32_1 f1984(.wen(f1984_wen), .wdata(f1984_wdata), .clk(f1984_clk), .rst(f1984_rst), .rdata(f1984_rdata));
  assign f1984_clk = clk;
  assign f1984_rst = rst;
  // Bindings to f1984

  // f1986
  logic [0:0] f1986_wen;
  logic [31:0] f1986_wdata;
  logic [0:0] f1986_clk;
  logic [0:0] f1986_rst;
  logic [31:0] f1986_rdata;
  sr_buffer_32_1 f1986(.wen(f1986_wen), .wdata(f1986_wdata), .clk(f1986_clk), .rst(f1986_rst), .rdata(f1986_rdata));
  assign f1986_clk = clk;
  assign f1986_rst = rst;
  // Bindings to f1986

  // f1988
  logic [0:0] f1988_wen;
  logic [31:0] f1988_wdata;
  logic [0:0] f1988_clk;
  logic [0:0] f1988_rst;
  logic [31:0] f1988_rdata;
  sr_buffer_32_1 f1988(.wen(f1988_wen), .wdata(f1988_wdata), .clk(f1988_clk), .rst(f1988_rst), .rdata(f1988_rdata));
  assign f1988_clk = clk;
  assign f1988_rst = rst;
  // Bindings to f1988

  // f1990
  logic [0:0] f1990_wen;
  logic [31:0] f1990_wdata;
  logic [0:0] f1990_clk;
  logic [0:0] f1990_rst;
  logic [31:0] f1990_rdata;
  sr_buffer_32_1 f1990(.wen(f1990_wen), .wdata(f1990_wdata), .clk(f1990_clk), .rst(f1990_rst), .rdata(f1990_rdata));
  assign f1990_clk = clk;
  assign f1990_rst = rst;
  // Bindings to f1990

  // f1992
  logic [0:0] f1992_wen;
  logic [31:0] f1992_wdata;
  logic [0:0] f1992_clk;
  logic [0:0] f1992_rst;
  logic [31:0] f1992_rdata;
  sr_buffer_32_1 f1992(.wen(f1992_wen), .wdata(f1992_wdata), .clk(f1992_clk), .rst(f1992_rst), .rdata(f1992_rdata));
  assign f1992_clk = clk;
  assign f1992_rst = rst;
  // Bindings to f1992

  // f1994
  logic [0:0] f1994_wen;
  logic [31:0] f1994_wdata;
  logic [0:0] f1994_clk;
  logic [0:0] f1994_rst;
  logic [31:0] f1994_rdata;
  sr_buffer_32_1 f1994(.wen(f1994_wen), .wdata(f1994_wdata), .clk(f1994_clk), .rst(f1994_rst), .rdata(f1994_rdata));
  assign f1994_clk = clk;
  assign f1994_rst = rst;
  // Bindings to f1994

  // f1996
  logic [0:0] f1996_wen;
  logic [31:0] f1996_wdata;
  logic [0:0] f1996_clk;
  logic [0:0] f1996_rst;
  logic [31:0] f1996_rdata;
  sr_buffer_32_1 f1996(.wen(f1996_wen), .wdata(f1996_wdata), .clk(f1996_clk), .rst(f1996_rst), .rdata(f1996_rdata));
  assign f1996_clk = clk;
  assign f1996_rst = rst;
  // Bindings to f1996

  // f1998
  logic [0:0] f1998_wen;
  logic [31:0] f1998_wdata;
  logic [0:0] f1998_clk;
  logic [0:0] f1998_rst;
  logic [31:0] f1998_rdata;
  sr_buffer_32_1 f1998(.wen(f1998_wen), .wdata(f1998_wdata), .clk(f1998_clk), .rst(f1998_rst), .rdata(f1998_rdata));
  assign f1998_clk = clk;
  assign f1998_rst = rst;
  // Bindings to f1998

  // f2000
  logic [0:0] f2000_wen;
  logic [31:0] f2000_wdata;
  logic [0:0] f2000_clk;
  logic [0:0] f2000_rst;
  logic [31:0] f2000_rdata;
  sr_buffer_32_1 f2000(.wen(f2000_wen), .wdata(f2000_wdata), .clk(f2000_clk), .rst(f2000_rst), .rdata(f2000_rdata));
  assign f2000_clk = clk;
  assign f2000_rst = rst;
  // Bindings to f2000

  // f2002
  logic [0:0] f2002_wen;
  logic [31:0] f2002_wdata;
  logic [0:0] f2002_clk;
  logic [0:0] f2002_rst;
  logic [31:0] f2002_rdata;
  sr_buffer_32_1 f2002(.wen(f2002_wen), .wdata(f2002_wdata), .clk(f2002_clk), .rst(f2002_rst), .rdata(f2002_rdata));
  assign f2002_clk = clk;
  assign f2002_rst = rst;
  // Bindings to f2002

  // f2004
  logic [0:0] f2004_wen;
  logic [31:0] f2004_wdata;
  logic [0:0] f2004_clk;
  logic [0:0] f2004_rst;
  logic [31:0] f2004_rdata;
  sr_buffer_32_1 f2004(.wen(f2004_wen), .wdata(f2004_wdata), .clk(f2004_clk), .rst(f2004_rst), .rdata(f2004_rdata));
  assign f2004_clk = clk;
  assign f2004_rst = rst;
  // Bindings to f2004

  // f2006
  logic [0:0] f2006_wen;
  logic [31:0] f2006_wdata;
  logic [0:0] f2006_clk;
  logic [0:0] f2006_rst;
  logic [31:0] f2006_rdata;
  sr_buffer_32_1 f2006(.wen(f2006_wen), .wdata(f2006_wdata), .clk(f2006_clk), .rst(f2006_rst), .rdata(f2006_rdata));
  assign f2006_clk = clk;
  assign f2006_rst = rst;
  // Bindings to f2006

  // f2008
  logic [0:0] f2008_wen;
  logic [31:0] f2008_wdata;
  logic [0:0] f2008_clk;
  logic [0:0] f2008_rst;
  logic [31:0] f2008_rdata;
  sr_buffer_32_1 f2008(.wen(f2008_wen), .wdata(f2008_wdata), .clk(f2008_clk), .rst(f2008_rst), .rdata(f2008_rdata));
  assign f2008_clk = clk;
  assign f2008_rst = rst;
  // Bindings to f2008

  // f2010
  logic [0:0] f2010_wen;
  logic [31:0] f2010_wdata;
  logic [0:0] f2010_clk;
  logic [0:0] f2010_rst;
  logic [31:0] f2010_rdata;
  sr_buffer_32_1 f2010(.wen(f2010_wen), .wdata(f2010_wdata), .clk(f2010_clk), .rst(f2010_rst), .rdata(f2010_rdata));
  assign f2010_clk = clk;
  assign f2010_rst = rst;
  // Bindings to f2010

  // f2012
  logic [0:0] f2012_wen;
  logic [31:0] f2012_wdata;
  logic [0:0] f2012_clk;
  logic [0:0] f2012_rst;
  logic [31:0] f2012_rdata;
  sr_buffer_32_1 f2012(.wen(f2012_wen), .wdata(f2012_wdata), .clk(f2012_clk), .rst(f2012_rst), .rdata(f2012_rdata));
  assign f2012_clk = clk;
  assign f2012_rst = rst;
  // Bindings to f2012

  // f2014
  logic [0:0] f2014_wen;
  logic [31:0] f2014_wdata;
  logic [0:0] f2014_clk;
  logic [0:0] f2014_rst;
  logic [31:0] f2014_rdata;
  sr_buffer_32_1 f2014(.wen(f2014_wen), .wdata(f2014_wdata), .clk(f2014_clk), .rst(f2014_rst), .rdata(f2014_rdata));
  assign f2014_clk = clk;
  assign f2014_rst = rst;
  // Bindings to f2014

  // f2016
  logic [0:0] f2016_wen;
  logic [31:0] f2016_wdata;
  logic [0:0] f2016_clk;
  logic [0:0] f2016_rst;
  logic [31:0] f2016_rdata;
  sr_buffer_32_1 f2016(.wen(f2016_wen), .wdata(f2016_wdata), .clk(f2016_clk), .rst(f2016_rst), .rdata(f2016_rdata));
  assign f2016_clk = clk;
  assign f2016_rst = rst;
  // Bindings to f2016

  // f2018
  logic [0:0] f2018_wen;
  logic [31:0] f2018_wdata;
  logic [0:0] f2018_clk;
  logic [0:0] f2018_rst;
  logic [31:0] f2018_rdata;
  sr_buffer_32_1 f2018(.wen(f2018_wen), .wdata(f2018_wdata), .clk(f2018_clk), .rst(f2018_rst), .rdata(f2018_rdata));
  assign f2018_clk = clk;
  assign f2018_rst = rst;
  // Bindings to f2018

  // f2020
  logic [0:0] f2020_wen;
  logic [31:0] f2020_wdata;
  logic [0:0] f2020_clk;
  logic [0:0] f2020_rst;
  logic [31:0] f2020_rdata;
  sr_buffer_32_1 f2020(.wen(f2020_wen), .wdata(f2020_wdata), .clk(f2020_clk), .rst(f2020_rst), .rdata(f2020_rdata));
  assign f2020_clk = clk;
  assign f2020_rst = rst;
  // Bindings to f2020

  // f2022
  logic [0:0] f2022_wen;
  logic [31:0] f2022_wdata;
  logic [0:0] f2022_clk;
  logic [0:0] f2022_rst;
  logic [31:0] f2022_rdata;
  sr_buffer_32_1 f2022(.wen(f2022_wen), .wdata(f2022_wdata), .clk(f2022_clk), .rst(f2022_rst), .rdata(f2022_rdata));
  assign f2022_clk = clk;
  assign f2022_rst = rst;
  // Bindings to f2022

  // f2024
  logic [0:0] f2024_wen;
  logic [31:0] f2024_wdata;
  logic [0:0] f2024_clk;
  logic [0:0] f2024_rst;
  logic [31:0] f2024_rdata;
  sr_buffer_32_1 f2024(.wen(f2024_wen), .wdata(f2024_wdata), .clk(f2024_clk), .rst(f2024_rst), .rdata(f2024_rdata));
  assign f2024_clk = clk;
  assign f2024_rst = rst;
  // Bindings to f2024

  // f2026
  logic [0:0] f2026_wen;
  logic [31:0] f2026_wdata;
  logic [0:0] f2026_clk;
  logic [0:0] f2026_rst;
  logic [31:0] f2026_rdata;
  sr_buffer_32_1 f2026(.wen(f2026_wen), .wdata(f2026_wdata), .clk(f2026_clk), .rst(f2026_rst), .rdata(f2026_rdata));
  assign f2026_clk = clk;
  assign f2026_rst = rst;
  // Bindings to f2026

  // f2028
  logic [0:0] f2028_wen;
  logic [31:0] f2028_wdata;
  logic [0:0] f2028_clk;
  logic [0:0] f2028_rst;
  logic [31:0] f2028_rdata;
  sr_buffer_32_1 f2028(.wen(f2028_wen), .wdata(f2028_wdata), .clk(f2028_clk), .rst(f2028_rst), .rdata(f2028_rdata));
  assign f2028_clk = clk;
  assign f2028_rst = rst;
  // Bindings to f2028

  // f2030
  logic [0:0] f2030_wen;
  logic [31:0] f2030_wdata;
  logic [0:0] f2030_clk;
  logic [0:0] f2030_rst;
  logic [31:0] f2030_rdata;
  sr_buffer_32_1 f2030(.wen(f2030_wen), .wdata(f2030_wdata), .clk(f2030_clk), .rst(f2030_rst), .rdata(f2030_rdata));
  assign f2030_clk = clk;
  assign f2030_rst = rst;
  // Bindings to f2030

  // f2032
  logic [0:0] f2032_wen;
  logic [31:0] f2032_wdata;
  logic [0:0] f2032_clk;
  logic [0:0] f2032_rst;
  logic [31:0] f2032_rdata;
  sr_buffer_32_1 f2032(.wen(f2032_wen), .wdata(f2032_wdata), .clk(f2032_clk), .rst(f2032_rst), .rdata(f2032_rdata));
  assign f2032_clk = clk;
  assign f2032_rst = rst;
  // Bindings to f2032

  // f2034
  logic [0:0] f2034_wen;
  logic [31:0] f2034_wdata;
  logic [0:0] f2034_clk;
  logic [0:0] f2034_rst;
  logic [31:0] f2034_rdata;
  sr_buffer_32_1 f2034(.wen(f2034_wen), .wdata(f2034_wdata), .clk(f2034_clk), .rst(f2034_rst), .rdata(f2034_rdata));
  assign f2034_clk = clk;
  assign f2034_rst = rst;
  // Bindings to f2034

  // f2036
  logic [0:0] f2036_wen;
  logic [31:0] f2036_wdata;
  logic [0:0] f2036_clk;
  logic [0:0] f2036_rst;
  logic [31:0] f2036_rdata;
  sr_buffer_32_1 f2036(.wen(f2036_wen), .wdata(f2036_wdata), .clk(f2036_clk), .rst(f2036_rst), .rdata(f2036_rdata));
  assign f2036_clk = clk;
  assign f2036_rst = rst;
  // Bindings to f2036

  // f2038
  logic [0:0] f2038_wen;
  logic [31:0] f2038_wdata;
  logic [0:0] f2038_clk;
  logic [0:0] f2038_rst;
  logic [31:0] f2038_rdata;
  sr_buffer_32_1 f2038(.wen(f2038_wen), .wdata(f2038_wdata), .clk(f2038_clk), .rst(f2038_rst), .rdata(f2038_rdata));
  assign f2038_clk = clk;
  assign f2038_rst = rst;
  // Bindings to f2038

  // f2040
  logic [0:0] f2040_wen;
  logic [31:0] f2040_wdata;
  logic [0:0] f2040_clk;
  logic [0:0] f2040_rst;
  logic [31:0] f2040_rdata;
  sr_buffer_32_1 f2040(.wen(f2040_wen), .wdata(f2040_wdata), .clk(f2040_clk), .rst(f2040_rst), .rdata(f2040_rdata));
  assign f2040_clk = clk;
  assign f2040_rst = rst;
  // Bindings to f2040

  // f2042
  logic [0:0] f2042_wen;
  logic [31:0] f2042_wdata;
  logic [0:0] f2042_clk;
  logic [0:0] f2042_rst;
  logic [31:0] f2042_rdata;
  sr_buffer_32_1 f2042(.wen(f2042_wen), .wdata(f2042_wdata), .clk(f2042_clk), .rst(f2042_rst), .rdata(f2042_rdata));
  assign f2042_clk = clk;
  assign f2042_rst = rst;
  // Bindings to f2042

  // f2044
  logic [0:0] f2044_wen;
  logic [31:0] f2044_wdata;
  logic [0:0] f2044_clk;
  logic [0:0] f2044_rst;
  logic [31:0] f2044_rdata;
  sr_buffer_32_1 f2044(.wen(f2044_wen), .wdata(f2044_wdata), .clk(f2044_clk), .rst(f2044_rst), .rdata(f2044_rdata));
  assign f2044_clk = clk;
  assign f2044_rst = rst;
  // Bindings to f2044

  // f2046
  logic [0:0] f2046_wen;
  logic [31:0] f2046_wdata;
  logic [0:0] f2046_clk;
  logic [0:0] f2046_rst;
  logic [31:0] f2046_rdata;
  sr_buffer_32_1 f2046(.wen(f2046_wen), .wdata(f2046_wdata), .clk(f2046_clk), .rst(f2046_rst), .rdata(f2046_rdata));
  assign f2046_clk = clk;
  assign f2046_rst = rst;
  // Bindings to f2046

  // f2048
  logic [0:0] f2048_wen;
  logic [31:0] f2048_wdata;
  logic [0:0] f2048_clk;
  logic [0:0] f2048_rst;
  logic [31:0] f2048_rdata;
  sr_buffer_32_1 f2048(.wen(f2048_wen), .wdata(f2048_wdata), .clk(f2048_clk), .rst(f2048_rst), .rdata(f2048_rdata));
  assign f2048_clk = clk;
  assign f2048_rst = rst;
  // Bindings to f2048

  // f2050
  logic [0:0] f2050_wen;
  logic [31:0] f2050_wdata;
  logic [0:0] f2050_clk;
  logic [0:0] f2050_rst;
  logic [31:0] f2050_rdata;
  sr_buffer_32_1 f2050(.wen(f2050_wen), .wdata(f2050_wdata), .clk(f2050_clk), .rst(f2050_rst), .rdata(f2050_rdata));
  assign f2050_clk = clk;
  assign f2050_rst = rst;
  // Bindings to f2050

  // f2052
  logic [0:0] f2052_wen;
  logic [31:0] f2052_wdata;
  logic [0:0] f2052_clk;
  logic [0:0] f2052_rst;
  logic [31:0] f2052_rdata;
  sr_buffer_32_1 f2052(.wen(f2052_wen), .wdata(f2052_wdata), .clk(f2052_clk), .rst(f2052_rst), .rdata(f2052_rdata));
  assign f2052_clk = clk;
  assign f2052_rst = rst;
  // Bindings to f2052

  // f2054
  logic [0:0] f2054_wen;
  logic [31:0] f2054_wdata;
  logic [0:0] f2054_clk;
  logic [0:0] f2054_rst;
  logic [31:0] f2054_rdata;
  sr_buffer_32_1 f2054(.wen(f2054_wen), .wdata(f2054_wdata), .clk(f2054_clk), .rst(f2054_rst), .rdata(f2054_rdata));
  assign f2054_clk = clk;
  assign f2054_rst = rst;
  // Bindings to f2054

  // f2056
  logic [0:0] f2056_wen;
  logic [31:0] f2056_wdata;
  logic [0:0] f2056_clk;
  logic [0:0] f2056_rst;
  logic [31:0] f2056_rdata;
  sr_buffer_32_1 f2056(.wen(f2056_wen), .wdata(f2056_wdata), .clk(f2056_clk), .rst(f2056_rst), .rdata(f2056_rdata));
  assign f2056_clk = clk;
  assign f2056_rst = rst;
  // Bindings to f2056

  // f2058
  logic [0:0] f2058_wen;
  logic [31:0] f2058_wdata;
  logic [0:0] f2058_clk;
  logic [0:0] f2058_rst;
  logic [31:0] f2058_rdata;
  sr_buffer_32_1 f2058(.wen(f2058_wen), .wdata(f2058_wdata), .clk(f2058_clk), .rst(f2058_rst), .rdata(f2058_rdata));
  assign f2058_clk = clk;
  assign f2058_rst = rst;
  // Bindings to f2058

  // f2060
  logic [0:0] f2060_wen;
  logic [31:0] f2060_wdata;
  logic [0:0] f2060_clk;
  logic [0:0] f2060_rst;
  logic [31:0] f2060_rdata;
  sr_buffer_32_1 f2060(.wen(f2060_wen), .wdata(f2060_wdata), .clk(f2060_clk), .rst(f2060_rst), .rdata(f2060_rdata));
  assign f2060_clk = clk;
  assign f2060_rst = rst;
  // Bindings to f2060

  // f2062
  logic [0:0] f2062_wen;
  logic [31:0] f2062_wdata;
  logic [0:0] f2062_clk;
  logic [0:0] f2062_rst;
  logic [31:0] f2062_rdata;
  sr_buffer_32_1 f2062(.wen(f2062_wen), .wdata(f2062_wdata), .clk(f2062_clk), .rst(f2062_rst), .rdata(f2062_rdata));
  assign f2062_clk = clk;
  assign f2062_rst = rst;
  // Bindings to f2062

  // f2064
  logic [0:0] f2064_wen;
  logic [31:0] f2064_wdata;
  logic [0:0] f2064_clk;
  logic [0:0] f2064_rst;
  logic [31:0] f2064_rdata;
  sr_buffer_32_1 f2064(.wen(f2064_wen), .wdata(f2064_wdata), .clk(f2064_clk), .rst(f2064_rst), .rdata(f2064_rdata));
  assign f2064_clk = clk;
  assign f2064_rst = rst;
  // Bindings to f2064

  // f2066
  logic [0:0] f2066_wen;
  logic [31:0] f2066_wdata;
  logic [0:0] f2066_clk;
  logic [0:0] f2066_rst;
  logic [31:0] f2066_rdata;
  sr_buffer_32_1 f2066(.wen(f2066_wen), .wdata(f2066_wdata), .clk(f2066_clk), .rst(f2066_rst), .rdata(f2066_rdata));
  assign f2066_clk = clk;
  assign f2066_rst = rst;
  // Bindings to f2066

  // f2068
  logic [0:0] f2068_wen;
  logic [31:0] f2068_wdata;
  logic [0:0] f2068_clk;
  logic [0:0] f2068_rst;
  logic [31:0] f2068_rdata;
  sr_buffer_32_1 f2068(.wen(f2068_wen), .wdata(f2068_wdata), .clk(f2068_clk), .rst(f2068_rst), .rdata(f2068_rdata));
  assign f2068_clk = clk;
  assign f2068_rst = rst;
  // Bindings to f2068

  // f2070
  logic [0:0] f2070_wen;
  logic [31:0] f2070_wdata;
  logic [0:0] f2070_clk;
  logic [0:0] f2070_rst;
  logic [31:0] f2070_rdata;
  sr_buffer_32_1 f2070(.wen(f2070_wen), .wdata(f2070_wdata), .clk(f2070_clk), .rst(f2070_rst), .rdata(f2070_rdata));
  assign f2070_clk = clk;
  assign f2070_rst = rst;
  // Bindings to f2070

  // f2072
  logic [0:0] f2072_wen;
  logic [31:0] f2072_wdata;
  logic [0:0] f2072_clk;
  logic [0:0] f2072_rst;
  logic [31:0] f2072_rdata;
  sr_buffer_32_1 f2072(.wen(f2072_wen), .wdata(f2072_wdata), .clk(f2072_clk), .rst(f2072_rst), .rdata(f2072_rdata));
  assign f2072_clk = clk;
  assign f2072_rst = rst;
  // Bindings to f2072

  // f2074
  logic [0:0] f2074_wen;
  logic [31:0] f2074_wdata;
  logic [0:0] f2074_clk;
  logic [0:0] f2074_rst;
  logic [31:0] f2074_rdata;
  sr_buffer_32_1 f2074(.wen(f2074_wen), .wdata(f2074_wdata), .clk(f2074_clk), .rst(f2074_rst), .rdata(f2074_rdata));
  assign f2074_clk = clk;
  assign f2074_rst = rst;
  // Bindings to f2074

  // f2076
  logic [0:0] f2076_wen;
  logic [31:0] f2076_wdata;
  logic [0:0] f2076_clk;
  logic [0:0] f2076_rst;
  logic [31:0] f2076_rdata;
  sr_buffer_32_1 f2076(.wen(f2076_wen), .wdata(f2076_wdata), .clk(f2076_clk), .rst(f2076_rst), .rdata(f2076_rdata));
  assign f2076_clk = clk;
  assign f2076_rst = rst;
  // Bindings to f2076

  // f2078
  logic [0:0] f2078_wen;
  logic [31:0] f2078_wdata;
  logic [0:0] f2078_clk;
  logic [0:0] f2078_rst;
  logic [31:0] f2078_rdata;
  sr_buffer_32_1 f2078(.wen(f2078_wen), .wdata(f2078_wdata), .clk(f2078_clk), .rst(f2078_rst), .rdata(f2078_rdata));
  assign f2078_clk = clk;
  assign f2078_rst = rst;
  // Bindings to f2078

  // f2080
  logic [0:0] f2080_wen;
  logic [31:0] f2080_wdata;
  logic [0:0] f2080_clk;
  logic [0:0] f2080_rst;
  logic [31:0] f2080_rdata;
  sr_buffer_32_1 f2080(.wen(f2080_wen), .wdata(f2080_wdata), .clk(f2080_clk), .rst(f2080_rst), .rdata(f2080_rdata));
  assign f2080_clk = clk;
  assign f2080_rst = rst;
  // Bindings to f2080

  // f2082
  logic [0:0] f2082_wen;
  logic [31:0] f2082_wdata;
  logic [0:0] f2082_clk;
  logic [0:0] f2082_rst;
  logic [31:0] f2082_rdata;
  sr_buffer_32_1 f2082(.wen(f2082_wen), .wdata(f2082_wdata), .clk(f2082_clk), .rst(f2082_rst), .rdata(f2082_rdata));
  assign f2082_clk = clk;
  assign f2082_rst = rst;
  // Bindings to f2082

  // f2084
  logic [0:0] f2084_wen;
  logic [31:0] f2084_wdata;
  logic [0:0] f2084_clk;
  logic [0:0] f2084_rst;
  logic [31:0] f2084_rdata;
  sr_buffer_32_1 f2084(.wen(f2084_wen), .wdata(f2084_wdata), .clk(f2084_clk), .rst(f2084_rst), .rdata(f2084_rdata));
  assign f2084_clk = clk;
  assign f2084_rst = rst;
  // Bindings to f2084

  // f2086
  logic [0:0] f2086_wen;
  logic [31:0] f2086_wdata;
  logic [0:0] f2086_clk;
  logic [0:0] f2086_rst;
  logic [31:0] f2086_rdata;
  sr_buffer_32_1 f2086(.wen(f2086_wen), .wdata(f2086_wdata), .clk(f2086_clk), .rst(f2086_rst), .rdata(f2086_rdata));
  assign f2086_clk = clk;
  assign f2086_rst = rst;
  // Bindings to f2086

  // f2088
  logic [0:0] f2088_wen;
  logic [31:0] f2088_wdata;
  logic [0:0] f2088_clk;
  logic [0:0] f2088_rst;
  logic [31:0] f2088_rdata;
  sr_buffer_32_1 f2088(.wen(f2088_wen), .wdata(f2088_wdata), .clk(f2088_clk), .rst(f2088_rst), .rdata(f2088_rdata));
  assign f2088_clk = clk;
  assign f2088_rst = rst;
  // Bindings to f2088

  // f2090
  logic [0:0] f2090_wen;
  logic [31:0] f2090_wdata;
  logic [0:0] f2090_clk;
  logic [0:0] f2090_rst;
  logic [31:0] f2090_rdata;
  sr_buffer_32_1 f2090(.wen(f2090_wen), .wdata(f2090_wdata), .clk(f2090_clk), .rst(f2090_rst), .rdata(f2090_rdata));
  assign f2090_clk = clk;
  assign f2090_rst = rst;
  // Bindings to f2090

  // f2092
  logic [0:0] f2092_wen;
  logic [31:0] f2092_wdata;
  logic [0:0] f2092_clk;
  logic [0:0] f2092_rst;
  logic [31:0] f2092_rdata;
  sr_buffer_32_1 f2092(.wen(f2092_wen), .wdata(f2092_wdata), .clk(f2092_clk), .rst(f2092_rst), .rdata(f2092_rdata));
  assign f2092_clk = clk;
  assign f2092_rst = rst;
  // Bindings to f2092

  // f2094
  logic [0:0] f2094_wen;
  logic [31:0] f2094_wdata;
  logic [0:0] f2094_clk;
  logic [0:0] f2094_rst;
  logic [31:0] f2094_rdata;
  sr_buffer_32_1 f2094(.wen(f2094_wen), .wdata(f2094_wdata), .clk(f2094_clk), .rst(f2094_rst), .rdata(f2094_rdata));
  assign f2094_clk = clk;
  assign f2094_rst = rst;
  // Bindings to f2094

  // f2096
  logic [0:0] f2096_wen;
  logic [31:0] f2096_wdata;
  logic [0:0] f2096_clk;
  logic [0:0] f2096_rst;
  logic [31:0] f2096_rdata;
  sr_buffer_32_1 f2096(.wen(f2096_wen), .wdata(f2096_wdata), .clk(f2096_clk), .rst(f2096_rst), .rdata(f2096_rdata));
  assign f2096_clk = clk;
  assign f2096_rst = rst;
  // Bindings to f2096

  // f2098
  logic [0:0] f2098_wen;
  logic [31:0] f2098_wdata;
  logic [0:0] f2098_clk;
  logic [0:0] f2098_rst;
  logic [31:0] f2098_rdata;
  sr_buffer_32_1 f2098(.wen(f2098_wen), .wdata(f2098_wdata), .clk(f2098_clk), .rst(f2098_rst), .rdata(f2098_rdata));
  assign f2098_clk = clk;
  assign f2098_rst = rst;
  // Bindings to f2098

  // f2100
  logic [0:0] f2100_wen;
  logic [31:0] f2100_wdata;
  logic [0:0] f2100_clk;
  logic [0:0] f2100_rst;
  logic [31:0] f2100_rdata;
  sr_buffer_32_1 f2100(.wen(f2100_wen), .wdata(f2100_wdata), .clk(f2100_clk), .rst(f2100_rst), .rdata(f2100_rdata));
  assign f2100_clk = clk;
  assign f2100_rst = rst;
  // Bindings to f2100

  // f2102
  logic [0:0] f2102_wen;
  logic [31:0] f2102_wdata;
  logic [0:0] f2102_clk;
  logic [0:0] f2102_rst;
  logic [31:0] f2102_rdata;
  sr_buffer_32_1 f2102(.wen(f2102_wen), .wdata(f2102_wdata), .clk(f2102_clk), .rst(f2102_rst), .rdata(f2102_rdata));
  assign f2102_clk = clk;
  assign f2102_rst = rst;
  // Bindings to f2102

  // f2104
  logic [0:0] f2104_wen;
  logic [31:0] f2104_wdata;
  logic [0:0] f2104_clk;
  logic [0:0] f2104_rst;
  logic [31:0] f2104_rdata;
  sr_buffer_32_1 f2104(.wen(f2104_wen), .wdata(f2104_wdata), .clk(f2104_clk), .rst(f2104_rst), .rdata(f2104_rdata));
  assign f2104_clk = clk;
  assign f2104_rst = rst;
  // Bindings to f2104

  // f2106
  logic [0:0] f2106_wen;
  logic [31:0] f2106_wdata;
  logic [0:0] f2106_clk;
  logic [0:0] f2106_rst;
  logic [31:0] f2106_rdata;
  sr_buffer_32_1 f2106(.wen(f2106_wen), .wdata(f2106_wdata), .clk(f2106_clk), .rst(f2106_rst), .rdata(f2106_rdata));
  assign f2106_clk = clk;
  assign f2106_rst = rst;
  // Bindings to f2106

  // f2108
  logic [0:0] f2108_wen;
  logic [31:0] f2108_wdata;
  logic [0:0] f2108_clk;
  logic [0:0] f2108_rst;
  logic [31:0] f2108_rdata;
  sr_buffer_32_1 f2108(.wen(f2108_wen), .wdata(f2108_wdata), .clk(f2108_clk), .rst(f2108_rst), .rdata(f2108_rdata));
  assign f2108_clk = clk;
  assign f2108_rst = rst;
  // Bindings to f2108

  // f2110
  logic [0:0] f2110_wen;
  logic [31:0] f2110_wdata;
  logic [0:0] f2110_clk;
  logic [0:0] f2110_rst;
  logic [31:0] f2110_rdata;
  sr_buffer_32_1 f2110(.wen(f2110_wen), .wdata(f2110_wdata), .clk(f2110_clk), .rst(f2110_rst), .rdata(f2110_rdata));
  assign f2110_clk = clk;
  assign f2110_rst = rst;
  // Bindings to f2110

  // f2112
  logic [0:0] f2112_wen;
  logic [31:0] f2112_wdata;
  logic [0:0] f2112_clk;
  logic [0:0] f2112_rst;
  logic [31:0] f2112_rdata;
  sr_buffer_32_1 f2112(.wen(f2112_wen), .wdata(f2112_wdata), .clk(f2112_clk), .rst(f2112_rst), .rdata(f2112_rdata));
  assign f2112_clk = clk;
  assign f2112_rst = rst;
  // Bindings to f2112

  // f2114
  logic [0:0] f2114_wen;
  logic [31:0] f2114_wdata;
  logic [0:0] f2114_clk;
  logic [0:0] f2114_rst;
  logic [31:0] f2114_rdata;
  sr_buffer_32_1 f2114(.wen(f2114_wen), .wdata(f2114_wdata), .clk(f2114_clk), .rst(f2114_rst), .rdata(f2114_rdata));
  assign f2114_clk = clk;
  assign f2114_rst = rst;
  // Bindings to f2114

  // f2116
  logic [0:0] f2116_wen;
  logic [31:0] f2116_wdata;
  logic [0:0] f2116_clk;
  logic [0:0] f2116_rst;
  logic [31:0] f2116_rdata;
  sr_buffer_32_1 f2116(.wen(f2116_wen), .wdata(f2116_wdata), .clk(f2116_clk), .rst(f2116_rst), .rdata(f2116_rdata));
  assign f2116_clk = clk;
  assign f2116_rst = rst;
  // Bindings to f2116

  // f2118
  logic [0:0] f2118_wen;
  logic [31:0] f2118_wdata;
  logic [0:0] f2118_clk;
  logic [0:0] f2118_rst;
  logic [31:0] f2118_rdata;
  sr_buffer_32_1 f2118(.wen(f2118_wen), .wdata(f2118_wdata), .clk(f2118_clk), .rst(f2118_rst), .rdata(f2118_rdata));
  assign f2118_clk = clk;
  assign f2118_rst = rst;
  // Bindings to f2118

  // f2120
  logic [0:0] f2120_wen;
  logic [31:0] f2120_wdata;
  logic [0:0] f2120_clk;
  logic [0:0] f2120_rst;
  logic [31:0] f2120_rdata;
  sr_buffer_32_1 f2120(.wen(f2120_wen), .wdata(f2120_wdata), .clk(f2120_clk), .rst(f2120_rst), .rdata(f2120_rdata));
  assign f2120_clk = clk;
  assign f2120_rst = rst;
  // Bindings to f2120

  // f2122
  logic [0:0] f2122_wen;
  logic [31:0] f2122_wdata;
  logic [0:0] f2122_clk;
  logic [0:0] f2122_rst;
  logic [31:0] f2122_rdata;
  sr_buffer_32_1 f2122(.wen(f2122_wen), .wdata(f2122_wdata), .clk(f2122_clk), .rst(f2122_rst), .rdata(f2122_rdata));
  assign f2122_clk = clk;
  assign f2122_rst = rst;
  // Bindings to f2122

  // f2124
  logic [0:0] f2124_wen;
  logic [31:0] f2124_wdata;
  logic [0:0] f2124_clk;
  logic [0:0] f2124_rst;
  logic [31:0] f2124_rdata;
  sr_buffer_32_1 f2124(.wen(f2124_wen), .wdata(f2124_wdata), .clk(f2124_clk), .rst(f2124_rst), .rdata(f2124_rdata));
  assign f2124_clk = clk;
  assign f2124_rst = rst;
  // Bindings to f2124

  // f2126
  logic [0:0] f2126_wen;
  logic [31:0] f2126_wdata;
  logic [0:0] f2126_clk;
  logic [0:0] f2126_rst;
  logic [31:0] f2126_rdata;
  sr_buffer_32_1 f2126(.wen(f2126_wen), .wdata(f2126_wdata), .clk(f2126_clk), .rst(f2126_rst), .rdata(f2126_rdata));
  assign f2126_clk = clk;
  assign f2126_rst = rst;
  // Bindings to f2126

  // f2128
  logic [0:0] f2128_wen;
  logic [31:0] f2128_wdata;
  logic [0:0] f2128_clk;
  logic [0:0] f2128_rst;
  logic [31:0] f2128_rdata;
  sr_buffer_32_1 f2128(.wen(f2128_wen), .wdata(f2128_wdata), .clk(f2128_clk), .rst(f2128_rst), .rdata(f2128_rdata));
  assign f2128_clk = clk;
  assign f2128_rst = rst;
  // Bindings to f2128

  // f2130
  logic [0:0] f2130_wen;
  logic [31:0] f2130_wdata;
  logic [0:0] f2130_clk;
  logic [0:0] f2130_rst;
  logic [31:0] f2130_rdata;
  sr_buffer_32_1 f2130(.wen(f2130_wen), .wdata(f2130_wdata), .clk(f2130_clk), .rst(f2130_rst), .rdata(f2130_rdata));
  assign f2130_clk = clk;
  assign f2130_rst = rst;
  // Bindings to f2130

  // f2132
  logic [0:0] f2132_wen;
  logic [31:0] f2132_wdata;
  logic [0:0] f2132_clk;
  logic [0:0] f2132_rst;
  logic [31:0] f2132_rdata;
  sr_buffer_32_1 f2132(.wen(f2132_wen), .wdata(f2132_wdata), .clk(f2132_clk), .rst(f2132_rst), .rdata(f2132_rdata));
  assign f2132_clk = clk;
  assign f2132_rst = rst;
  // Bindings to f2132

  // f2134
  logic [0:0] f2134_wen;
  logic [31:0] f2134_wdata;
  logic [0:0] f2134_clk;
  logic [0:0] f2134_rst;
  logic [31:0] f2134_rdata;
  sr_buffer_32_1 f2134(.wen(f2134_wen), .wdata(f2134_wdata), .clk(f2134_clk), .rst(f2134_rst), .rdata(f2134_rdata));
  assign f2134_clk = clk;
  assign f2134_rst = rst;
  // Bindings to f2134

  // f2136
  logic [0:0] f2136_wen;
  logic [31:0] f2136_wdata;
  logic [0:0] f2136_clk;
  logic [0:0] f2136_rst;
  logic [31:0] f2136_rdata;
  sr_buffer_32_1 f2136(.wen(f2136_wen), .wdata(f2136_wdata), .clk(f2136_clk), .rst(f2136_rst), .rdata(f2136_rdata));
  assign f2136_clk = clk;
  assign f2136_rst = rst;
  // Bindings to f2136

  // f2138
  logic [0:0] f2138_wen;
  logic [31:0] f2138_wdata;
  logic [0:0] f2138_clk;
  logic [0:0] f2138_rst;
  logic [31:0] f2138_rdata;
  sr_buffer_32_1 f2138(.wen(f2138_wen), .wdata(f2138_wdata), .clk(f2138_clk), .rst(f2138_rst), .rdata(f2138_rdata));
  assign f2138_clk = clk;
  assign f2138_rst = rst;
  // Bindings to f2138

  // f2140
  logic [0:0] f2140_wen;
  logic [31:0] f2140_wdata;
  logic [0:0] f2140_clk;
  logic [0:0] f2140_rst;
  logic [31:0] f2140_rdata;
  sr_buffer_32_1 f2140(.wen(f2140_wen), .wdata(f2140_wdata), .clk(f2140_clk), .rst(f2140_rst), .rdata(f2140_rdata));
  assign f2140_clk = clk;
  assign f2140_rst = rst;
  // Bindings to f2140

  // f2142
  logic [0:0] f2142_wen;
  logic [31:0] f2142_wdata;
  logic [0:0] f2142_clk;
  logic [0:0] f2142_rst;
  logic [31:0] f2142_rdata;
  sr_buffer_32_1 f2142(.wen(f2142_wen), .wdata(f2142_wdata), .clk(f2142_clk), .rst(f2142_rst), .rdata(f2142_rdata));
  assign f2142_clk = clk;
  assign f2142_rst = rst;
  // Bindings to f2142

  // f2144
  logic [0:0] f2144_wen;
  logic [31:0] f2144_wdata;
  logic [0:0] f2144_clk;
  logic [0:0] f2144_rst;
  logic [31:0] f2144_rdata;
  sr_buffer_32_1 f2144(.wen(f2144_wen), .wdata(f2144_wdata), .clk(f2144_clk), .rst(f2144_rst), .rdata(f2144_rdata));
  assign f2144_clk = clk;
  assign f2144_rst = rst;
  // Bindings to f2144

  // f2146
  logic [0:0] f2146_wen;
  logic [31:0] f2146_wdata;
  logic [0:0] f2146_clk;
  logic [0:0] f2146_rst;
  logic [31:0] f2146_rdata;
  sr_buffer_32_1 f2146(.wen(f2146_wen), .wdata(f2146_wdata), .clk(f2146_clk), .rst(f2146_rst), .rdata(f2146_rdata));
  assign f2146_clk = clk;
  assign f2146_rst = rst;
  // Bindings to f2146

  // f2148
  logic [0:0] f2148_wen;
  logic [31:0] f2148_wdata;
  logic [0:0] f2148_clk;
  logic [0:0] f2148_rst;
  logic [31:0] f2148_rdata;
  sr_buffer_32_1 f2148(.wen(f2148_wen), .wdata(f2148_wdata), .clk(f2148_clk), .rst(f2148_rst), .rdata(f2148_rdata));
  assign f2148_clk = clk;
  assign f2148_rst = rst;
  // Bindings to f2148

  // f2150
  logic [0:0] f2150_wen;
  logic [31:0] f2150_wdata;
  logic [0:0] f2150_clk;
  logic [0:0] f2150_rst;
  logic [31:0] f2150_rdata;
  sr_buffer_32_1 f2150(.wen(f2150_wen), .wdata(f2150_wdata), .clk(f2150_clk), .rst(f2150_rst), .rdata(f2150_rdata));
  assign f2150_clk = clk;
  assign f2150_rst = rst;
  // Bindings to f2150

  // f2152
  logic [0:0] f2152_wen;
  logic [31:0] f2152_wdata;
  logic [0:0] f2152_clk;
  logic [0:0] f2152_rst;
  logic [31:0] f2152_rdata;
  sr_buffer_32_1 f2152(.wen(f2152_wen), .wdata(f2152_wdata), .clk(f2152_clk), .rst(f2152_rst), .rdata(f2152_rdata));
  assign f2152_clk = clk;
  assign f2152_rst = rst;
  // Bindings to f2152

  // f2154
  logic [0:0] f2154_wen;
  logic [31:0] f2154_wdata;
  logic [0:0] f2154_clk;
  logic [0:0] f2154_rst;
  logic [31:0] f2154_rdata;
  sr_buffer_32_1 f2154(.wen(f2154_wen), .wdata(f2154_wdata), .clk(f2154_clk), .rst(f2154_rst), .rdata(f2154_rdata));
  assign f2154_clk = clk;
  assign f2154_rst = rst;
  // Bindings to f2154

  // f2156
  logic [0:0] f2156_wen;
  logic [31:0] f2156_wdata;
  logic [0:0] f2156_clk;
  logic [0:0] f2156_rst;
  logic [31:0] f2156_rdata;
  sr_buffer_32_1 f2156(.wen(f2156_wen), .wdata(f2156_wdata), .clk(f2156_clk), .rst(f2156_rst), .rdata(f2156_rdata));
  assign f2156_clk = clk;
  assign f2156_rst = rst;
  // Bindings to f2156

  // f2158
  logic [0:0] f2158_wen;
  logic [31:0] f2158_wdata;
  logic [0:0] f2158_clk;
  logic [0:0] f2158_rst;
  logic [31:0] f2158_rdata;
  sr_buffer_32_1 f2158(.wen(f2158_wen), .wdata(f2158_wdata), .clk(f2158_clk), .rst(f2158_rst), .rdata(f2158_rdata));
  assign f2158_clk = clk;
  assign f2158_rst = rst;
  // Bindings to f2158

  // f2160
  logic [0:0] f2160_wen;
  logic [31:0] f2160_wdata;
  logic [0:0] f2160_clk;
  logic [0:0] f2160_rst;
  logic [31:0] f2160_rdata;
  sr_buffer_32_1 f2160(.wen(f2160_wen), .wdata(f2160_wdata), .clk(f2160_clk), .rst(f2160_rst), .rdata(f2160_rdata));
  assign f2160_clk = clk;
  assign f2160_rst = rst;
  // Bindings to f2160

  // f2162
  logic [0:0] f2162_wen;
  logic [31:0] f2162_wdata;
  logic [0:0] f2162_clk;
  logic [0:0] f2162_rst;
  logic [31:0] f2162_rdata;
  sr_buffer_32_1 f2162(.wen(f2162_wen), .wdata(f2162_wdata), .clk(f2162_clk), .rst(f2162_rst), .rdata(f2162_rdata));
  assign f2162_clk = clk;
  assign f2162_rst = rst;
  // Bindings to f2162

  // f2164
  logic [0:0] f2164_wen;
  logic [31:0] f2164_wdata;
  logic [0:0] f2164_clk;
  logic [0:0] f2164_rst;
  logic [31:0] f2164_rdata;
  sr_buffer_32_1 f2164(.wen(f2164_wen), .wdata(f2164_wdata), .clk(f2164_clk), .rst(f2164_rst), .rdata(f2164_rdata));
  assign f2164_clk = clk;
  assign f2164_rst = rst;
  // Bindings to f2164

  // f2166
  logic [0:0] f2166_wen;
  logic [31:0] f2166_wdata;
  logic [0:0] f2166_clk;
  logic [0:0] f2166_rst;
  logic [31:0] f2166_rdata;
  sr_buffer_32_1 f2166(.wen(f2166_wen), .wdata(f2166_wdata), .clk(f2166_clk), .rst(f2166_rst), .rdata(f2166_rdata));
  assign f2166_clk = clk;
  assign f2166_rst = rst;
  // Bindings to f2166

  // f2168
  logic [0:0] f2168_wen;
  logic [31:0] f2168_wdata;
  logic [0:0] f2168_clk;
  logic [0:0] f2168_rst;
  logic [31:0] f2168_rdata;
  sr_buffer_32_1 f2168(.wen(f2168_wen), .wdata(f2168_wdata), .clk(f2168_clk), .rst(f2168_rst), .rdata(f2168_rdata));
  assign f2168_clk = clk;
  assign f2168_rst = rst;
  // Bindings to f2168

  // f2170
  logic [0:0] f2170_wen;
  logic [31:0] f2170_wdata;
  logic [0:0] f2170_clk;
  logic [0:0] f2170_rst;
  logic [31:0] f2170_rdata;
  sr_buffer_32_1 f2170(.wen(f2170_wen), .wdata(f2170_wdata), .clk(f2170_clk), .rst(f2170_rst), .rdata(f2170_rdata));
  assign f2170_clk = clk;
  assign f2170_rst = rst;
  // Bindings to f2170

  // f2172
  logic [0:0] f2172_wen;
  logic [31:0] f2172_wdata;
  logic [0:0] f2172_clk;
  logic [0:0] f2172_rst;
  logic [31:0] f2172_rdata;
  sr_buffer_32_1 f2172(.wen(f2172_wen), .wdata(f2172_wdata), .clk(f2172_clk), .rst(f2172_rst), .rdata(f2172_rdata));
  assign f2172_clk = clk;
  assign f2172_rst = rst;
  // Bindings to f2172

  // f2174
  logic [0:0] f2174_wen;
  logic [31:0] f2174_wdata;
  logic [0:0] f2174_clk;
  logic [0:0] f2174_rst;
  logic [31:0] f2174_rdata;
  sr_buffer_32_1 f2174(.wen(f2174_wen), .wdata(f2174_wdata), .clk(f2174_clk), .rst(f2174_rst), .rdata(f2174_rdata));
  assign f2174_clk = clk;
  assign f2174_rst = rst;
  // Bindings to f2174

  // f2176
  logic [0:0] f2176_wen;
  logic [31:0] f2176_wdata;
  logic [0:0] f2176_clk;
  logic [0:0] f2176_rst;
  logic [31:0] f2176_rdata;
  sr_buffer_32_1 f2176(.wen(f2176_wen), .wdata(f2176_wdata), .clk(f2176_clk), .rst(f2176_rst), .rdata(f2176_rdata));
  assign f2176_clk = clk;
  assign f2176_rst = rst;
  // Bindings to f2176

  // f2178
  logic [0:0] f2178_wen;
  logic [31:0] f2178_wdata;
  logic [0:0] f2178_clk;
  logic [0:0] f2178_rst;
  logic [31:0] f2178_rdata;
  sr_buffer_32_1 f2178(.wen(f2178_wen), .wdata(f2178_wdata), .clk(f2178_clk), .rst(f2178_rst), .rdata(f2178_rdata));
  assign f2178_clk = clk;
  assign f2178_rst = rst;
  // Bindings to f2178

  // f2180
  logic [0:0] f2180_wen;
  logic [31:0] f2180_wdata;
  logic [0:0] f2180_clk;
  logic [0:0] f2180_rst;
  logic [31:0] f2180_rdata;
  sr_buffer_32_1 f2180(.wen(f2180_wen), .wdata(f2180_wdata), .clk(f2180_clk), .rst(f2180_rst), .rdata(f2180_rdata));
  assign f2180_clk = clk;
  assign f2180_rst = rst;
  // Bindings to f2180

  // f2182
  logic [0:0] f2182_wen;
  logic [31:0] f2182_wdata;
  logic [0:0] f2182_clk;
  logic [0:0] f2182_rst;
  logic [31:0] f2182_rdata;
  sr_buffer_32_1 f2182(.wen(f2182_wen), .wdata(f2182_wdata), .clk(f2182_clk), .rst(f2182_rst), .rdata(f2182_rdata));
  assign f2182_clk = clk;
  assign f2182_rst = rst;
  // Bindings to f2182

  // f2184
  logic [0:0] f2184_wen;
  logic [31:0] f2184_wdata;
  logic [0:0] f2184_clk;
  logic [0:0] f2184_rst;
  logic [31:0] f2184_rdata;
  sr_buffer_32_1 f2184(.wen(f2184_wen), .wdata(f2184_wdata), .clk(f2184_clk), .rst(f2184_rst), .rdata(f2184_rdata));
  assign f2184_clk = clk;
  assign f2184_rst = rst;
  // Bindings to f2184

  // f2186
  logic [0:0] f2186_wen;
  logic [31:0] f2186_wdata;
  logic [0:0] f2186_clk;
  logic [0:0] f2186_rst;
  logic [31:0] f2186_rdata;
  sr_buffer_32_1 f2186(.wen(f2186_wen), .wdata(f2186_wdata), .clk(f2186_clk), .rst(f2186_rst), .rdata(f2186_rdata));
  assign f2186_clk = clk;
  assign f2186_rst = rst;
  // Bindings to f2186

  // f2188
  logic [0:0] f2188_wen;
  logic [31:0] f2188_wdata;
  logic [0:0] f2188_clk;
  logic [0:0] f2188_rst;
  logic [31:0] f2188_rdata;
  sr_buffer_32_1 f2188(.wen(f2188_wen), .wdata(f2188_wdata), .clk(f2188_clk), .rst(f2188_rst), .rdata(f2188_rdata));
  assign f2188_clk = clk;
  assign f2188_rst = rst;
  // Bindings to f2188

  // f2190
  logic [0:0] f2190_wen;
  logic [31:0] f2190_wdata;
  logic [0:0] f2190_clk;
  logic [0:0] f2190_rst;
  logic [31:0] f2190_rdata;
  sr_buffer_32_1 f2190(.wen(f2190_wen), .wdata(f2190_wdata), .clk(f2190_clk), .rst(f2190_rst), .rdata(f2190_rdata));
  assign f2190_clk = clk;
  assign f2190_rst = rst;
  // Bindings to f2190

  // f2192
  logic [0:0] f2192_wen;
  logic [31:0] f2192_wdata;
  logic [0:0] f2192_clk;
  logic [0:0] f2192_rst;
  logic [31:0] f2192_rdata;
  sr_buffer_32_1 f2192(.wen(f2192_wen), .wdata(f2192_wdata), .clk(f2192_clk), .rst(f2192_rst), .rdata(f2192_rdata));
  assign f2192_clk = clk;
  assign f2192_rst = rst;
  // Bindings to f2192

  // f2194
  logic [0:0] f2194_wen;
  logic [31:0] f2194_wdata;
  logic [0:0] f2194_clk;
  logic [0:0] f2194_rst;
  logic [31:0] f2194_rdata;
  sr_buffer_32_1 f2194(.wen(f2194_wen), .wdata(f2194_wdata), .clk(f2194_clk), .rst(f2194_rst), .rdata(f2194_rdata));
  assign f2194_clk = clk;
  assign f2194_rst = rst;
  // Bindings to f2194

  // f2196
  logic [0:0] f2196_wen;
  logic [31:0] f2196_wdata;
  logic [0:0] f2196_clk;
  logic [0:0] f2196_rst;
  logic [31:0] f2196_rdata;
  sr_buffer_32_1 f2196(.wen(f2196_wen), .wdata(f2196_wdata), .clk(f2196_clk), .rst(f2196_rst), .rdata(f2196_rdata));
  assign f2196_clk = clk;
  assign f2196_rst = rst;
  // Bindings to f2196

  // f2198
  logic [0:0] f2198_wen;
  logic [31:0] f2198_wdata;
  logic [0:0] f2198_clk;
  logic [0:0] f2198_rst;
  logic [31:0] f2198_rdata;
  sr_buffer_32_1 f2198(.wen(f2198_wen), .wdata(f2198_wdata), .clk(f2198_clk), .rst(f2198_rst), .rdata(f2198_rdata));
  assign f2198_clk = clk;
  assign f2198_rst = rst;
  // Bindings to f2198

  // f2200
  logic [0:0] f2200_wen;
  logic [31:0] f2200_wdata;
  logic [0:0] f2200_clk;
  logic [0:0] f2200_rst;
  logic [31:0] f2200_rdata;
  sr_buffer_32_1 f2200(.wen(f2200_wen), .wdata(f2200_wdata), .clk(f2200_clk), .rst(f2200_rst), .rdata(f2200_rdata));
  assign f2200_clk = clk;
  assign f2200_rst = rst;
  // Bindings to f2200

  // f2202
  logic [0:0] f2202_wen;
  logic [31:0] f2202_wdata;
  logic [0:0] f2202_clk;
  logic [0:0] f2202_rst;
  logic [31:0] f2202_rdata;
  sr_buffer_32_1 f2202(.wen(f2202_wen), .wdata(f2202_wdata), .clk(f2202_clk), .rst(f2202_rst), .rdata(f2202_rdata));
  assign f2202_clk = clk;
  assign f2202_rst = rst;
  // Bindings to f2202

  // f2204
  logic [0:0] f2204_wen;
  logic [31:0] f2204_wdata;
  logic [0:0] f2204_clk;
  logic [0:0] f2204_rst;
  logic [31:0] f2204_rdata;
  sr_buffer_32_1 f2204(.wen(f2204_wen), .wdata(f2204_wdata), .clk(f2204_clk), .rst(f2204_rst), .rdata(f2204_rdata));
  assign f2204_clk = clk;
  assign f2204_rst = rst;
  // Bindings to f2204

  // f2206
  logic [0:0] f2206_wen;
  logic [31:0] f2206_wdata;
  logic [0:0] f2206_clk;
  logic [0:0] f2206_rst;
  logic [31:0] f2206_rdata;
  sr_buffer_32_1 f2206(.wen(f2206_wen), .wdata(f2206_wdata), .clk(f2206_clk), .rst(f2206_rst), .rdata(f2206_rdata));
  assign f2206_clk = clk;
  assign f2206_rst = rst;
  // Bindings to f2206

  // f2208
  logic [0:0] f2208_wen;
  logic [31:0] f2208_wdata;
  logic [0:0] f2208_clk;
  logic [0:0] f2208_rst;
  logic [31:0] f2208_rdata;
  sr_buffer_32_1 f2208(.wen(f2208_wen), .wdata(f2208_wdata), .clk(f2208_clk), .rst(f2208_rst), .rdata(f2208_rdata));
  assign f2208_clk = clk;
  assign f2208_rst = rst;
  // Bindings to f2208

  // f2210
  logic [0:0] f2210_wen;
  logic [31:0] f2210_wdata;
  logic [0:0] f2210_clk;
  logic [0:0] f2210_rst;
  logic [31:0] f2210_rdata;
  sr_buffer_32_1 f2210(.wen(f2210_wen), .wdata(f2210_wdata), .clk(f2210_clk), .rst(f2210_rst), .rdata(f2210_rdata));
  assign f2210_clk = clk;
  assign f2210_rst = rst;
  // Bindings to f2210

  // f2212
  logic [0:0] f2212_wen;
  logic [31:0] f2212_wdata;
  logic [0:0] f2212_clk;
  logic [0:0] f2212_rst;
  logic [31:0] f2212_rdata;
  sr_buffer_32_1 f2212(.wen(f2212_wen), .wdata(f2212_wdata), .clk(f2212_clk), .rst(f2212_rst), .rdata(f2212_rdata));
  assign f2212_clk = clk;
  assign f2212_rst = rst;
  // Bindings to f2212

  // f2214
  logic [0:0] f2214_wen;
  logic [31:0] f2214_wdata;
  logic [0:0] f2214_clk;
  logic [0:0] f2214_rst;
  logic [31:0] f2214_rdata;
  sr_buffer_32_1 f2214(.wen(f2214_wen), .wdata(f2214_wdata), .clk(f2214_clk), .rst(f2214_rst), .rdata(f2214_rdata));
  assign f2214_clk = clk;
  assign f2214_rst = rst;
  // Bindings to f2214

  // f2216
  logic [0:0] f2216_wen;
  logic [31:0] f2216_wdata;
  logic [0:0] f2216_clk;
  logic [0:0] f2216_rst;
  logic [31:0] f2216_rdata;
  sr_buffer_32_1 f2216(.wen(f2216_wen), .wdata(f2216_wdata), .clk(f2216_clk), .rst(f2216_rst), .rdata(f2216_rdata));
  assign f2216_clk = clk;
  assign f2216_rst = rst;
  // Bindings to f2216

  // f2218
  logic [0:0] f2218_wen;
  logic [31:0] f2218_wdata;
  logic [0:0] f2218_clk;
  logic [0:0] f2218_rst;
  logic [31:0] f2218_rdata;
  sr_buffer_32_1 f2218(.wen(f2218_wen), .wdata(f2218_wdata), .clk(f2218_clk), .rst(f2218_rst), .rdata(f2218_rdata));
  assign f2218_clk = clk;
  assign f2218_rst = rst;
  // Bindings to f2218

  // f2220
  logic [0:0] f2220_wen;
  logic [31:0] f2220_wdata;
  logic [0:0] f2220_clk;
  logic [0:0] f2220_rst;
  logic [31:0] f2220_rdata;
  sr_buffer_32_1 f2220(.wen(f2220_wen), .wdata(f2220_wdata), .clk(f2220_clk), .rst(f2220_rst), .rdata(f2220_rdata));
  assign f2220_clk = clk;
  assign f2220_rst = rst;
  // Bindings to f2220

  // f2222
  logic [0:0] f2222_wen;
  logic [31:0] f2222_wdata;
  logic [0:0] f2222_clk;
  logic [0:0] f2222_rst;
  logic [31:0] f2222_rdata;
  sr_buffer_32_1 f2222(.wen(f2222_wen), .wdata(f2222_wdata), .clk(f2222_clk), .rst(f2222_rst), .rdata(f2222_rdata));
  assign f2222_clk = clk;
  assign f2222_rst = rst;
  // Bindings to f2222

  // f2224
  logic [0:0] f2224_wen;
  logic [31:0] f2224_wdata;
  logic [0:0] f2224_clk;
  logic [0:0] f2224_rst;
  logic [31:0] f2224_rdata;
  sr_buffer_32_1 f2224(.wen(f2224_wen), .wdata(f2224_wdata), .clk(f2224_clk), .rst(f2224_rst), .rdata(f2224_rdata));
  assign f2224_clk = clk;
  assign f2224_rst = rst;
  // Bindings to f2224

  // f2226
  logic [0:0] f2226_wen;
  logic [31:0] f2226_wdata;
  logic [0:0] f2226_clk;
  logic [0:0] f2226_rst;
  logic [31:0] f2226_rdata;
  sr_buffer_32_1 f2226(.wen(f2226_wen), .wdata(f2226_wdata), .clk(f2226_clk), .rst(f2226_rst), .rdata(f2226_rdata));
  assign f2226_clk = clk;
  assign f2226_rst = rst;
  // Bindings to f2226

  // f2228
  logic [0:0] f2228_wen;
  logic [31:0] f2228_wdata;
  logic [0:0] f2228_clk;
  logic [0:0] f2228_rst;
  logic [31:0] f2228_rdata;
  sr_buffer_32_1 f2228(.wen(f2228_wen), .wdata(f2228_wdata), .clk(f2228_clk), .rst(f2228_rst), .rdata(f2228_rdata));
  assign f2228_clk = clk;
  assign f2228_rst = rst;
  // Bindings to f2228

  // f2230
  logic [0:0] f2230_wen;
  logic [31:0] f2230_wdata;
  logic [0:0] f2230_clk;
  logic [0:0] f2230_rst;
  logic [31:0] f2230_rdata;
  sr_buffer_32_1 f2230(.wen(f2230_wen), .wdata(f2230_wdata), .clk(f2230_clk), .rst(f2230_rst), .rdata(f2230_rdata));
  assign f2230_clk = clk;
  assign f2230_rst = rst;
  // Bindings to f2230

  // f2232
  logic [0:0] f2232_wen;
  logic [31:0] f2232_wdata;
  logic [0:0] f2232_clk;
  logic [0:0] f2232_rst;
  logic [31:0] f2232_rdata;
  sr_buffer_32_1 f2232(.wen(f2232_wen), .wdata(f2232_wdata), .clk(f2232_clk), .rst(f2232_rst), .rdata(f2232_rdata));
  assign f2232_clk = clk;
  assign f2232_rst = rst;
  // Bindings to f2232

  // f2234
  logic [0:0] f2234_wen;
  logic [31:0] f2234_wdata;
  logic [0:0] f2234_clk;
  logic [0:0] f2234_rst;
  logic [31:0] f2234_rdata;
  sr_buffer_32_1 f2234(.wen(f2234_wen), .wdata(f2234_wdata), .clk(f2234_clk), .rst(f2234_rst), .rdata(f2234_rdata));
  assign f2234_clk = clk;
  assign f2234_rst = rst;
  // Bindings to f2234

  // f2236
  logic [0:0] f2236_wen;
  logic [31:0] f2236_wdata;
  logic [0:0] f2236_clk;
  logic [0:0] f2236_rst;
  logic [31:0] f2236_rdata;
  sr_buffer_32_1 f2236(.wen(f2236_wen), .wdata(f2236_wdata), .clk(f2236_clk), .rst(f2236_rst), .rdata(f2236_rdata));
  assign f2236_clk = clk;
  assign f2236_rst = rst;
  // Bindings to f2236

  // f2238
  logic [0:0] f2238_wen;
  logic [31:0] f2238_wdata;
  logic [0:0] f2238_clk;
  logic [0:0] f2238_rst;
  logic [31:0] f2238_rdata;
  sr_buffer_32_1 f2238(.wen(f2238_wen), .wdata(f2238_wdata), .clk(f2238_clk), .rst(f2238_rst), .rdata(f2238_rdata));
  assign f2238_clk = clk;
  assign f2238_rst = rst;
  // Bindings to f2238

  // f2240
  logic [0:0] f2240_wen;
  logic [31:0] f2240_wdata;
  logic [0:0] f2240_clk;
  logic [0:0] f2240_rst;
  logic [31:0] f2240_rdata;
  sr_buffer_32_1 f2240(.wen(f2240_wen), .wdata(f2240_wdata), .clk(f2240_clk), .rst(f2240_rst), .rdata(f2240_rdata));
  assign f2240_clk = clk;
  assign f2240_rst = rst;
  // Bindings to f2240

  // f2242
  logic [0:0] f2242_wen;
  logic [31:0] f2242_wdata;
  logic [0:0] f2242_clk;
  logic [0:0] f2242_rst;
  logic [31:0] f2242_rdata;
  sr_buffer_32_1 f2242(.wen(f2242_wen), .wdata(f2242_wdata), .clk(f2242_clk), .rst(f2242_rst), .rdata(f2242_rdata));
  assign f2242_clk = clk;
  assign f2242_rst = rst;
  // Bindings to f2242

  // f2244
  logic [0:0] f2244_wen;
  logic [31:0] f2244_wdata;
  logic [0:0] f2244_clk;
  logic [0:0] f2244_rst;
  logic [31:0] f2244_rdata;
  sr_buffer_32_1 f2244(.wen(f2244_wen), .wdata(f2244_wdata), .clk(f2244_clk), .rst(f2244_rst), .rdata(f2244_rdata));
  assign f2244_clk = clk;
  assign f2244_rst = rst;
  // Bindings to f2244

  // f2246
  logic [0:0] f2246_wen;
  logic [31:0] f2246_wdata;
  logic [0:0] f2246_clk;
  logic [0:0] f2246_rst;
  logic [31:0] f2246_rdata;
  sr_buffer_32_1 f2246(.wen(f2246_wen), .wdata(f2246_wdata), .clk(f2246_clk), .rst(f2246_rst), .rdata(f2246_rdata));
  assign f2246_clk = clk;
  assign f2246_rst = rst;
  // Bindings to f2246

  // f2248
  logic [0:0] f2248_wen;
  logic [31:0] f2248_wdata;
  logic [0:0] f2248_clk;
  logic [0:0] f2248_rst;
  logic [31:0] f2248_rdata;
  sr_buffer_32_1 f2248(.wen(f2248_wen), .wdata(f2248_wdata), .clk(f2248_clk), .rst(f2248_rst), .rdata(f2248_rdata));
  assign f2248_clk = clk;
  assign f2248_rst = rst;
  // Bindings to f2248

  // f2250
  logic [0:0] f2250_wen;
  logic [31:0] f2250_wdata;
  logic [0:0] f2250_clk;
  logic [0:0] f2250_rst;
  logic [31:0] f2250_rdata;
  sr_buffer_32_1 f2250(.wen(f2250_wen), .wdata(f2250_wdata), .clk(f2250_clk), .rst(f2250_rst), .rdata(f2250_rdata));
  assign f2250_clk = clk;
  assign f2250_rst = rst;
  // Bindings to f2250

  // f2252
  logic [0:0] f2252_wen;
  logic [31:0] f2252_wdata;
  logic [0:0] f2252_clk;
  logic [0:0] f2252_rst;
  logic [31:0] f2252_rdata;
  sr_buffer_32_1 f2252(.wen(f2252_wen), .wdata(f2252_wdata), .clk(f2252_clk), .rst(f2252_rst), .rdata(f2252_rdata));
  assign f2252_clk = clk;
  assign f2252_rst = rst;
  // Bindings to f2252

  // f2254
  logic [0:0] f2254_wen;
  logic [31:0] f2254_wdata;
  logic [0:0] f2254_clk;
  logic [0:0] f2254_rst;
  logic [31:0] f2254_rdata;
  sr_buffer_32_1 f2254(.wen(f2254_wen), .wdata(f2254_wdata), .clk(f2254_clk), .rst(f2254_rst), .rdata(f2254_rdata));
  assign f2254_clk = clk;
  assign f2254_rst = rst;
  // Bindings to f2254

  // f2256
  logic [0:0] f2256_wen;
  logic [31:0] f2256_wdata;
  logic [0:0] f2256_clk;
  logic [0:0] f2256_rst;
  logic [31:0] f2256_rdata;
  sr_buffer_32_1 f2256(.wen(f2256_wen), .wdata(f2256_wdata), .clk(f2256_clk), .rst(f2256_rst), .rdata(f2256_rdata));
  assign f2256_clk = clk;
  assign f2256_rst = rst;
  // Bindings to f2256

  // f2258
  logic [0:0] f2258_wen;
  logic [31:0] f2258_wdata;
  logic [0:0] f2258_clk;
  logic [0:0] f2258_rst;
  logic [31:0] f2258_rdata;
  sr_buffer_32_1 f2258(.wen(f2258_wen), .wdata(f2258_wdata), .clk(f2258_clk), .rst(f2258_rst), .rdata(f2258_rdata));
  assign f2258_clk = clk;
  assign f2258_rst = rst;
  // Bindings to f2258

  // f2260
  logic [0:0] f2260_wen;
  logic [31:0] f2260_wdata;
  logic [0:0] f2260_clk;
  logic [0:0] f2260_rst;
  logic [31:0] f2260_rdata;
  sr_buffer_32_1 f2260(.wen(f2260_wen), .wdata(f2260_wdata), .clk(f2260_clk), .rst(f2260_rst), .rdata(f2260_rdata));
  assign f2260_clk = clk;
  assign f2260_rst = rst;
  // Bindings to f2260

  // f2262
  logic [0:0] f2262_wen;
  logic [31:0] f2262_wdata;
  logic [0:0] f2262_clk;
  logic [0:0] f2262_rst;
  logic [31:0] f2262_rdata;
  sr_buffer_32_1 f2262(.wen(f2262_wen), .wdata(f2262_wdata), .clk(f2262_clk), .rst(f2262_rst), .rdata(f2262_rdata));
  assign f2262_clk = clk;
  assign f2262_rst = rst;
  // Bindings to f2262

  // f2264
  logic [0:0] f2264_wen;
  logic [31:0] f2264_wdata;
  logic [0:0] f2264_clk;
  logic [0:0] f2264_rst;
  logic [31:0] f2264_rdata;
  sr_buffer_32_1 f2264(.wen(f2264_wen), .wdata(f2264_wdata), .clk(f2264_clk), .rst(f2264_rst), .rdata(f2264_rdata));
  assign f2264_clk = clk;
  assign f2264_rst = rst;
  // Bindings to f2264

  // f2266
  logic [0:0] f2266_wen;
  logic [31:0] f2266_wdata;
  logic [0:0] f2266_clk;
  logic [0:0] f2266_rst;
  logic [31:0] f2266_rdata;
  sr_buffer_32_1 f2266(.wen(f2266_wen), .wdata(f2266_wdata), .clk(f2266_clk), .rst(f2266_rst), .rdata(f2266_rdata));
  assign f2266_clk = clk;
  assign f2266_rst = rst;
  // Bindings to f2266

  // f2268
  logic [0:0] f2268_wen;
  logic [31:0] f2268_wdata;
  logic [0:0] f2268_clk;
  logic [0:0] f2268_rst;
  logic [31:0] f2268_rdata;
  sr_buffer_32_1 f2268(.wen(f2268_wen), .wdata(f2268_wdata), .clk(f2268_clk), .rst(f2268_rst), .rdata(f2268_rdata));
  assign f2268_clk = clk;
  assign f2268_rst = rst;
  // Bindings to f2268

  // f2270
  logic [0:0] f2270_wen;
  logic [31:0] f2270_wdata;
  logic [0:0] f2270_clk;
  logic [0:0] f2270_rst;
  logic [31:0] f2270_rdata;
  sr_buffer_32_1 f2270(.wen(f2270_wen), .wdata(f2270_wdata), .clk(f2270_clk), .rst(f2270_rst), .rdata(f2270_rdata));
  assign f2270_clk = clk;
  assign f2270_rst = rst;
  // Bindings to f2270

  // f2272
  logic [0:0] f2272_wen;
  logic [31:0] f2272_wdata;
  logic [0:0] f2272_clk;
  logic [0:0] f2272_rst;
  logic [31:0] f2272_rdata;
  sr_buffer_32_1 f2272(.wen(f2272_wen), .wdata(f2272_wdata), .clk(f2272_clk), .rst(f2272_rst), .rdata(f2272_rdata));
  assign f2272_clk = clk;
  assign f2272_rst = rst;
  // Bindings to f2272

  // f2274
  logic [0:0] f2274_wen;
  logic [31:0] f2274_wdata;
  logic [0:0] f2274_clk;
  logic [0:0] f2274_rst;
  logic [31:0] f2274_rdata;
  sr_buffer_32_1 f2274(.wen(f2274_wen), .wdata(f2274_wdata), .clk(f2274_clk), .rst(f2274_rst), .rdata(f2274_rdata));
  assign f2274_clk = clk;
  assign f2274_rst = rst;
  // Bindings to f2274

  // f2276
  logic [0:0] f2276_wen;
  logic [31:0] f2276_wdata;
  logic [0:0] f2276_clk;
  logic [0:0] f2276_rst;
  logic [31:0] f2276_rdata;
  sr_buffer_32_1 f2276(.wen(f2276_wen), .wdata(f2276_wdata), .clk(f2276_clk), .rst(f2276_rst), .rdata(f2276_rdata));
  assign f2276_clk = clk;
  assign f2276_rst = rst;
  // Bindings to f2276

  // f2278
  logic [0:0] f2278_wen;
  logic [31:0] f2278_wdata;
  logic [0:0] f2278_clk;
  logic [0:0] f2278_rst;
  logic [31:0] f2278_rdata;
  sr_buffer_32_1 f2278(.wen(f2278_wen), .wdata(f2278_wdata), .clk(f2278_clk), .rst(f2278_rst), .rdata(f2278_rdata));
  assign f2278_clk = clk;
  assign f2278_rst = rst;
  // Bindings to f2278

  // f2280
  logic [0:0] f2280_wen;
  logic [31:0] f2280_wdata;
  logic [0:0] f2280_clk;
  logic [0:0] f2280_rst;
  logic [31:0] f2280_rdata;
  sr_buffer_32_1 f2280(.wen(f2280_wen), .wdata(f2280_wdata), .clk(f2280_clk), .rst(f2280_rst), .rdata(f2280_rdata));
  assign f2280_clk = clk;
  assign f2280_rst = rst;
  // Bindings to f2280

  // f2282
  logic [0:0] f2282_wen;
  logic [31:0] f2282_wdata;
  logic [0:0] f2282_clk;
  logic [0:0] f2282_rst;
  logic [31:0] f2282_rdata;
  sr_buffer_32_1 f2282(.wen(f2282_wen), .wdata(f2282_wdata), .clk(f2282_clk), .rst(f2282_rst), .rdata(f2282_rdata));
  assign f2282_clk = clk;
  assign f2282_rst = rst;
  // Bindings to f2282

  // f2284
  logic [0:0] f2284_wen;
  logic [31:0] f2284_wdata;
  logic [0:0] f2284_clk;
  logic [0:0] f2284_rst;
  logic [31:0] f2284_rdata;
  sr_buffer_32_1 f2284(.wen(f2284_wen), .wdata(f2284_wdata), .clk(f2284_clk), .rst(f2284_rst), .rdata(f2284_rdata));
  assign f2284_clk = clk;
  assign f2284_rst = rst;
  // Bindings to f2284

  // f2286
  logic [0:0] f2286_wen;
  logic [31:0] f2286_wdata;
  logic [0:0] f2286_clk;
  logic [0:0] f2286_rst;
  logic [31:0] f2286_rdata;
  sr_buffer_32_1 f2286(.wen(f2286_wen), .wdata(f2286_wdata), .clk(f2286_clk), .rst(f2286_rst), .rdata(f2286_rdata));
  assign f2286_clk = clk;
  assign f2286_rst = rst;
  // Bindings to f2286

  // f2288
  logic [0:0] f2288_wen;
  logic [31:0] f2288_wdata;
  logic [0:0] f2288_clk;
  logic [0:0] f2288_rst;
  logic [31:0] f2288_rdata;
  sr_buffer_32_1 f2288(.wen(f2288_wen), .wdata(f2288_wdata), .clk(f2288_clk), .rst(f2288_rst), .rdata(f2288_rdata));
  assign f2288_clk = clk;
  assign f2288_rst = rst;
  // Bindings to f2288

  // f2290
  logic [0:0] f2290_wen;
  logic [31:0] f2290_wdata;
  logic [0:0] f2290_clk;
  logic [0:0] f2290_rst;
  logic [31:0] f2290_rdata;
  sr_buffer_32_1 f2290(.wen(f2290_wen), .wdata(f2290_wdata), .clk(f2290_clk), .rst(f2290_rst), .rdata(f2290_rdata));
  assign f2290_clk = clk;
  assign f2290_rst = rst;
  // Bindings to f2290

  // f2292
  logic [0:0] f2292_wen;
  logic [31:0] f2292_wdata;
  logic [0:0] f2292_clk;
  logic [0:0] f2292_rst;
  logic [31:0] f2292_rdata;
  sr_buffer_32_1 f2292(.wen(f2292_wen), .wdata(f2292_wdata), .clk(f2292_clk), .rst(f2292_rst), .rdata(f2292_rdata));
  assign f2292_clk = clk;
  assign f2292_rst = rst;
  // Bindings to f2292

  // f2294
  logic [0:0] f2294_wen;
  logic [31:0] f2294_wdata;
  logic [0:0] f2294_clk;
  logic [0:0] f2294_rst;
  logic [31:0] f2294_rdata;
  sr_buffer_32_1 f2294(.wen(f2294_wen), .wdata(f2294_wdata), .clk(f2294_clk), .rst(f2294_rst), .rdata(f2294_rdata));
  assign f2294_clk = clk;
  assign f2294_rst = rst;
  // Bindings to f2294

  // f2296
  logic [0:0] f2296_wen;
  logic [31:0] f2296_wdata;
  logic [0:0] f2296_clk;
  logic [0:0] f2296_rst;
  logic [31:0] f2296_rdata;
  sr_buffer_32_1 f2296(.wen(f2296_wen), .wdata(f2296_wdata), .clk(f2296_clk), .rst(f2296_rst), .rdata(f2296_rdata));
  assign f2296_clk = clk;
  assign f2296_rst = rst;
  // Bindings to f2296

  // f2298
  logic [0:0] f2298_wen;
  logic [31:0] f2298_wdata;
  logic [0:0] f2298_clk;
  logic [0:0] f2298_rst;
  logic [31:0] f2298_rdata;
  sr_buffer_32_1 f2298(.wen(f2298_wen), .wdata(f2298_wdata), .clk(f2298_clk), .rst(f2298_rst), .rdata(f2298_rdata));
  assign f2298_clk = clk;
  assign f2298_rst = rst;
  // Bindings to f2298

  // f2300
  logic [0:0] f2300_wen;
  logic [31:0] f2300_wdata;
  logic [0:0] f2300_clk;
  logic [0:0] f2300_rst;
  logic [31:0] f2300_rdata;
  sr_buffer_32_1 f2300(.wen(f2300_wen), .wdata(f2300_wdata), .clk(f2300_clk), .rst(f2300_rst), .rdata(f2300_rdata));
  assign f2300_clk = clk;
  assign f2300_rst = rst;
  // Bindings to f2300

  // f2302
  logic [0:0] f2302_wen;
  logic [31:0] f2302_wdata;
  logic [0:0] f2302_clk;
  logic [0:0] f2302_rst;
  logic [31:0] f2302_rdata;
  sr_buffer_32_1 f2302(.wen(f2302_wen), .wdata(f2302_wdata), .clk(f2302_clk), .rst(f2302_rst), .rdata(f2302_rdata));
  assign f2302_clk = clk;
  assign f2302_rst = rst;
  // Bindings to f2302

  // f2304
  logic [0:0] f2304_wen;
  logic [31:0] f2304_wdata;
  logic [0:0] f2304_clk;
  logic [0:0] f2304_rst;
  logic [31:0] f2304_rdata;
  sr_buffer_32_1 f2304(.wen(f2304_wen), .wdata(f2304_wdata), .clk(f2304_clk), .rst(f2304_rst), .rdata(f2304_rdata));
  assign f2304_clk = clk;
  assign f2304_rst = rst;
  // Bindings to f2304

  // f2306
  logic [0:0] f2306_wen;
  logic [31:0] f2306_wdata;
  logic [0:0] f2306_clk;
  logic [0:0] f2306_rst;
  logic [31:0] f2306_rdata;
  sr_buffer_32_1 f2306(.wen(f2306_wen), .wdata(f2306_wdata), .clk(f2306_clk), .rst(f2306_rst), .rdata(f2306_rdata));
  assign f2306_clk = clk;
  assign f2306_rst = rst;
  // Bindings to f2306

  // f2308
  logic [0:0] f2308_wen;
  logic [31:0] f2308_wdata;
  logic [0:0] f2308_clk;
  logic [0:0] f2308_rst;
  logic [31:0] f2308_rdata;
  sr_buffer_32_1 f2308(.wen(f2308_wen), .wdata(f2308_wdata), .clk(f2308_clk), .rst(f2308_rst), .rdata(f2308_rdata));
  assign f2308_clk = clk;
  assign f2308_rst = rst;
  // Bindings to f2308

  // f2310
  logic [0:0] f2310_wen;
  logic [31:0] f2310_wdata;
  logic [0:0] f2310_clk;
  logic [0:0] f2310_rst;
  logic [31:0] f2310_rdata;
  sr_buffer_32_1 f2310(.wen(f2310_wen), .wdata(f2310_wdata), .clk(f2310_clk), .rst(f2310_rst), .rdata(f2310_rdata));
  assign f2310_clk = clk;
  assign f2310_rst = rst;
  // Bindings to f2310

  // f2312
  logic [0:0] f2312_wen;
  logic [31:0] f2312_wdata;
  logic [0:0] f2312_clk;
  logic [0:0] f2312_rst;
  logic [31:0] f2312_rdata;
  sr_buffer_32_1 f2312(.wen(f2312_wen), .wdata(f2312_wdata), .clk(f2312_clk), .rst(f2312_rst), .rdata(f2312_rdata));
  assign f2312_clk = clk;
  assign f2312_rst = rst;
  // Bindings to f2312

  // f2314
  logic [0:0] f2314_wen;
  logic [31:0] f2314_wdata;
  logic [0:0] f2314_clk;
  logic [0:0] f2314_rst;
  logic [31:0] f2314_rdata;
  sr_buffer_32_1 f2314(.wen(f2314_wen), .wdata(f2314_wdata), .clk(f2314_clk), .rst(f2314_rst), .rdata(f2314_rdata));
  assign f2314_clk = clk;
  assign f2314_rst = rst;
  // Bindings to f2314

  // f2316
  logic [0:0] f2316_wen;
  logic [31:0] f2316_wdata;
  logic [0:0] f2316_clk;
  logic [0:0] f2316_rst;
  logic [31:0] f2316_rdata;
  sr_buffer_32_1 f2316(.wen(f2316_wen), .wdata(f2316_wdata), .clk(f2316_clk), .rst(f2316_rst), .rdata(f2316_rdata));
  assign f2316_clk = clk;
  assign f2316_rst = rst;
  // Bindings to f2316

  // f2318
  logic [0:0] f2318_wen;
  logic [31:0] f2318_wdata;
  logic [0:0] f2318_clk;
  logic [0:0] f2318_rst;
  logic [31:0] f2318_rdata;
  sr_buffer_32_1 f2318(.wen(f2318_wen), .wdata(f2318_wdata), .clk(f2318_clk), .rst(f2318_rst), .rdata(f2318_rdata));
  assign f2318_clk = clk;
  assign f2318_rst = rst;
  // Bindings to f2318

  // f2320
  logic [0:0] f2320_wen;
  logic [31:0] f2320_wdata;
  logic [0:0] f2320_clk;
  logic [0:0] f2320_rst;
  logic [31:0] f2320_rdata;
  sr_buffer_32_1 f2320(.wen(f2320_wen), .wdata(f2320_wdata), .clk(f2320_clk), .rst(f2320_rst), .rdata(f2320_rdata));
  assign f2320_clk = clk;
  assign f2320_rst = rst;
  // Bindings to f2320

  // f2322
  logic [0:0] f2322_wen;
  logic [31:0] f2322_wdata;
  logic [0:0] f2322_clk;
  logic [0:0] f2322_rst;
  logic [31:0] f2322_rdata;
  sr_buffer_32_1 f2322(.wen(f2322_wen), .wdata(f2322_wdata), .clk(f2322_clk), .rst(f2322_rst), .rdata(f2322_rdata));
  assign f2322_clk = clk;
  assign f2322_rst = rst;
  // Bindings to f2322

  // f2324
  logic [0:0] f2324_wen;
  logic [31:0] f2324_wdata;
  logic [0:0] f2324_clk;
  logic [0:0] f2324_rst;
  logic [31:0] f2324_rdata;
  sr_buffer_32_1 f2324(.wen(f2324_wen), .wdata(f2324_wdata), .clk(f2324_clk), .rst(f2324_rst), .rdata(f2324_rdata));
  assign f2324_clk = clk;
  assign f2324_rst = rst;
  // Bindings to f2324

  // f2326
  logic [0:0] f2326_wen;
  logic [31:0] f2326_wdata;
  logic [0:0] f2326_clk;
  logic [0:0] f2326_rst;
  logic [31:0] f2326_rdata;
  sr_buffer_32_1 f2326(.wen(f2326_wen), .wdata(f2326_wdata), .clk(f2326_clk), .rst(f2326_rst), .rdata(f2326_rdata));
  assign f2326_clk = clk;
  assign f2326_rst = rst;
  // Bindings to f2326

  // f2328
  logic [0:0] f2328_wen;
  logic [31:0] f2328_wdata;
  logic [0:0] f2328_clk;
  logic [0:0] f2328_rst;
  logic [31:0] f2328_rdata;
  sr_buffer_32_1 f2328(.wen(f2328_wen), .wdata(f2328_wdata), .clk(f2328_clk), .rst(f2328_rst), .rdata(f2328_rdata));
  assign f2328_clk = clk;
  assign f2328_rst = rst;
  // Bindings to f2328

  // f2330
  logic [0:0] f2330_wen;
  logic [31:0] f2330_wdata;
  logic [0:0] f2330_clk;
  logic [0:0] f2330_rst;
  logic [31:0] f2330_rdata;
  sr_buffer_32_1 f2330(.wen(f2330_wen), .wdata(f2330_wdata), .clk(f2330_clk), .rst(f2330_rst), .rdata(f2330_rdata));
  assign f2330_clk = clk;
  assign f2330_rst = rst;
  // Bindings to f2330

  // f2332
  logic [0:0] f2332_wen;
  logic [31:0] f2332_wdata;
  logic [0:0] f2332_clk;
  logic [0:0] f2332_rst;
  logic [31:0] f2332_rdata;
  sr_buffer_32_1 f2332(.wen(f2332_wen), .wdata(f2332_wdata), .clk(f2332_clk), .rst(f2332_rst), .rdata(f2332_rdata));
  assign f2332_clk = clk;
  assign f2332_rst = rst;
  // Bindings to f2332

  // f2334
  logic [0:0] f2334_wen;
  logic [31:0] f2334_wdata;
  logic [0:0] f2334_clk;
  logic [0:0] f2334_rst;
  logic [31:0] f2334_rdata;
  sr_buffer_32_1 f2334(.wen(f2334_wen), .wdata(f2334_wdata), .clk(f2334_clk), .rst(f2334_rst), .rdata(f2334_rdata));
  assign f2334_clk = clk;
  assign f2334_rst = rst;
  // Bindings to f2334

  // f2336
  logic [0:0] f2336_wen;
  logic [31:0] f2336_wdata;
  logic [0:0] f2336_clk;
  logic [0:0] f2336_rst;
  logic [31:0] f2336_rdata;
  sr_buffer_32_1 f2336(.wen(f2336_wen), .wdata(f2336_wdata), .clk(f2336_clk), .rst(f2336_rst), .rdata(f2336_rdata));
  assign f2336_clk = clk;
  assign f2336_rst = rst;
  // Bindings to f2336

  // f2338
  logic [0:0] f2338_wen;
  logic [31:0] f2338_wdata;
  logic [0:0] f2338_clk;
  logic [0:0] f2338_rst;
  logic [31:0] f2338_rdata;
  sr_buffer_32_1 f2338(.wen(f2338_wen), .wdata(f2338_wdata), .clk(f2338_clk), .rst(f2338_rst), .rdata(f2338_rdata));
  assign f2338_clk = clk;
  assign f2338_rst = rst;
  // Bindings to f2338

  // f2340
  logic [0:0] f2340_wen;
  logic [31:0] f2340_wdata;
  logic [0:0] f2340_clk;
  logic [0:0] f2340_rst;
  logic [31:0] f2340_rdata;
  sr_buffer_32_1 f2340(.wen(f2340_wen), .wdata(f2340_wdata), .clk(f2340_clk), .rst(f2340_rst), .rdata(f2340_rdata));
  assign f2340_clk = clk;
  assign f2340_rst = rst;
  // Bindings to f2340

  // f2342
  logic [0:0] f2342_wen;
  logic [31:0] f2342_wdata;
  logic [0:0] f2342_clk;
  logic [0:0] f2342_rst;
  logic [31:0] f2342_rdata;
  sr_buffer_32_1 f2342(.wen(f2342_wen), .wdata(f2342_wdata), .clk(f2342_clk), .rst(f2342_rst), .rdata(f2342_rdata));
  assign f2342_clk = clk;
  assign f2342_rst = rst;
  // Bindings to f2342

  // f2344
  logic [0:0] f2344_wen;
  logic [31:0] f2344_wdata;
  logic [0:0] f2344_clk;
  logic [0:0] f2344_rst;
  logic [31:0] f2344_rdata;
  sr_buffer_32_1 f2344(.wen(f2344_wen), .wdata(f2344_wdata), .clk(f2344_clk), .rst(f2344_rst), .rdata(f2344_rdata));
  assign f2344_clk = clk;
  assign f2344_rst = rst;
  // Bindings to f2344

  // f2346
  logic [0:0] f2346_wen;
  logic [31:0] f2346_wdata;
  logic [0:0] f2346_clk;
  logic [0:0] f2346_rst;
  logic [31:0] f2346_rdata;
  sr_buffer_32_1 f2346(.wen(f2346_wen), .wdata(f2346_wdata), .clk(f2346_clk), .rst(f2346_rst), .rdata(f2346_rdata));
  assign f2346_clk = clk;
  assign f2346_rst = rst;
  // Bindings to f2346

  // f2348
  logic [0:0] f2348_wen;
  logic [31:0] f2348_wdata;
  logic [0:0] f2348_clk;
  logic [0:0] f2348_rst;
  logic [31:0] f2348_rdata;
  sr_buffer_32_1 f2348(.wen(f2348_wen), .wdata(f2348_wdata), .clk(f2348_clk), .rst(f2348_rst), .rdata(f2348_rdata));
  assign f2348_clk = clk;
  assign f2348_rst = rst;
  // Bindings to f2348

  // f2350
  logic [0:0] f2350_wen;
  logic [31:0] f2350_wdata;
  logic [0:0] f2350_clk;
  logic [0:0] f2350_rst;
  logic [31:0] f2350_rdata;
  sr_buffer_32_1 f2350(.wen(f2350_wen), .wdata(f2350_wdata), .clk(f2350_clk), .rst(f2350_rst), .rdata(f2350_rdata));
  assign f2350_clk = clk;
  assign f2350_rst = rst;
  // Bindings to f2350

  // f2352
  logic [0:0] f2352_wen;
  logic [31:0] f2352_wdata;
  logic [0:0] f2352_clk;
  logic [0:0] f2352_rst;
  logic [31:0] f2352_rdata;
  sr_buffer_32_1 f2352(.wen(f2352_wen), .wdata(f2352_wdata), .clk(f2352_clk), .rst(f2352_rst), .rdata(f2352_rdata));
  assign f2352_clk = clk;
  assign f2352_rst = rst;
  // Bindings to f2352

  // f2354
  logic [0:0] f2354_wen;
  logic [31:0] f2354_wdata;
  logic [0:0] f2354_clk;
  logic [0:0] f2354_rst;
  logic [31:0] f2354_rdata;
  sr_buffer_32_1 f2354(.wen(f2354_wen), .wdata(f2354_wdata), .clk(f2354_clk), .rst(f2354_rst), .rdata(f2354_rdata));
  assign f2354_clk = clk;
  assign f2354_rst = rst;
  // Bindings to f2354

  // f2356
  logic [0:0] f2356_wen;
  logic [31:0] f2356_wdata;
  logic [0:0] f2356_clk;
  logic [0:0] f2356_rst;
  logic [31:0] f2356_rdata;
  sr_buffer_32_1 f2356(.wen(f2356_wen), .wdata(f2356_wdata), .clk(f2356_clk), .rst(f2356_rst), .rdata(f2356_rdata));
  assign f2356_clk = clk;
  assign f2356_rst = rst;
  // Bindings to f2356

  // f2358
  logic [0:0] f2358_wen;
  logic [31:0] f2358_wdata;
  logic [0:0] f2358_clk;
  logic [0:0] f2358_rst;
  logic [31:0] f2358_rdata;
  sr_buffer_32_1 f2358(.wen(f2358_wen), .wdata(f2358_wdata), .clk(f2358_clk), .rst(f2358_rst), .rdata(f2358_rdata));
  assign f2358_clk = clk;
  assign f2358_rst = rst;
  // Bindings to f2358

  // f2360
  logic [0:0] f2360_wen;
  logic [31:0] f2360_wdata;
  logic [0:0] f2360_clk;
  logic [0:0] f2360_rst;
  logic [31:0] f2360_rdata;
  sr_buffer_32_1 f2360(.wen(f2360_wen), .wdata(f2360_wdata), .clk(f2360_clk), .rst(f2360_rst), .rdata(f2360_rdata));
  assign f2360_clk = clk;
  assign f2360_rst = rst;
  // Bindings to f2360

  // f2362
  logic [0:0] f2362_wen;
  logic [31:0] f2362_wdata;
  logic [0:0] f2362_clk;
  logic [0:0] f2362_rst;
  logic [31:0] f2362_rdata;
  sr_buffer_32_1 f2362(.wen(f2362_wen), .wdata(f2362_wdata), .clk(f2362_clk), .rst(f2362_rst), .rdata(f2362_rdata));
  assign f2362_clk = clk;
  assign f2362_rst = rst;
  // Bindings to f2362

  // f2364
  logic [0:0] f2364_wen;
  logic [31:0] f2364_wdata;
  logic [0:0] f2364_clk;
  logic [0:0] f2364_rst;
  logic [31:0] f2364_rdata;
  sr_buffer_32_1 f2364(.wen(f2364_wen), .wdata(f2364_wdata), .clk(f2364_clk), .rst(f2364_rst), .rdata(f2364_rdata));
  assign f2364_clk = clk;
  assign f2364_rst = rst;
  // Bindings to f2364

  // f2366
  logic [0:0] f2366_wen;
  logic [31:0] f2366_wdata;
  logic [0:0] f2366_clk;
  logic [0:0] f2366_rst;
  logic [31:0] f2366_rdata;
  sr_buffer_32_1 f2366(.wen(f2366_wen), .wdata(f2366_wdata), .clk(f2366_clk), .rst(f2366_rst), .rdata(f2366_rdata));
  assign f2366_clk = clk;
  assign f2366_rst = rst;
  // Bindings to f2366

  // f2368
  logic [0:0] f2368_wen;
  logic [31:0] f2368_wdata;
  logic [0:0] f2368_clk;
  logic [0:0] f2368_rst;
  logic [31:0] f2368_rdata;
  sr_buffer_32_1 f2368(.wen(f2368_wen), .wdata(f2368_wdata), .clk(f2368_clk), .rst(f2368_rst), .rdata(f2368_rdata));
  assign f2368_clk = clk;
  assign f2368_rst = rst;
  // Bindings to f2368

  // f2370
  logic [0:0] f2370_wen;
  logic [31:0] f2370_wdata;
  logic [0:0] f2370_clk;
  logic [0:0] f2370_rst;
  logic [31:0] f2370_rdata;
  sr_buffer_32_1 f2370(.wen(f2370_wen), .wdata(f2370_wdata), .clk(f2370_clk), .rst(f2370_rst), .rdata(f2370_rdata));
  assign f2370_clk = clk;
  assign f2370_rst = rst;
  // Bindings to f2370

  // f2372
  logic [0:0] f2372_wen;
  logic [31:0] f2372_wdata;
  logic [0:0] f2372_clk;
  logic [0:0] f2372_rst;
  logic [31:0] f2372_rdata;
  sr_buffer_32_1 f2372(.wen(f2372_wen), .wdata(f2372_wdata), .clk(f2372_clk), .rst(f2372_rst), .rdata(f2372_rdata));
  assign f2372_clk = clk;
  assign f2372_rst = rst;
  // Bindings to f2372

  // f2374
  logic [0:0] f2374_wen;
  logic [31:0] f2374_wdata;
  logic [0:0] f2374_clk;
  logic [0:0] f2374_rst;
  logic [31:0] f2374_rdata;
  sr_buffer_32_1 f2374(.wen(f2374_wen), .wdata(f2374_wdata), .clk(f2374_clk), .rst(f2374_rst), .rdata(f2374_rdata));
  assign f2374_clk = clk;
  assign f2374_rst = rst;
  // Bindings to f2374

  // f2376
  logic [0:0] f2376_wen;
  logic [31:0] f2376_wdata;
  logic [0:0] f2376_clk;
  logic [0:0] f2376_rst;
  logic [31:0] f2376_rdata;
  sr_buffer_32_1 f2376(.wen(f2376_wen), .wdata(f2376_wdata), .clk(f2376_clk), .rst(f2376_rst), .rdata(f2376_rdata));
  assign f2376_clk = clk;
  assign f2376_rst = rst;
  // Bindings to f2376

  // f2378
  logic [0:0] f2378_wen;
  logic [31:0] f2378_wdata;
  logic [0:0] f2378_clk;
  logic [0:0] f2378_rst;
  logic [31:0] f2378_rdata;
  sr_buffer_32_1 f2378(.wen(f2378_wen), .wdata(f2378_wdata), .clk(f2378_clk), .rst(f2378_rst), .rdata(f2378_rdata));
  assign f2378_clk = clk;
  assign f2378_rst = rst;
  // Bindings to f2378

  // f2380
  logic [0:0] f2380_wen;
  logic [31:0] f2380_wdata;
  logic [0:0] f2380_clk;
  logic [0:0] f2380_rst;
  logic [31:0] f2380_rdata;
  sr_buffer_32_1 f2380(.wen(f2380_wen), .wdata(f2380_wdata), .clk(f2380_clk), .rst(f2380_rst), .rdata(f2380_rdata));
  assign f2380_clk = clk;
  assign f2380_rst = rst;
  // Bindings to f2380

  // f2382
  logic [0:0] f2382_wen;
  logic [31:0] f2382_wdata;
  logic [0:0] f2382_clk;
  logic [0:0] f2382_rst;
  logic [31:0] f2382_rdata;
  sr_buffer_32_1 f2382(.wen(f2382_wen), .wdata(f2382_wdata), .clk(f2382_clk), .rst(f2382_rst), .rdata(f2382_rdata));
  assign f2382_clk = clk;
  assign f2382_rst = rst;
  // Bindings to f2382

  // f2384
  logic [0:0] f2384_wen;
  logic [31:0] f2384_wdata;
  logic [0:0] f2384_clk;
  logic [0:0] f2384_rst;
  logic [31:0] f2384_rdata;
  sr_buffer_32_1 f2384(.wen(f2384_wen), .wdata(f2384_wdata), .clk(f2384_clk), .rst(f2384_rst), .rdata(f2384_rdata));
  assign f2384_clk = clk;
  assign f2384_rst = rst;
  // Bindings to f2384

  // f2386
  logic [0:0] f2386_wen;
  logic [31:0] f2386_wdata;
  logic [0:0] f2386_clk;
  logic [0:0] f2386_rst;
  logic [31:0] f2386_rdata;
  sr_buffer_32_1 f2386(.wen(f2386_wen), .wdata(f2386_wdata), .clk(f2386_clk), .rst(f2386_rst), .rdata(f2386_rdata));
  assign f2386_clk = clk;
  assign f2386_rst = rst;
  // Bindings to f2386

  // f2388
  logic [0:0] f2388_wen;
  logic [31:0] f2388_wdata;
  logic [0:0] f2388_clk;
  logic [0:0] f2388_rst;
  logic [31:0] f2388_rdata;
  sr_buffer_32_1 f2388(.wen(f2388_wen), .wdata(f2388_wdata), .clk(f2388_clk), .rst(f2388_rst), .rdata(f2388_rdata));
  assign f2388_clk = clk;
  assign f2388_rst = rst;
  // Bindings to f2388

  // f2390
  logic [0:0] f2390_wen;
  logic [31:0] f2390_wdata;
  logic [0:0] f2390_clk;
  logic [0:0] f2390_rst;
  logic [31:0] f2390_rdata;
  sr_buffer_32_1 f2390(.wen(f2390_wen), .wdata(f2390_wdata), .clk(f2390_clk), .rst(f2390_rst), .rdata(f2390_rdata));
  assign f2390_clk = clk;
  assign f2390_rst = rst;
  // Bindings to f2390

  // f2392
  logic [0:0] f2392_wen;
  logic [31:0] f2392_wdata;
  logic [0:0] f2392_clk;
  logic [0:0] f2392_rst;
  logic [31:0] f2392_rdata;
  sr_buffer_32_1 f2392(.wen(f2392_wen), .wdata(f2392_wdata), .clk(f2392_clk), .rst(f2392_rst), .rdata(f2392_rdata));
  assign f2392_clk = clk;
  assign f2392_rst = rst;
  // Bindings to f2392

  // f2394
  logic [0:0] f2394_wen;
  logic [31:0] f2394_wdata;
  logic [0:0] f2394_clk;
  logic [0:0] f2394_rst;
  logic [31:0] f2394_rdata;
  sr_buffer_32_1 f2394(.wen(f2394_wen), .wdata(f2394_wdata), .clk(f2394_clk), .rst(f2394_rst), .rdata(f2394_rdata));
  assign f2394_clk = clk;
  assign f2394_rst = rst;
  // Bindings to f2394

  // f2396
  logic [0:0] f2396_wen;
  logic [31:0] f2396_wdata;
  logic [0:0] f2396_clk;
  logic [0:0] f2396_rst;
  logic [31:0] f2396_rdata;
  sr_buffer_32_1 f2396(.wen(f2396_wen), .wdata(f2396_wdata), .clk(f2396_clk), .rst(f2396_rst), .rdata(f2396_rdata));
  assign f2396_clk = clk;
  assign f2396_rst = rst;
  // Bindings to f2396

  // f2398
  logic [0:0] f2398_wen;
  logic [31:0] f2398_wdata;
  logic [0:0] f2398_clk;
  logic [0:0] f2398_rst;
  logic [31:0] f2398_rdata;
  sr_buffer_32_1 f2398(.wen(f2398_wen), .wdata(f2398_wdata), .clk(f2398_clk), .rst(f2398_rst), .rdata(f2398_rdata));
  assign f2398_clk = clk;
  assign f2398_rst = rst;
  // Bindings to f2398

  // f2400
  logic [0:0] f2400_wen;
  logic [31:0] f2400_wdata;
  logic [0:0] f2400_clk;
  logic [0:0] f2400_rst;
  logic [31:0] f2400_rdata;
  sr_buffer_32_1 f2400(.wen(f2400_wen), .wdata(f2400_wdata), .clk(f2400_clk), .rst(f2400_rst), .rdata(f2400_rdata));
  assign f2400_clk = clk;
  assign f2400_rst = rst;
  // Bindings to f2400

  // f2402
  logic [0:0] f2402_wen;
  logic [31:0] f2402_wdata;
  logic [0:0] f2402_clk;
  logic [0:0] f2402_rst;
  logic [31:0] f2402_rdata;
  sr_buffer_32_1 f2402(.wen(f2402_wen), .wdata(f2402_wdata), .clk(f2402_clk), .rst(f2402_rst), .rdata(f2402_rdata));
  assign f2402_clk = clk;
  assign f2402_rst = rst;
  // Bindings to f2402

  // f2404
  logic [0:0] f2404_wen;
  logic [31:0] f2404_wdata;
  logic [0:0] f2404_clk;
  logic [0:0] f2404_rst;
  logic [31:0] f2404_rdata;
  sr_buffer_32_1 f2404(.wen(f2404_wen), .wdata(f2404_wdata), .clk(f2404_clk), .rst(f2404_rst), .rdata(f2404_rdata));
  assign f2404_clk = clk;
  assign f2404_rst = rst;
  // Bindings to f2404

  // f2406
  logic [0:0] f2406_wen;
  logic [31:0] f2406_wdata;
  logic [0:0] f2406_clk;
  logic [0:0] f2406_rst;
  logic [31:0] f2406_rdata;
  sr_buffer_32_1 f2406(.wen(f2406_wen), .wdata(f2406_wdata), .clk(f2406_clk), .rst(f2406_rst), .rdata(f2406_rdata));
  assign f2406_clk = clk;
  assign f2406_rst = rst;
  // Bindings to f2406

  // f2408
  logic [0:0] f2408_wen;
  logic [31:0] f2408_wdata;
  logic [0:0] f2408_clk;
  logic [0:0] f2408_rst;
  logic [31:0] f2408_rdata;
  sr_buffer_32_1 f2408(.wen(f2408_wen), .wdata(f2408_wdata), .clk(f2408_clk), .rst(f2408_rst), .rdata(f2408_rdata));
  assign f2408_clk = clk;
  assign f2408_rst = rst;
  // Bindings to f2408

  // f2410
  logic [0:0] f2410_wen;
  logic [31:0] f2410_wdata;
  logic [0:0] f2410_clk;
  logic [0:0] f2410_rst;
  logic [31:0] f2410_rdata;
  sr_buffer_32_1 f2410(.wen(f2410_wen), .wdata(f2410_wdata), .clk(f2410_clk), .rst(f2410_rst), .rdata(f2410_rdata));
  assign f2410_clk = clk;
  assign f2410_rst = rst;
  // Bindings to f2410

  // f2412
  logic [0:0] f2412_wen;
  logic [31:0] f2412_wdata;
  logic [0:0] f2412_clk;
  logic [0:0] f2412_rst;
  logic [31:0] f2412_rdata;
  sr_buffer_32_1 f2412(.wen(f2412_wen), .wdata(f2412_wdata), .clk(f2412_clk), .rst(f2412_rst), .rdata(f2412_rdata));
  assign f2412_clk = clk;
  assign f2412_rst = rst;
  // Bindings to f2412

  // f2414
  logic [0:0] f2414_wen;
  logic [31:0] f2414_wdata;
  logic [0:0] f2414_clk;
  logic [0:0] f2414_rst;
  logic [31:0] f2414_rdata;
  sr_buffer_32_1 f2414(.wen(f2414_wen), .wdata(f2414_wdata), .clk(f2414_clk), .rst(f2414_rst), .rdata(f2414_rdata));
  assign f2414_clk = clk;
  assign f2414_rst = rst;
  // Bindings to f2414

  // f2416
  logic [0:0] f2416_wen;
  logic [31:0] f2416_wdata;
  logic [0:0] f2416_clk;
  logic [0:0] f2416_rst;
  logic [31:0] f2416_rdata;
  sr_buffer_32_1 f2416(.wen(f2416_wen), .wdata(f2416_wdata), .clk(f2416_clk), .rst(f2416_rst), .rdata(f2416_rdata));
  assign f2416_clk = clk;
  assign f2416_rst = rst;
  // Bindings to f2416

  // f2418
  logic [0:0] f2418_wen;
  logic [31:0] f2418_wdata;
  logic [0:0] f2418_clk;
  logic [0:0] f2418_rst;
  logic [31:0] f2418_rdata;
  sr_buffer_32_1 f2418(.wen(f2418_wen), .wdata(f2418_wdata), .clk(f2418_clk), .rst(f2418_rst), .rdata(f2418_rdata));
  assign f2418_clk = clk;
  assign f2418_rst = rst;
  // Bindings to f2418

  // f2420
  logic [0:0] f2420_wen;
  logic [31:0] f2420_wdata;
  logic [0:0] f2420_clk;
  logic [0:0] f2420_rst;
  logic [31:0] f2420_rdata;
  sr_buffer_32_1 f2420(.wen(f2420_wen), .wdata(f2420_wdata), .clk(f2420_clk), .rst(f2420_rst), .rdata(f2420_rdata));
  assign f2420_clk = clk;
  assign f2420_rst = rst;
  // Bindings to f2420

  // f2422
  logic [0:0] f2422_wen;
  logic [31:0] f2422_wdata;
  logic [0:0] f2422_clk;
  logic [0:0] f2422_rst;
  logic [31:0] f2422_rdata;
  sr_buffer_32_1 f2422(.wen(f2422_wen), .wdata(f2422_wdata), .clk(f2422_clk), .rst(f2422_rst), .rdata(f2422_rdata));
  assign f2422_clk = clk;
  assign f2422_rst = rst;
  // Bindings to f2422

  // f2424
  logic [0:0] f2424_wen;
  logic [31:0] f2424_wdata;
  logic [0:0] f2424_clk;
  logic [0:0] f2424_rst;
  logic [31:0] f2424_rdata;
  sr_buffer_32_1 f2424(.wen(f2424_wen), .wdata(f2424_wdata), .clk(f2424_clk), .rst(f2424_rst), .rdata(f2424_rdata));
  assign f2424_clk = clk;
  assign f2424_rst = rst;
  // Bindings to f2424

  // f2426
  logic [0:0] f2426_wen;
  logic [31:0] f2426_wdata;
  logic [0:0] f2426_clk;
  logic [0:0] f2426_rst;
  logic [31:0] f2426_rdata;
  sr_buffer_32_1 f2426(.wen(f2426_wen), .wdata(f2426_wdata), .clk(f2426_clk), .rst(f2426_rst), .rdata(f2426_rdata));
  assign f2426_clk = clk;
  assign f2426_rst = rst;
  // Bindings to f2426

  // f2428
  logic [0:0] f2428_wen;
  logic [31:0] f2428_wdata;
  logic [0:0] f2428_clk;
  logic [0:0] f2428_rst;
  logic [31:0] f2428_rdata;
  sr_buffer_32_1 f2428(.wen(f2428_wen), .wdata(f2428_wdata), .clk(f2428_clk), .rst(f2428_rst), .rdata(f2428_rdata));
  assign f2428_clk = clk;
  assign f2428_rst = rst;
  // Bindings to f2428

  // f2430
  logic [0:0] f2430_wen;
  logic [31:0] f2430_wdata;
  logic [0:0] f2430_clk;
  logic [0:0] f2430_rst;
  logic [31:0] f2430_rdata;
  sr_buffer_32_1 f2430(.wen(f2430_wen), .wdata(f2430_wdata), .clk(f2430_clk), .rst(f2430_rst), .rdata(f2430_rdata));
  assign f2430_clk = clk;
  assign f2430_rst = rst;
  // Bindings to f2430

  // f2432
  logic [0:0] f2432_wen;
  logic [31:0] f2432_wdata;
  logic [0:0] f2432_clk;
  logic [0:0] f2432_rst;
  logic [31:0] f2432_rdata;
  sr_buffer_32_1 f2432(.wen(f2432_wen), .wdata(f2432_wdata), .clk(f2432_clk), .rst(f2432_rst), .rdata(f2432_rdata));
  assign f2432_clk = clk;
  assign f2432_rst = rst;
  // Bindings to f2432

  // f2434
  logic [0:0] f2434_wen;
  logic [31:0] f2434_wdata;
  logic [0:0] f2434_clk;
  logic [0:0] f2434_rst;
  logic [31:0] f2434_rdata;
  sr_buffer_32_1 f2434(.wen(f2434_wen), .wdata(f2434_wdata), .clk(f2434_clk), .rst(f2434_rst), .rdata(f2434_rdata));
  assign f2434_clk = clk;
  assign f2434_rst = rst;
  // Bindings to f2434

  // f2436
  logic [0:0] f2436_wen;
  logic [31:0] f2436_wdata;
  logic [0:0] f2436_clk;
  logic [0:0] f2436_rst;
  logic [31:0] f2436_rdata;
  sr_buffer_32_1 f2436(.wen(f2436_wen), .wdata(f2436_wdata), .clk(f2436_clk), .rst(f2436_rst), .rdata(f2436_rdata));
  assign f2436_clk = clk;
  assign f2436_rst = rst;
  // Bindings to f2436

  // f2438
  logic [0:0] f2438_wen;
  logic [31:0] f2438_wdata;
  logic [0:0] f2438_clk;
  logic [0:0] f2438_rst;
  logic [31:0] f2438_rdata;
  sr_buffer_32_1 f2438(.wen(f2438_wen), .wdata(f2438_wdata), .clk(f2438_clk), .rst(f2438_rst), .rdata(f2438_rdata));
  assign f2438_clk = clk;
  assign f2438_rst = rst;
  // Bindings to f2438

  // f2440
  logic [0:0] f2440_wen;
  logic [31:0] f2440_wdata;
  logic [0:0] f2440_clk;
  logic [0:0] f2440_rst;
  logic [31:0] f2440_rdata;
  sr_buffer_32_1 f2440(.wen(f2440_wen), .wdata(f2440_wdata), .clk(f2440_clk), .rst(f2440_rst), .rdata(f2440_rdata));
  assign f2440_clk = clk;
  assign f2440_rst = rst;
  // Bindings to f2440

  // f2442
  logic [0:0] f2442_wen;
  logic [31:0] f2442_wdata;
  logic [0:0] f2442_clk;
  logic [0:0] f2442_rst;
  logic [31:0] f2442_rdata;
  sr_buffer_32_1 f2442(.wen(f2442_wen), .wdata(f2442_wdata), .clk(f2442_clk), .rst(f2442_rst), .rdata(f2442_rdata));
  assign f2442_clk = clk;
  assign f2442_rst = rst;
  // Bindings to f2442

  // f2444
  logic [0:0] f2444_wen;
  logic [31:0] f2444_wdata;
  logic [0:0] f2444_clk;
  logic [0:0] f2444_rst;
  logic [31:0] f2444_rdata;
  sr_buffer_32_1 f2444(.wen(f2444_wen), .wdata(f2444_wdata), .clk(f2444_clk), .rst(f2444_rst), .rdata(f2444_rdata));
  assign f2444_clk = clk;
  assign f2444_rst = rst;
  // Bindings to f2444

  // f2446
  logic [0:0] f2446_wen;
  logic [31:0] f2446_wdata;
  logic [0:0] f2446_clk;
  logic [0:0] f2446_rst;
  logic [31:0] f2446_rdata;
  sr_buffer_32_1 f2446(.wen(f2446_wen), .wdata(f2446_wdata), .clk(f2446_clk), .rst(f2446_rst), .rdata(f2446_rdata));
  assign f2446_clk = clk;
  assign f2446_rst = rst;
  // Bindings to f2446

  // f2448
  logic [0:0] f2448_wen;
  logic [31:0] f2448_wdata;
  logic [0:0] f2448_clk;
  logic [0:0] f2448_rst;
  logic [31:0] f2448_rdata;
  sr_buffer_32_1 f2448(.wen(f2448_wen), .wdata(f2448_wdata), .clk(f2448_clk), .rst(f2448_rst), .rdata(f2448_rdata));
  assign f2448_clk = clk;
  assign f2448_rst = rst;
  // Bindings to f2448

  // f2450
  logic [0:0] f2450_wen;
  logic [31:0] f2450_wdata;
  logic [0:0] f2450_clk;
  logic [0:0] f2450_rst;
  logic [31:0] f2450_rdata;
  sr_buffer_32_1 f2450(.wen(f2450_wen), .wdata(f2450_wdata), .clk(f2450_clk), .rst(f2450_rst), .rdata(f2450_rdata));
  assign f2450_clk = clk;
  assign f2450_rst = rst;
  // Bindings to f2450

  // f2452
  logic [0:0] f2452_wen;
  logic [31:0] f2452_wdata;
  logic [0:0] f2452_clk;
  logic [0:0] f2452_rst;
  logic [31:0] f2452_rdata;
  sr_buffer_32_1 f2452(.wen(f2452_wen), .wdata(f2452_wdata), .clk(f2452_clk), .rst(f2452_rst), .rdata(f2452_rdata));
  assign f2452_clk = clk;
  assign f2452_rst = rst;
  // Bindings to f2452

  // f2454
  logic [0:0] f2454_wen;
  logic [31:0] f2454_wdata;
  logic [0:0] f2454_clk;
  logic [0:0] f2454_rst;
  logic [31:0] f2454_rdata;
  sr_buffer_32_1 f2454(.wen(f2454_wen), .wdata(f2454_wdata), .clk(f2454_clk), .rst(f2454_rst), .rdata(f2454_rdata));
  assign f2454_clk = clk;
  assign f2454_rst = rst;
  // Bindings to f2454

  // f2456
  logic [0:0] f2456_wen;
  logic [31:0] f2456_wdata;
  logic [0:0] f2456_clk;
  logic [0:0] f2456_rst;
  logic [31:0] f2456_rdata;
  sr_buffer_32_1 f2456(.wen(f2456_wen), .wdata(f2456_wdata), .clk(f2456_clk), .rst(f2456_rst), .rdata(f2456_rdata));
  assign f2456_clk = clk;
  assign f2456_rst = rst;
  // Bindings to f2456

  // f2458
  logic [0:0] f2458_wen;
  logic [31:0] f2458_wdata;
  logic [0:0] f2458_clk;
  logic [0:0] f2458_rst;
  logic [31:0] f2458_rdata;
  sr_buffer_32_1 f2458(.wen(f2458_wen), .wdata(f2458_wdata), .clk(f2458_clk), .rst(f2458_rst), .rdata(f2458_rdata));
  assign f2458_clk = clk;
  assign f2458_rst = rst;
  // Bindings to f2458

  // f2460
  logic [0:0] f2460_wen;
  logic [31:0] f2460_wdata;
  logic [0:0] f2460_clk;
  logic [0:0] f2460_rst;
  logic [31:0] f2460_rdata;
  sr_buffer_32_1 f2460(.wen(f2460_wen), .wdata(f2460_wdata), .clk(f2460_clk), .rst(f2460_rst), .rdata(f2460_rdata));
  assign f2460_clk = clk;
  assign f2460_rst = rst;
  // Bindings to f2460

  // f2462
  logic [0:0] f2462_wen;
  logic [31:0] f2462_wdata;
  logic [0:0] f2462_clk;
  logic [0:0] f2462_rst;
  logic [31:0] f2462_rdata;
  sr_buffer_32_1 f2462(.wen(f2462_wen), .wdata(f2462_wdata), .clk(f2462_clk), .rst(f2462_rst), .rdata(f2462_rdata));
  assign f2462_clk = clk;
  assign f2462_rst = rst;
  // Bindings to f2462

  // f2464
  logic [0:0] f2464_wen;
  logic [31:0] f2464_wdata;
  logic [0:0] f2464_clk;
  logic [0:0] f2464_rst;
  logic [31:0] f2464_rdata;
  sr_buffer_32_1 f2464(.wen(f2464_wen), .wdata(f2464_wdata), .clk(f2464_clk), .rst(f2464_rst), .rdata(f2464_rdata));
  assign f2464_clk = clk;
  assign f2464_rst = rst;
  // Bindings to f2464

  // f2466
  logic [0:0] f2466_wen;
  logic [31:0] f2466_wdata;
  logic [0:0] f2466_clk;
  logic [0:0] f2466_rst;
  logic [31:0] f2466_rdata;
  sr_buffer_32_1 f2466(.wen(f2466_wen), .wdata(f2466_wdata), .clk(f2466_clk), .rst(f2466_rst), .rdata(f2466_rdata));
  assign f2466_clk = clk;
  assign f2466_rst = rst;
  // Bindings to f2466

  // f2468
  logic [0:0] f2468_wen;
  logic [31:0] f2468_wdata;
  logic [0:0] f2468_clk;
  logic [0:0] f2468_rst;
  logic [31:0] f2468_rdata;
  sr_buffer_32_1 f2468(.wen(f2468_wen), .wdata(f2468_wdata), .clk(f2468_clk), .rst(f2468_rst), .rdata(f2468_rdata));
  assign f2468_clk = clk;
  assign f2468_rst = rst;
  // Bindings to f2468

  // f2470
  logic [0:0] f2470_wen;
  logic [31:0] f2470_wdata;
  logic [0:0] f2470_clk;
  logic [0:0] f2470_rst;
  logic [31:0] f2470_rdata;
  sr_buffer_32_1 f2470(.wen(f2470_wen), .wdata(f2470_wdata), .clk(f2470_clk), .rst(f2470_rst), .rdata(f2470_rdata));
  assign f2470_clk = clk;
  assign f2470_rst = rst;
  // Bindings to f2470

  // f2472
  logic [0:0] f2472_wen;
  logic [31:0] f2472_wdata;
  logic [0:0] f2472_clk;
  logic [0:0] f2472_rst;
  logic [31:0] f2472_rdata;
  sr_buffer_32_1 f2472(.wen(f2472_wen), .wdata(f2472_wdata), .clk(f2472_clk), .rst(f2472_rst), .rdata(f2472_rdata));
  assign f2472_clk = clk;
  assign f2472_rst = rst;
  // Bindings to f2472

  // f2474
  logic [0:0] f2474_wen;
  logic [31:0] f2474_wdata;
  logic [0:0] f2474_clk;
  logic [0:0] f2474_rst;
  logic [31:0] f2474_rdata;
  sr_buffer_32_1 f2474(.wen(f2474_wen), .wdata(f2474_wdata), .clk(f2474_clk), .rst(f2474_rst), .rdata(f2474_rdata));
  assign f2474_clk = clk;
  assign f2474_rst = rst;
  // Bindings to f2474

  // f2476
  logic [0:0] f2476_wen;
  logic [31:0] f2476_wdata;
  logic [0:0] f2476_clk;
  logic [0:0] f2476_rst;
  logic [31:0] f2476_rdata;
  sr_buffer_32_1 f2476(.wen(f2476_wen), .wdata(f2476_wdata), .clk(f2476_clk), .rst(f2476_rst), .rdata(f2476_rdata));
  assign f2476_clk = clk;
  assign f2476_rst = rst;
  // Bindings to f2476

  // f2478
  logic [0:0] f2478_wen;
  logic [31:0] f2478_wdata;
  logic [0:0] f2478_clk;
  logic [0:0] f2478_rst;
  logic [31:0] f2478_rdata;
  sr_buffer_32_1 f2478(.wen(f2478_wen), .wdata(f2478_wdata), .clk(f2478_clk), .rst(f2478_rst), .rdata(f2478_rdata));
  assign f2478_clk = clk;
  assign f2478_rst = rst;
  // Bindings to f2478

  // f2480
  logic [0:0] f2480_wen;
  logic [31:0] f2480_wdata;
  logic [0:0] f2480_clk;
  logic [0:0] f2480_rst;
  logic [31:0] f2480_rdata;
  sr_buffer_32_1 f2480(.wen(f2480_wen), .wdata(f2480_wdata), .clk(f2480_clk), .rst(f2480_rst), .rdata(f2480_rdata));
  assign f2480_clk = clk;
  assign f2480_rst = rst;
  // Bindings to f2480

  // f2482
  logic [0:0] f2482_wen;
  logic [31:0] f2482_wdata;
  logic [0:0] f2482_clk;
  logic [0:0] f2482_rst;
  logic [31:0] f2482_rdata;
  sr_buffer_32_1 f2482(.wen(f2482_wen), .wdata(f2482_wdata), .clk(f2482_clk), .rst(f2482_rst), .rdata(f2482_rdata));
  assign f2482_clk = clk;
  assign f2482_rst = rst;
  // Bindings to f2482

  // f2484
  logic [0:0] f2484_wen;
  logic [31:0] f2484_wdata;
  logic [0:0] f2484_clk;
  logic [0:0] f2484_rst;
  logic [31:0] f2484_rdata;
  sr_buffer_32_1 f2484(.wen(f2484_wen), .wdata(f2484_wdata), .clk(f2484_clk), .rst(f2484_rst), .rdata(f2484_rdata));
  assign f2484_clk = clk;
  assign f2484_rst = rst;
  // Bindings to f2484

  // f2486
  logic [0:0] f2486_wen;
  logic [31:0] f2486_wdata;
  logic [0:0] f2486_clk;
  logic [0:0] f2486_rst;
  logic [31:0] f2486_rdata;
  sr_buffer_32_1 f2486(.wen(f2486_wen), .wdata(f2486_wdata), .clk(f2486_clk), .rst(f2486_rst), .rdata(f2486_rdata));
  assign f2486_clk = clk;
  assign f2486_rst = rst;
  // Bindings to f2486

  // f2488
  logic [0:0] f2488_wen;
  logic [31:0] f2488_wdata;
  logic [0:0] f2488_clk;
  logic [0:0] f2488_rst;
  logic [31:0] f2488_rdata;
  sr_buffer_32_1 f2488(.wen(f2488_wen), .wdata(f2488_wdata), .clk(f2488_clk), .rst(f2488_rst), .rdata(f2488_rdata));
  assign f2488_clk = clk;
  assign f2488_rst = rst;
  // Bindings to f2488

  // f2490
  logic [0:0] f2490_wen;
  logic [31:0] f2490_wdata;
  logic [0:0] f2490_clk;
  logic [0:0] f2490_rst;
  logic [31:0] f2490_rdata;
  sr_buffer_32_1 f2490(.wen(f2490_wen), .wdata(f2490_wdata), .clk(f2490_clk), .rst(f2490_rst), .rdata(f2490_rdata));
  assign f2490_clk = clk;
  assign f2490_rst = rst;
  // Bindings to f2490

  // f2492
  logic [0:0] f2492_wen;
  logic [31:0] f2492_wdata;
  logic [0:0] f2492_clk;
  logic [0:0] f2492_rst;
  logic [31:0] f2492_rdata;
  sr_buffer_32_1 f2492(.wen(f2492_wen), .wdata(f2492_wdata), .clk(f2492_clk), .rst(f2492_rst), .rdata(f2492_rdata));
  assign f2492_clk = clk;
  assign f2492_rst = rst;
  // Bindings to f2492

  // f2494
  logic [0:0] f2494_wen;
  logic [31:0] f2494_wdata;
  logic [0:0] f2494_clk;
  logic [0:0] f2494_rst;
  logic [31:0] f2494_rdata;
  sr_buffer_32_1 f2494(.wen(f2494_wen), .wdata(f2494_wdata), .clk(f2494_clk), .rst(f2494_rst), .rdata(f2494_rdata));
  assign f2494_clk = clk;
  assign f2494_rst = rst;
  // Bindings to f2494

  // f2496
  logic [0:0] f2496_wen;
  logic [31:0] f2496_wdata;
  logic [0:0] f2496_clk;
  logic [0:0] f2496_rst;
  logic [31:0] f2496_rdata;
  sr_buffer_32_1 f2496(.wen(f2496_wen), .wdata(f2496_wdata), .clk(f2496_clk), .rst(f2496_rst), .rdata(f2496_rdata));
  assign f2496_clk = clk;
  assign f2496_rst = rst;
  // Bindings to f2496

  // f2498
  logic [0:0] f2498_wen;
  logic [31:0] f2498_wdata;
  logic [0:0] f2498_clk;
  logic [0:0] f2498_rst;
  logic [31:0] f2498_rdata;
  sr_buffer_32_1 f2498(.wen(f2498_wen), .wdata(f2498_wdata), .clk(f2498_clk), .rst(f2498_rst), .rdata(f2498_rdata));
  assign f2498_clk = clk;
  assign f2498_rst = rst;
  // Bindings to f2498

  // f2500
  logic [0:0] f2500_wen;
  logic [31:0] f2500_wdata;
  logic [0:0] f2500_clk;
  logic [0:0] f2500_rst;
  logic [31:0] f2500_rdata;
  sr_buffer_32_1 f2500(.wen(f2500_wen), .wdata(f2500_wdata), .clk(f2500_clk), .rst(f2500_rst), .rdata(f2500_rdata));
  assign f2500_clk = clk;
  assign f2500_rst = rst;
  // Bindings to f2500

  // f2502
  logic [0:0] f2502_wen;
  logic [31:0] f2502_wdata;
  logic [0:0] f2502_clk;
  logic [0:0] f2502_rst;
  logic [31:0] f2502_rdata;
  sr_buffer_32_1 f2502(.wen(f2502_wen), .wdata(f2502_wdata), .clk(f2502_clk), .rst(f2502_rst), .rdata(f2502_rdata));
  assign f2502_clk = clk;
  assign f2502_rst = rst;
  // Bindings to f2502

  // f2504
  logic [0:0] f2504_wen;
  logic [31:0] f2504_wdata;
  logic [0:0] f2504_clk;
  logic [0:0] f2504_rst;
  logic [31:0] f2504_rdata;
  sr_buffer_32_1 f2504(.wen(f2504_wen), .wdata(f2504_wdata), .clk(f2504_clk), .rst(f2504_rst), .rdata(f2504_rdata));
  assign f2504_clk = clk;
  assign f2504_rst = rst;
  // Bindings to f2504

  // f2506
  logic [0:0] f2506_wen;
  logic [31:0] f2506_wdata;
  logic [0:0] f2506_clk;
  logic [0:0] f2506_rst;
  logic [31:0] f2506_rdata;
  sr_buffer_32_1 f2506(.wen(f2506_wen), .wdata(f2506_wdata), .clk(f2506_clk), .rst(f2506_rst), .rdata(f2506_rdata));
  assign f2506_clk = clk;
  assign f2506_rst = rst;
  // Bindings to f2506

  // f2508
  logic [0:0] f2508_wen;
  logic [31:0] f2508_wdata;
  logic [0:0] f2508_clk;
  logic [0:0] f2508_rst;
  logic [31:0] f2508_rdata;
  sr_buffer_32_1 f2508(.wen(f2508_wen), .wdata(f2508_wdata), .clk(f2508_clk), .rst(f2508_rst), .rdata(f2508_rdata));
  assign f2508_clk = clk;
  assign f2508_rst = rst;
  // Bindings to f2508

  // f2510
  logic [0:0] f2510_wen;
  logic [31:0] f2510_wdata;
  logic [0:0] f2510_clk;
  logic [0:0] f2510_rst;
  logic [31:0] f2510_rdata;
  sr_buffer_32_1 f2510(.wen(f2510_wen), .wdata(f2510_wdata), .clk(f2510_clk), .rst(f2510_rst), .rdata(f2510_rdata));
  assign f2510_clk = clk;
  assign f2510_rst = rst;
  // Bindings to f2510

  // f2512
  logic [0:0] f2512_wen;
  logic [31:0] f2512_wdata;
  logic [0:0] f2512_clk;
  logic [0:0] f2512_rst;
  logic [31:0] f2512_rdata;
  sr_buffer_32_1 f2512(.wen(f2512_wen), .wdata(f2512_wdata), .clk(f2512_clk), .rst(f2512_rst), .rdata(f2512_rdata));
  assign f2512_clk = clk;
  assign f2512_rst = rst;
  // Bindings to f2512

  // f2514
  logic [0:0] f2514_wen;
  logic [31:0] f2514_wdata;
  logic [0:0] f2514_clk;
  logic [0:0] f2514_rst;
  logic [31:0] f2514_rdata;
  sr_buffer_32_1 f2514(.wen(f2514_wen), .wdata(f2514_wdata), .clk(f2514_clk), .rst(f2514_rst), .rdata(f2514_rdata));
  assign f2514_clk = clk;
  assign f2514_rst = rst;
  // Bindings to f2514

  // f2516
  logic [0:0] f2516_wen;
  logic [31:0] f2516_wdata;
  logic [0:0] f2516_clk;
  logic [0:0] f2516_rst;
  logic [31:0] f2516_rdata;
  sr_buffer_32_1 f2516(.wen(f2516_wen), .wdata(f2516_wdata), .clk(f2516_clk), .rst(f2516_rst), .rdata(f2516_rdata));
  assign f2516_clk = clk;
  assign f2516_rst = rst;
  // Bindings to f2516

  // f2518
  logic [0:0] f2518_wen;
  logic [31:0] f2518_wdata;
  logic [0:0] f2518_clk;
  logic [0:0] f2518_rst;
  logic [31:0] f2518_rdata;
  sr_buffer_32_1 f2518(.wen(f2518_wen), .wdata(f2518_wdata), .clk(f2518_clk), .rst(f2518_rst), .rdata(f2518_rdata));
  assign f2518_clk = clk;
  assign f2518_rst = rst;
  // Bindings to f2518

  // f2520
  logic [0:0] f2520_wen;
  logic [31:0] f2520_wdata;
  logic [0:0] f2520_clk;
  logic [0:0] f2520_rst;
  logic [31:0] f2520_rdata;
  sr_buffer_32_1 f2520(.wen(f2520_wen), .wdata(f2520_wdata), .clk(f2520_clk), .rst(f2520_rst), .rdata(f2520_rdata));
  assign f2520_clk = clk;
  assign f2520_rst = rst;
  // Bindings to f2520

  // f2522
  logic [0:0] f2522_wen;
  logic [31:0] f2522_wdata;
  logic [0:0] f2522_clk;
  logic [0:0] f2522_rst;
  logic [31:0] f2522_rdata;
  sr_buffer_32_1 f2522(.wen(f2522_wen), .wdata(f2522_wdata), .clk(f2522_clk), .rst(f2522_rst), .rdata(f2522_rdata));
  assign f2522_clk = clk;
  assign f2522_rst = rst;
  // Bindings to f2522

  // f2524
  logic [0:0] f2524_wen;
  logic [31:0] f2524_wdata;
  logic [0:0] f2524_clk;
  logic [0:0] f2524_rst;
  logic [31:0] f2524_rdata;
  sr_buffer_32_1 f2524(.wen(f2524_wen), .wdata(f2524_wdata), .clk(f2524_clk), .rst(f2524_rst), .rdata(f2524_rdata));
  assign f2524_clk = clk;
  assign f2524_rst = rst;
  // Bindings to f2524

  // f2526
  logic [0:0] f2526_wen;
  logic [31:0] f2526_wdata;
  logic [0:0] f2526_clk;
  logic [0:0] f2526_rst;
  logic [31:0] f2526_rdata;
  sr_buffer_32_1 f2526(.wen(f2526_wen), .wdata(f2526_wdata), .clk(f2526_clk), .rst(f2526_rst), .rdata(f2526_rdata));
  assign f2526_clk = clk;
  assign f2526_rst = rst;
  // Bindings to f2526

  // f2528
  logic [0:0] f2528_wen;
  logic [31:0] f2528_wdata;
  logic [0:0] f2528_clk;
  logic [0:0] f2528_rst;
  logic [31:0] f2528_rdata;
  sr_buffer_32_1 f2528(.wen(f2528_wen), .wdata(f2528_wdata), .clk(f2528_clk), .rst(f2528_rst), .rdata(f2528_rdata));
  assign f2528_clk = clk;
  assign f2528_rst = rst;
  // Bindings to f2528

  // f2530
  logic [0:0] f2530_wen;
  logic [31:0] f2530_wdata;
  logic [0:0] f2530_clk;
  logic [0:0] f2530_rst;
  logic [31:0] f2530_rdata;
  sr_buffer_32_1 f2530(.wen(f2530_wen), .wdata(f2530_wdata), .clk(f2530_clk), .rst(f2530_rst), .rdata(f2530_rdata));
  assign f2530_clk = clk;
  assign f2530_rst = rst;
  // Bindings to f2530

  // f772
  logic [0:0] f772_wen;
  logic [31:0] f772_wdata;
  logic [0:0] f772_clk;
  logic [0:0] f772_rst;
  logic [31:0] f772_rdata;
  sr_buffer_32_1 f772(.wen(f772_wen), .wdata(f772_wdata), .clk(f772_clk), .rst(f772_rst), .rdata(f772_rdata));
  assign f772_clk = clk;
  assign f772_rst = rst;
  // Bindings to f772

  // f774
  logic [0:0] f774_wen;
  logic [31:0] f774_wdata;
  logic [0:0] f774_clk;
  logic [0:0] f774_rst;
  logic [31:0] f774_rdata;
  sr_buffer_32_1 f774(.wen(f774_wen), .wdata(f774_wdata), .clk(f774_clk), .rst(f774_rst), .rdata(f774_rdata));
  assign f774_clk = clk;
  assign f774_rst = rst;
  // Bindings to f774

  // f776
  logic [0:0] f776_wen;
  logic [31:0] f776_wdata;
  logic [0:0] f776_clk;
  logic [0:0] f776_rst;
  logic [31:0] f776_rdata;
  sr_buffer_32_1 f776(.wen(f776_wen), .wdata(f776_wdata), .clk(f776_clk), .rst(f776_rst), .rdata(f776_rdata));
  assign f776_clk = clk;
  assign f776_rst = rst;
  // Bindings to f776

  // f778
  logic [0:0] f778_wen;
  logic [31:0] f778_wdata;
  logic [0:0] f778_clk;
  logic [0:0] f778_rst;
  logic [31:0] f778_rdata;
  sr_buffer_32_1 f778(.wen(f778_wen), .wdata(f778_wdata), .clk(f778_clk), .rst(f778_rst), .rdata(f778_rdata));
  assign f778_clk = clk;
  assign f778_rst = rst;
  // Bindings to f778

  // f780
  logic [0:0] f780_wen;
  logic [31:0] f780_wdata;
  logic [0:0] f780_clk;
  logic [0:0] f780_rst;
  logic [31:0] f780_rdata;
  sr_buffer_32_1 f780(.wen(f780_wen), .wdata(f780_wdata), .clk(f780_clk), .rst(f780_rst), .rdata(f780_rdata));
  assign f780_clk = clk;
  assign f780_rst = rst;
  // Bindings to f780

  // f782
  logic [0:0] f782_wen;
  logic [31:0] f782_wdata;
  logic [0:0] f782_clk;
  logic [0:0] f782_rst;
  logic [31:0] f782_rdata;
  sr_buffer_32_1 f782(.wen(f782_wen), .wdata(f782_wdata), .clk(f782_clk), .rst(f782_rst), .rdata(f782_rdata));
  assign f782_clk = clk;
  assign f782_rst = rst;
  // Bindings to f782

  // f784
  logic [0:0] f784_wen;
  logic [31:0] f784_wdata;
  logic [0:0] f784_clk;
  logic [0:0] f784_rst;
  logic [31:0] f784_rdata;
  sr_buffer_32_1 f784(.wen(f784_wen), .wdata(f784_wdata), .clk(f784_clk), .rst(f784_rst), .rdata(f784_rdata));
  assign f784_clk = clk;
  assign f784_rst = rst;
  // Bindings to f784

  // f786
  logic [0:0] f786_wen;
  logic [31:0] f786_wdata;
  logic [0:0] f786_clk;
  logic [0:0] f786_rst;
  logic [31:0] f786_rdata;
  sr_buffer_32_1 f786(.wen(f786_wen), .wdata(f786_wdata), .clk(f786_clk), .rst(f786_rst), .rdata(f786_rdata));
  assign f786_clk = clk;
  assign f786_rst = rst;
  // Bindings to f786

  // f788
  logic [0:0] f788_wen;
  logic [31:0] f788_wdata;
  logic [0:0] f788_clk;
  logic [0:0] f788_rst;
  logic [31:0] f788_rdata;
  sr_buffer_32_1 f788(.wen(f788_wen), .wdata(f788_wdata), .clk(f788_clk), .rst(f788_rst), .rdata(f788_rdata));
  assign f788_clk = clk;
  assign f788_rst = rst;
  // Bindings to f788

  // f790
  logic [0:0] f790_wen;
  logic [31:0] f790_wdata;
  logic [0:0] f790_clk;
  logic [0:0] f790_rst;
  logic [31:0] f790_rdata;
  sr_buffer_32_1 f790(.wen(f790_wen), .wdata(f790_wdata), .clk(f790_clk), .rst(f790_rst), .rdata(f790_rdata));
  assign f790_clk = clk;
  assign f790_rst = rst;
  // Bindings to f790

  // f792
  logic [0:0] f792_wen;
  logic [31:0] f792_wdata;
  logic [0:0] f792_clk;
  logic [0:0] f792_rst;
  logic [31:0] f792_rdata;
  sr_buffer_32_1 f792(.wen(f792_wen), .wdata(f792_wdata), .clk(f792_clk), .rst(f792_rst), .rdata(f792_rdata));
  assign f792_clk = clk;
  assign f792_rst = rst;
  // Bindings to f792

  // f794
  logic [0:0] f794_wen;
  logic [31:0] f794_wdata;
  logic [0:0] f794_clk;
  logic [0:0] f794_rst;
  logic [31:0] f794_rdata;
  sr_buffer_32_1 f794(.wen(f794_wen), .wdata(f794_wdata), .clk(f794_clk), .rst(f794_rst), .rdata(f794_rdata));
  assign f794_clk = clk;
  assign f794_rst = rst;
  // Bindings to f794

  // f796
  logic [0:0] f796_wen;
  logic [31:0] f796_wdata;
  logic [0:0] f796_clk;
  logic [0:0] f796_rst;
  logic [31:0] f796_rdata;
  sr_buffer_32_1 f796(.wen(f796_wen), .wdata(f796_wdata), .clk(f796_clk), .rst(f796_rst), .rdata(f796_rdata));
  assign f796_clk = clk;
  assign f796_rst = rst;
  // Bindings to f796

  // f798
  logic [0:0] f798_wen;
  logic [31:0] f798_wdata;
  logic [0:0] f798_clk;
  logic [0:0] f798_rst;
  logic [31:0] f798_rdata;
  sr_buffer_32_1 f798(.wen(f798_wen), .wdata(f798_wdata), .clk(f798_clk), .rst(f798_rst), .rdata(f798_rdata));
  assign f798_clk = clk;
  assign f798_rst = rst;
  // Bindings to f798

  // f800
  logic [0:0] f800_wen;
  logic [31:0] f800_wdata;
  logic [0:0] f800_clk;
  logic [0:0] f800_rst;
  logic [31:0] f800_rdata;
  sr_buffer_32_1 f800(.wen(f800_wen), .wdata(f800_wdata), .clk(f800_clk), .rst(f800_rst), .rdata(f800_rdata));
  assign f800_clk = clk;
  assign f800_rst = rst;
  // Bindings to f800

  // f802
  logic [0:0] f802_wen;
  logic [31:0] f802_wdata;
  logic [0:0] f802_clk;
  logic [0:0] f802_rst;
  logic [31:0] f802_rdata;
  sr_buffer_32_1 f802(.wen(f802_wen), .wdata(f802_wdata), .clk(f802_clk), .rst(f802_rst), .rdata(f802_rdata));
  assign f802_clk = clk;
  assign f802_rst = rst;
  // Bindings to f802

  // f804
  logic [0:0] f804_wen;
  logic [31:0] f804_wdata;
  logic [0:0] f804_clk;
  logic [0:0] f804_rst;
  logic [31:0] f804_rdata;
  sr_buffer_32_1 f804(.wen(f804_wen), .wdata(f804_wdata), .clk(f804_clk), .rst(f804_rst), .rdata(f804_rdata));
  assign f804_clk = clk;
  assign f804_rst = rst;
  // Bindings to f804

  // f806
  logic [0:0] f806_wen;
  logic [31:0] f806_wdata;
  logic [0:0] f806_clk;
  logic [0:0] f806_rst;
  logic [31:0] f806_rdata;
  sr_buffer_32_1 f806(.wen(f806_wen), .wdata(f806_wdata), .clk(f806_clk), .rst(f806_rst), .rdata(f806_rdata));
  assign f806_clk = clk;
  assign f806_rst = rst;
  // Bindings to f806

  // f808
  logic [0:0] f808_wen;
  logic [31:0] f808_wdata;
  logic [0:0] f808_clk;
  logic [0:0] f808_rst;
  logic [31:0] f808_rdata;
  sr_buffer_32_1 f808(.wen(f808_wen), .wdata(f808_wdata), .clk(f808_clk), .rst(f808_rst), .rdata(f808_rdata));
  assign f808_clk = clk;
  assign f808_rst = rst;
  // Bindings to f808

  // f810
  logic [0:0] f810_wen;
  logic [31:0] f810_wdata;
  logic [0:0] f810_clk;
  logic [0:0] f810_rst;
  logic [31:0] f810_rdata;
  sr_buffer_32_1 f810(.wen(f810_wen), .wdata(f810_wdata), .clk(f810_clk), .rst(f810_rst), .rdata(f810_rdata));
  assign f810_clk = clk;
  assign f810_rst = rst;
  // Bindings to f810

  // f812
  logic [0:0] f812_wen;
  logic [31:0] f812_wdata;
  logic [0:0] f812_clk;
  logic [0:0] f812_rst;
  logic [31:0] f812_rdata;
  sr_buffer_32_1 f812(.wen(f812_wen), .wdata(f812_wdata), .clk(f812_clk), .rst(f812_rst), .rdata(f812_rdata));
  assign f812_clk = clk;
  assign f812_rst = rst;
  // Bindings to f812

  // f814
  logic [0:0] f814_wen;
  logic [31:0] f814_wdata;
  logic [0:0] f814_clk;
  logic [0:0] f814_rst;
  logic [31:0] f814_rdata;
  sr_buffer_32_1 f814(.wen(f814_wen), .wdata(f814_wdata), .clk(f814_clk), .rst(f814_rst), .rdata(f814_rdata));
  assign f814_clk = clk;
  assign f814_rst = rst;
  // Bindings to f814

  // f816
  logic [0:0] f816_wen;
  logic [31:0] f816_wdata;
  logic [0:0] f816_clk;
  logic [0:0] f816_rst;
  logic [31:0] f816_rdata;
  sr_buffer_32_1 f816(.wen(f816_wen), .wdata(f816_wdata), .clk(f816_clk), .rst(f816_rst), .rdata(f816_rdata));
  assign f816_clk = clk;
  assign f816_rst = rst;
  // Bindings to f816

  // f818
  logic [0:0] f818_wen;
  logic [31:0] f818_wdata;
  logic [0:0] f818_clk;
  logic [0:0] f818_rst;
  logic [31:0] f818_rdata;
  sr_buffer_32_1 f818(.wen(f818_wen), .wdata(f818_wdata), .clk(f818_clk), .rst(f818_rst), .rdata(f818_rdata));
  assign f818_clk = clk;
  assign f818_rst = rst;
  // Bindings to f818

  // f820
  logic [0:0] f820_wen;
  logic [31:0] f820_wdata;
  logic [0:0] f820_clk;
  logic [0:0] f820_rst;
  logic [31:0] f820_rdata;
  sr_buffer_32_1 f820(.wen(f820_wen), .wdata(f820_wdata), .clk(f820_clk), .rst(f820_rst), .rdata(f820_rdata));
  assign f820_clk = clk;
  assign f820_rst = rst;
  // Bindings to f820

  // f822
  logic [0:0] f822_wen;
  logic [31:0] f822_wdata;
  logic [0:0] f822_clk;
  logic [0:0] f822_rst;
  logic [31:0] f822_rdata;
  sr_buffer_32_1 f822(.wen(f822_wen), .wdata(f822_wdata), .clk(f822_clk), .rst(f822_rst), .rdata(f822_rdata));
  assign f822_clk = clk;
  assign f822_rst = rst;
  // Bindings to f822

  // f824
  logic [0:0] f824_wen;
  logic [31:0] f824_wdata;
  logic [0:0] f824_clk;
  logic [0:0] f824_rst;
  logic [31:0] f824_rdata;
  sr_buffer_32_1 f824(.wen(f824_wen), .wdata(f824_wdata), .clk(f824_clk), .rst(f824_rst), .rdata(f824_rdata));
  assign f824_clk = clk;
  assign f824_rst = rst;
  // Bindings to f824

  // f826
  logic [0:0] f826_wen;
  logic [31:0] f826_wdata;
  logic [0:0] f826_clk;
  logic [0:0] f826_rst;
  logic [31:0] f826_rdata;
  sr_buffer_32_1 f826(.wen(f826_wen), .wdata(f826_wdata), .clk(f826_clk), .rst(f826_rst), .rdata(f826_rdata));
  assign f826_clk = clk;
  assign f826_rst = rst;
  // Bindings to f826

  // f828
  logic [0:0] f828_wen;
  logic [31:0] f828_wdata;
  logic [0:0] f828_clk;
  logic [0:0] f828_rst;
  logic [31:0] f828_rdata;
  sr_buffer_32_1 f828(.wen(f828_wen), .wdata(f828_wdata), .clk(f828_clk), .rst(f828_rst), .rdata(f828_rdata));
  assign f828_clk = clk;
  assign f828_rst = rst;
  // Bindings to f828

  // f830
  logic [0:0] f830_wen;
  logic [31:0] f830_wdata;
  logic [0:0] f830_clk;
  logic [0:0] f830_rst;
  logic [31:0] f830_rdata;
  sr_buffer_32_1 f830(.wen(f830_wen), .wdata(f830_wdata), .clk(f830_clk), .rst(f830_rst), .rdata(f830_rdata));
  assign f830_clk = clk;
  assign f830_rst = rst;
  // Bindings to f830

  // f832
  logic [0:0] f832_wen;
  logic [31:0] f832_wdata;
  logic [0:0] f832_clk;
  logic [0:0] f832_rst;
  logic [31:0] f832_rdata;
  sr_buffer_32_1 f832(.wen(f832_wen), .wdata(f832_wdata), .clk(f832_clk), .rst(f832_rst), .rdata(f832_rdata));
  assign f832_clk = clk;
  assign f832_rst = rst;
  // Bindings to f832

  // f834
  logic [0:0] f834_wen;
  logic [31:0] f834_wdata;
  logic [0:0] f834_clk;
  logic [0:0] f834_rst;
  logic [31:0] f834_rdata;
  sr_buffer_32_1 f834(.wen(f834_wen), .wdata(f834_wdata), .clk(f834_clk), .rst(f834_rst), .rdata(f834_rdata));
  assign f834_clk = clk;
  assign f834_rst = rst;
  // Bindings to f834

  // f836
  logic [0:0] f836_wen;
  logic [31:0] f836_wdata;
  logic [0:0] f836_clk;
  logic [0:0] f836_rst;
  logic [31:0] f836_rdata;
  sr_buffer_32_1 f836(.wen(f836_wen), .wdata(f836_wdata), .clk(f836_clk), .rst(f836_rst), .rdata(f836_rdata));
  assign f836_clk = clk;
  assign f836_rst = rst;
  // Bindings to f836

  // f838
  logic [0:0] f838_wen;
  logic [31:0] f838_wdata;
  logic [0:0] f838_clk;
  logic [0:0] f838_rst;
  logic [31:0] f838_rdata;
  sr_buffer_32_1 f838(.wen(f838_wen), .wdata(f838_wdata), .clk(f838_clk), .rst(f838_rst), .rdata(f838_rdata));
  assign f838_clk = clk;
  assign f838_rst = rst;
  // Bindings to f838

  // f840
  logic [0:0] f840_wen;
  logic [31:0] f840_wdata;
  logic [0:0] f840_clk;
  logic [0:0] f840_rst;
  logic [31:0] f840_rdata;
  sr_buffer_32_1 f840(.wen(f840_wen), .wdata(f840_wdata), .clk(f840_clk), .rst(f840_rst), .rdata(f840_rdata));
  assign f840_clk = clk;
  assign f840_rst = rst;
  // Bindings to f840

  // f842
  logic [0:0] f842_wen;
  logic [31:0] f842_wdata;
  logic [0:0] f842_clk;
  logic [0:0] f842_rst;
  logic [31:0] f842_rdata;
  sr_buffer_32_1 f842(.wen(f842_wen), .wdata(f842_wdata), .clk(f842_clk), .rst(f842_rst), .rdata(f842_rdata));
  assign f842_clk = clk;
  assign f842_rst = rst;
  // Bindings to f842

  // f844
  logic [0:0] f844_wen;
  logic [31:0] f844_wdata;
  logic [0:0] f844_clk;
  logic [0:0] f844_rst;
  logic [31:0] f844_rdata;
  sr_buffer_32_1 f844(.wen(f844_wen), .wdata(f844_wdata), .clk(f844_clk), .rst(f844_rst), .rdata(f844_rdata));
  assign f844_clk = clk;
  assign f844_rst = rst;
  // Bindings to f844

  // f846
  logic [0:0] f846_wen;
  logic [31:0] f846_wdata;
  logic [0:0] f846_clk;
  logic [0:0] f846_rst;
  logic [31:0] f846_rdata;
  sr_buffer_32_1 f846(.wen(f846_wen), .wdata(f846_wdata), .clk(f846_clk), .rst(f846_rst), .rdata(f846_rdata));
  assign f846_clk = clk;
  assign f846_rst = rst;
  // Bindings to f846

  // f848
  logic [0:0] f848_wen;
  logic [31:0] f848_wdata;
  logic [0:0] f848_clk;
  logic [0:0] f848_rst;
  logic [31:0] f848_rdata;
  sr_buffer_32_1 f848(.wen(f848_wen), .wdata(f848_wdata), .clk(f848_clk), .rst(f848_rst), .rdata(f848_rdata));
  assign f848_clk = clk;
  assign f848_rst = rst;
  // Bindings to f848

  // f850
  logic [0:0] f850_wen;
  logic [31:0] f850_wdata;
  logic [0:0] f850_clk;
  logic [0:0] f850_rst;
  logic [31:0] f850_rdata;
  sr_buffer_32_1 f850(.wen(f850_wen), .wdata(f850_wdata), .clk(f850_clk), .rst(f850_rst), .rdata(f850_rdata));
  assign f850_clk = clk;
  assign f850_rst = rst;
  // Bindings to f850

  // f852
  logic [0:0] f852_wen;
  logic [31:0] f852_wdata;
  logic [0:0] f852_clk;
  logic [0:0] f852_rst;
  logic [31:0] f852_rdata;
  sr_buffer_32_1 f852(.wen(f852_wen), .wdata(f852_wdata), .clk(f852_clk), .rst(f852_rst), .rdata(f852_rdata));
  assign f852_clk = clk;
  assign f852_rst = rst;
  // Bindings to f852

  // f854
  logic [0:0] f854_wen;
  logic [31:0] f854_wdata;
  logic [0:0] f854_clk;
  logic [0:0] f854_rst;
  logic [31:0] f854_rdata;
  sr_buffer_32_1 f854(.wen(f854_wen), .wdata(f854_wdata), .clk(f854_clk), .rst(f854_rst), .rdata(f854_rdata));
  assign f854_clk = clk;
  assign f854_rst = rst;
  // Bindings to f854

  // f856
  logic [0:0] f856_wen;
  logic [31:0] f856_wdata;
  logic [0:0] f856_clk;
  logic [0:0] f856_rst;
  logic [31:0] f856_rdata;
  sr_buffer_32_1 f856(.wen(f856_wen), .wdata(f856_wdata), .clk(f856_clk), .rst(f856_rst), .rdata(f856_rdata));
  assign f856_clk = clk;
  assign f856_rst = rst;
  // Bindings to f856

  // f858
  logic [0:0] f858_wen;
  logic [31:0] f858_wdata;
  logic [0:0] f858_clk;
  logic [0:0] f858_rst;
  logic [31:0] f858_rdata;
  sr_buffer_32_1 f858(.wen(f858_wen), .wdata(f858_wdata), .clk(f858_clk), .rst(f858_rst), .rdata(f858_rdata));
  assign f858_clk = clk;
  assign f858_rst = rst;
  // Bindings to f858

  // f860
  logic [0:0] f860_wen;
  logic [31:0] f860_wdata;
  logic [0:0] f860_clk;
  logic [0:0] f860_rst;
  logic [31:0] f860_rdata;
  sr_buffer_32_1 f860(.wen(f860_wen), .wdata(f860_wdata), .clk(f860_clk), .rst(f860_rst), .rdata(f860_rdata));
  assign f860_clk = clk;
  assign f860_rst = rst;
  // Bindings to f860

  // f862
  logic [0:0] f862_wen;
  logic [31:0] f862_wdata;
  logic [0:0] f862_clk;
  logic [0:0] f862_rst;
  logic [31:0] f862_rdata;
  sr_buffer_32_1 f862(.wen(f862_wen), .wdata(f862_wdata), .clk(f862_clk), .rst(f862_rst), .rdata(f862_rdata));
  assign f862_clk = clk;
  assign f862_rst = rst;
  // Bindings to f862

  // f864
  logic [0:0] f864_wen;
  logic [31:0] f864_wdata;
  logic [0:0] f864_clk;
  logic [0:0] f864_rst;
  logic [31:0] f864_rdata;
  sr_buffer_32_1 f864(.wen(f864_wen), .wdata(f864_wdata), .clk(f864_clk), .rst(f864_rst), .rdata(f864_rdata));
  assign f864_clk = clk;
  assign f864_rst = rst;
  // Bindings to f864

  // f866
  logic [0:0] f866_wen;
  logic [31:0] f866_wdata;
  logic [0:0] f866_clk;
  logic [0:0] f866_rst;
  logic [31:0] f866_rdata;
  sr_buffer_32_1 f866(.wen(f866_wen), .wdata(f866_wdata), .clk(f866_clk), .rst(f866_rst), .rdata(f866_rdata));
  assign f866_clk = clk;
  assign f866_rst = rst;
  // Bindings to f866

  // f868
  logic [0:0] f868_wen;
  logic [31:0] f868_wdata;
  logic [0:0] f868_clk;
  logic [0:0] f868_rst;
  logic [31:0] f868_rdata;
  sr_buffer_32_1 f868(.wen(f868_wen), .wdata(f868_wdata), .clk(f868_clk), .rst(f868_rst), .rdata(f868_rdata));
  assign f868_clk = clk;
  assign f868_rst = rst;
  // Bindings to f868

  // f870
  logic [0:0] f870_wen;
  logic [31:0] f870_wdata;
  logic [0:0] f870_clk;
  logic [0:0] f870_rst;
  logic [31:0] f870_rdata;
  sr_buffer_32_1 f870(.wen(f870_wen), .wdata(f870_wdata), .clk(f870_clk), .rst(f870_rst), .rdata(f870_rdata));
  assign f870_clk = clk;
  assign f870_rst = rst;
  // Bindings to f870

  // f872
  logic [0:0] f872_wen;
  logic [31:0] f872_wdata;
  logic [0:0] f872_clk;
  logic [0:0] f872_rst;
  logic [31:0] f872_rdata;
  sr_buffer_32_1 f872(.wen(f872_wen), .wdata(f872_wdata), .clk(f872_clk), .rst(f872_rst), .rdata(f872_rdata));
  assign f872_clk = clk;
  assign f872_rst = rst;
  // Bindings to f872

  // f874
  logic [0:0] f874_wen;
  logic [31:0] f874_wdata;
  logic [0:0] f874_clk;
  logic [0:0] f874_rst;
  logic [31:0] f874_rdata;
  sr_buffer_32_1 f874(.wen(f874_wen), .wdata(f874_wdata), .clk(f874_clk), .rst(f874_rst), .rdata(f874_rdata));
  assign f874_clk = clk;
  assign f874_rst = rst;
  // Bindings to f874

  // f876
  logic [0:0] f876_wen;
  logic [31:0] f876_wdata;
  logic [0:0] f876_clk;
  logic [0:0] f876_rst;
  logic [31:0] f876_rdata;
  sr_buffer_32_1 f876(.wen(f876_wen), .wdata(f876_wdata), .clk(f876_clk), .rst(f876_rst), .rdata(f876_rdata));
  assign f876_clk = clk;
  assign f876_rst = rst;
  // Bindings to f876

  // f878
  logic [0:0] f878_wen;
  logic [31:0] f878_wdata;
  logic [0:0] f878_clk;
  logic [0:0] f878_rst;
  logic [31:0] f878_rdata;
  sr_buffer_32_1 f878(.wen(f878_wen), .wdata(f878_wdata), .clk(f878_clk), .rst(f878_rst), .rdata(f878_rdata));
  assign f878_clk = clk;
  assign f878_rst = rst;
  // Bindings to f878

  // f880
  logic [0:0] f880_wen;
  logic [31:0] f880_wdata;
  logic [0:0] f880_clk;
  logic [0:0] f880_rst;
  logic [31:0] f880_rdata;
  sr_buffer_32_1 f880(.wen(f880_wen), .wdata(f880_wdata), .clk(f880_clk), .rst(f880_rst), .rdata(f880_rdata));
  assign f880_clk = clk;
  assign f880_rst = rst;
  // Bindings to f880

  // f882
  logic [0:0] f882_wen;
  logic [31:0] f882_wdata;
  logic [0:0] f882_clk;
  logic [0:0] f882_rst;
  logic [31:0] f882_rdata;
  sr_buffer_32_1 f882(.wen(f882_wen), .wdata(f882_wdata), .clk(f882_clk), .rst(f882_rst), .rdata(f882_rdata));
  assign f882_clk = clk;
  assign f882_rst = rst;
  // Bindings to f882

  // f884
  logic [0:0] f884_wen;
  logic [31:0] f884_wdata;
  logic [0:0] f884_clk;
  logic [0:0] f884_rst;
  logic [31:0] f884_rdata;
  sr_buffer_32_1 f884(.wen(f884_wen), .wdata(f884_wdata), .clk(f884_clk), .rst(f884_rst), .rdata(f884_rdata));
  assign f884_clk = clk;
  assign f884_rst = rst;
  // Bindings to f884

  // f886
  logic [0:0] f886_wen;
  logic [31:0] f886_wdata;
  logic [0:0] f886_clk;
  logic [0:0] f886_rst;
  logic [31:0] f886_rdata;
  sr_buffer_32_1 f886(.wen(f886_wen), .wdata(f886_wdata), .clk(f886_clk), .rst(f886_rst), .rdata(f886_rdata));
  assign f886_clk = clk;
  assign f886_rst = rst;
  // Bindings to f886

  // f888
  logic [0:0] f888_wen;
  logic [31:0] f888_wdata;
  logic [0:0] f888_clk;
  logic [0:0] f888_rst;
  logic [31:0] f888_rdata;
  sr_buffer_32_1 f888(.wen(f888_wen), .wdata(f888_wdata), .clk(f888_clk), .rst(f888_rst), .rdata(f888_rdata));
  assign f888_clk = clk;
  assign f888_rst = rst;
  // Bindings to f888

  // f890
  logic [0:0] f890_wen;
  logic [31:0] f890_wdata;
  logic [0:0] f890_clk;
  logic [0:0] f890_rst;
  logic [31:0] f890_rdata;
  sr_buffer_32_1 f890(.wen(f890_wen), .wdata(f890_wdata), .clk(f890_clk), .rst(f890_rst), .rdata(f890_rdata));
  assign f890_clk = clk;
  assign f890_rst = rst;
  // Bindings to f890

  // f892
  logic [0:0] f892_wen;
  logic [31:0] f892_wdata;
  logic [0:0] f892_clk;
  logic [0:0] f892_rst;
  logic [31:0] f892_rdata;
  sr_buffer_32_1 f892(.wen(f892_wen), .wdata(f892_wdata), .clk(f892_clk), .rst(f892_rst), .rdata(f892_rdata));
  assign f892_clk = clk;
  assign f892_rst = rst;
  // Bindings to f892

  // f894
  logic [0:0] f894_wen;
  logic [31:0] f894_wdata;
  logic [0:0] f894_clk;
  logic [0:0] f894_rst;
  logic [31:0] f894_rdata;
  sr_buffer_32_1 f894(.wen(f894_wen), .wdata(f894_wdata), .clk(f894_clk), .rst(f894_rst), .rdata(f894_rdata));
  assign f894_clk = clk;
  assign f894_rst = rst;
  // Bindings to f894

  // f896
  logic [0:0] f896_wen;
  logic [31:0] f896_wdata;
  logic [0:0] f896_clk;
  logic [0:0] f896_rst;
  logic [31:0] f896_rdata;
  sr_buffer_32_1 f896(.wen(f896_wen), .wdata(f896_wdata), .clk(f896_clk), .rst(f896_rst), .rdata(f896_rdata));
  assign f896_clk = clk;
  assign f896_rst = rst;
  // Bindings to f896

  // f898
  logic [0:0] f898_wen;
  logic [31:0] f898_wdata;
  logic [0:0] f898_clk;
  logic [0:0] f898_rst;
  logic [31:0] f898_rdata;
  sr_buffer_32_1 f898(.wen(f898_wen), .wdata(f898_wdata), .clk(f898_clk), .rst(f898_rst), .rdata(f898_rdata));
  assign f898_clk = clk;
  assign f898_rst = rst;
  // Bindings to f898

  // f900
  logic [0:0] f900_wen;
  logic [31:0] f900_wdata;
  logic [0:0] f900_clk;
  logic [0:0] f900_rst;
  logic [31:0] f900_rdata;
  sr_buffer_32_1 f900(.wen(f900_wen), .wdata(f900_wdata), .clk(f900_clk), .rst(f900_rst), .rdata(f900_rdata));
  assign f900_clk = clk;
  assign f900_rst = rst;
  // Bindings to f900

  // f902
  logic [0:0] f902_wen;
  logic [31:0] f902_wdata;
  logic [0:0] f902_clk;
  logic [0:0] f902_rst;
  logic [31:0] f902_rdata;
  sr_buffer_32_1 f902(.wen(f902_wen), .wdata(f902_wdata), .clk(f902_clk), .rst(f902_rst), .rdata(f902_rdata));
  assign f902_clk = clk;
  assign f902_rst = rst;
  // Bindings to f902

  // f904
  logic [0:0] f904_wen;
  logic [31:0] f904_wdata;
  logic [0:0] f904_clk;
  logic [0:0] f904_rst;
  logic [31:0] f904_rdata;
  sr_buffer_32_1 f904(.wen(f904_wen), .wdata(f904_wdata), .clk(f904_clk), .rst(f904_rst), .rdata(f904_rdata));
  assign f904_clk = clk;
  assign f904_rst = rst;
  // Bindings to f904

  // f906
  logic [0:0] f906_wen;
  logic [31:0] f906_wdata;
  logic [0:0] f906_clk;
  logic [0:0] f906_rst;
  logic [31:0] f906_rdata;
  sr_buffer_32_1 f906(.wen(f906_wen), .wdata(f906_wdata), .clk(f906_clk), .rst(f906_rst), .rdata(f906_rdata));
  assign f906_clk = clk;
  assign f906_rst = rst;
  // Bindings to f906

  // f908
  logic [0:0] f908_wen;
  logic [31:0] f908_wdata;
  logic [0:0] f908_clk;
  logic [0:0] f908_rst;
  logic [31:0] f908_rdata;
  sr_buffer_32_1 f908(.wen(f908_wen), .wdata(f908_wdata), .clk(f908_clk), .rst(f908_rst), .rdata(f908_rdata));
  assign f908_clk = clk;
  assign f908_rst = rst;
  // Bindings to f908

  // f910
  logic [0:0] f910_wen;
  logic [31:0] f910_wdata;
  logic [0:0] f910_clk;
  logic [0:0] f910_rst;
  logic [31:0] f910_rdata;
  sr_buffer_32_1 f910(.wen(f910_wen), .wdata(f910_wdata), .clk(f910_clk), .rst(f910_rst), .rdata(f910_rdata));
  assign f910_clk = clk;
  assign f910_rst = rst;
  // Bindings to f910

  // f912
  logic [0:0] f912_wen;
  logic [31:0] f912_wdata;
  logic [0:0] f912_clk;
  logic [0:0] f912_rst;
  logic [31:0] f912_rdata;
  sr_buffer_32_1 f912(.wen(f912_wen), .wdata(f912_wdata), .clk(f912_clk), .rst(f912_rst), .rdata(f912_rdata));
  assign f912_clk = clk;
  assign f912_rst = rst;
  // Bindings to f912

  // f914
  logic [0:0] f914_wen;
  logic [31:0] f914_wdata;
  logic [0:0] f914_clk;
  logic [0:0] f914_rst;
  logic [31:0] f914_rdata;
  sr_buffer_32_1 f914(.wen(f914_wen), .wdata(f914_wdata), .clk(f914_clk), .rst(f914_rst), .rdata(f914_rdata));
  assign f914_clk = clk;
  assign f914_rst = rst;
  // Bindings to f914

  // f916
  logic [0:0] f916_wen;
  logic [31:0] f916_wdata;
  logic [0:0] f916_clk;
  logic [0:0] f916_rst;
  logic [31:0] f916_rdata;
  sr_buffer_32_1 f916(.wen(f916_wen), .wdata(f916_wdata), .clk(f916_clk), .rst(f916_rst), .rdata(f916_rdata));
  assign f916_clk = clk;
  assign f916_rst = rst;
  // Bindings to f916

  // f918
  logic [0:0] f918_wen;
  logic [31:0] f918_wdata;
  logic [0:0] f918_clk;
  logic [0:0] f918_rst;
  logic [31:0] f918_rdata;
  sr_buffer_32_1 f918(.wen(f918_wen), .wdata(f918_wdata), .clk(f918_clk), .rst(f918_rst), .rdata(f918_rdata));
  assign f918_clk = clk;
  assign f918_rst = rst;
  // Bindings to f918

  // f920
  logic [0:0] f920_wen;
  logic [31:0] f920_wdata;
  logic [0:0] f920_clk;
  logic [0:0] f920_rst;
  logic [31:0] f920_rdata;
  sr_buffer_32_1 f920(.wen(f920_wen), .wdata(f920_wdata), .clk(f920_clk), .rst(f920_rst), .rdata(f920_rdata));
  assign f920_clk = clk;
  assign f920_rst = rst;
  // Bindings to f920

  // f922
  logic [0:0] f922_wen;
  logic [31:0] f922_wdata;
  logic [0:0] f922_clk;
  logic [0:0] f922_rst;
  logic [31:0] f922_rdata;
  sr_buffer_32_1 f922(.wen(f922_wen), .wdata(f922_wdata), .clk(f922_clk), .rst(f922_rst), .rdata(f922_rdata));
  assign f922_clk = clk;
  assign f922_rst = rst;
  // Bindings to f922

  // f924
  logic [0:0] f924_wen;
  logic [31:0] f924_wdata;
  logic [0:0] f924_clk;
  logic [0:0] f924_rst;
  logic [31:0] f924_rdata;
  sr_buffer_32_1 f924(.wen(f924_wen), .wdata(f924_wdata), .clk(f924_clk), .rst(f924_rst), .rdata(f924_rdata));
  assign f924_clk = clk;
  assign f924_rst = rst;
  // Bindings to f924

  // f926
  logic [0:0] f926_wen;
  logic [31:0] f926_wdata;
  logic [0:0] f926_clk;
  logic [0:0] f926_rst;
  logic [31:0] f926_rdata;
  sr_buffer_32_1 f926(.wen(f926_wen), .wdata(f926_wdata), .clk(f926_clk), .rst(f926_rst), .rdata(f926_rdata));
  assign f926_clk = clk;
  assign f926_rst = rst;
  // Bindings to f926

  // f928
  logic [0:0] f928_wen;
  logic [31:0] f928_wdata;
  logic [0:0] f928_clk;
  logic [0:0] f928_rst;
  logic [31:0] f928_rdata;
  sr_buffer_32_1 f928(.wen(f928_wen), .wdata(f928_wdata), .clk(f928_clk), .rst(f928_rst), .rdata(f928_rdata));
  assign f928_clk = clk;
  assign f928_rst = rst;
  // Bindings to f928

  // f930
  logic [0:0] f930_wen;
  logic [31:0] f930_wdata;
  logic [0:0] f930_clk;
  logic [0:0] f930_rst;
  logic [31:0] f930_rdata;
  sr_buffer_32_1 f930(.wen(f930_wen), .wdata(f930_wdata), .clk(f930_clk), .rst(f930_rst), .rdata(f930_rdata));
  assign f930_clk = clk;
  assign f930_rst = rst;
  // Bindings to f930

  // f932
  logic [0:0] f932_wen;
  logic [31:0] f932_wdata;
  logic [0:0] f932_clk;
  logic [0:0] f932_rst;
  logic [31:0] f932_rdata;
  sr_buffer_32_1 f932(.wen(f932_wen), .wdata(f932_wdata), .clk(f932_clk), .rst(f932_rst), .rdata(f932_rdata));
  assign f932_clk = clk;
  assign f932_rst = rst;
  // Bindings to f932

  // f934
  logic [0:0] f934_wen;
  logic [31:0] f934_wdata;
  logic [0:0] f934_clk;
  logic [0:0] f934_rst;
  logic [31:0] f934_rdata;
  sr_buffer_32_1 f934(.wen(f934_wen), .wdata(f934_wdata), .clk(f934_clk), .rst(f934_rst), .rdata(f934_rdata));
  assign f934_clk = clk;
  assign f934_rst = rst;
  // Bindings to f934

  // f936
  logic [0:0] f936_wen;
  logic [31:0] f936_wdata;
  logic [0:0] f936_clk;
  logic [0:0] f936_rst;
  logic [31:0] f936_rdata;
  sr_buffer_32_1 f936(.wen(f936_wen), .wdata(f936_wdata), .clk(f936_clk), .rst(f936_rst), .rdata(f936_rdata));
  assign f936_clk = clk;
  assign f936_rst = rst;
  // Bindings to f936

  // f938
  logic [0:0] f938_wen;
  logic [31:0] f938_wdata;
  logic [0:0] f938_clk;
  logic [0:0] f938_rst;
  logic [31:0] f938_rdata;
  sr_buffer_32_1 f938(.wen(f938_wen), .wdata(f938_wdata), .clk(f938_clk), .rst(f938_rst), .rdata(f938_rdata));
  assign f938_clk = clk;
  assign f938_rst = rst;
  // Bindings to f938

  // f940
  logic [0:0] f940_wen;
  logic [31:0] f940_wdata;
  logic [0:0] f940_clk;
  logic [0:0] f940_rst;
  logic [31:0] f940_rdata;
  sr_buffer_32_1 f940(.wen(f940_wen), .wdata(f940_wdata), .clk(f940_clk), .rst(f940_rst), .rdata(f940_rdata));
  assign f940_clk = clk;
  assign f940_rst = rst;
  // Bindings to f940

  // f942
  logic [0:0] f942_wen;
  logic [31:0] f942_wdata;
  logic [0:0] f942_clk;
  logic [0:0] f942_rst;
  logic [31:0] f942_rdata;
  sr_buffer_32_1 f942(.wen(f942_wen), .wdata(f942_wdata), .clk(f942_clk), .rst(f942_rst), .rdata(f942_rdata));
  assign f942_clk = clk;
  assign f942_rst = rst;
  // Bindings to f942

  // f944
  logic [0:0] f944_wen;
  logic [31:0] f944_wdata;
  logic [0:0] f944_clk;
  logic [0:0] f944_rst;
  logic [31:0] f944_rdata;
  sr_buffer_32_1 f944(.wen(f944_wen), .wdata(f944_wdata), .clk(f944_clk), .rst(f944_rst), .rdata(f944_rdata));
  assign f944_clk = clk;
  assign f944_rst = rst;
  // Bindings to f944

  // f946
  logic [0:0] f946_wen;
  logic [31:0] f946_wdata;
  logic [0:0] f946_clk;
  logic [0:0] f946_rst;
  logic [31:0] f946_rdata;
  sr_buffer_32_1 f946(.wen(f946_wen), .wdata(f946_wdata), .clk(f946_clk), .rst(f946_rst), .rdata(f946_rdata));
  assign f946_clk = clk;
  assign f946_rst = rst;
  // Bindings to f946

  // f948
  logic [0:0] f948_wen;
  logic [31:0] f948_wdata;
  logic [0:0] f948_clk;
  logic [0:0] f948_rst;
  logic [31:0] f948_rdata;
  sr_buffer_32_1 f948(.wen(f948_wen), .wdata(f948_wdata), .clk(f948_clk), .rst(f948_rst), .rdata(f948_rdata));
  assign f948_clk = clk;
  assign f948_rst = rst;
  // Bindings to f948

  // f950
  logic [0:0] f950_wen;
  logic [31:0] f950_wdata;
  logic [0:0] f950_clk;
  logic [0:0] f950_rst;
  logic [31:0] f950_rdata;
  sr_buffer_32_1 f950(.wen(f950_wen), .wdata(f950_wdata), .clk(f950_clk), .rst(f950_rst), .rdata(f950_rdata));
  assign f950_clk = clk;
  assign f950_rst = rst;
  // Bindings to f950

  // f952
  logic [0:0] f952_wen;
  logic [31:0] f952_wdata;
  logic [0:0] f952_clk;
  logic [0:0] f952_rst;
  logic [31:0] f952_rdata;
  sr_buffer_32_1 f952(.wen(f952_wen), .wdata(f952_wdata), .clk(f952_clk), .rst(f952_rst), .rdata(f952_rdata));
  assign f952_clk = clk;
  assign f952_rst = rst;
  // Bindings to f952

  // f954
  logic [0:0] f954_wen;
  logic [31:0] f954_wdata;
  logic [0:0] f954_clk;
  logic [0:0] f954_rst;
  logic [31:0] f954_rdata;
  sr_buffer_32_1 f954(.wen(f954_wen), .wdata(f954_wdata), .clk(f954_clk), .rst(f954_rst), .rdata(f954_rdata));
  assign f954_clk = clk;
  assign f954_rst = rst;
  // Bindings to f954

  // f956
  logic [0:0] f956_wen;
  logic [31:0] f956_wdata;
  logic [0:0] f956_clk;
  logic [0:0] f956_rst;
  logic [31:0] f956_rdata;
  sr_buffer_32_1 f956(.wen(f956_wen), .wdata(f956_wdata), .clk(f956_clk), .rst(f956_rst), .rdata(f956_rdata));
  assign f956_clk = clk;
  assign f956_rst = rst;
  // Bindings to f956

  // f958
  logic [0:0] f958_wen;
  logic [31:0] f958_wdata;
  logic [0:0] f958_clk;
  logic [0:0] f958_rst;
  logic [31:0] f958_rdata;
  sr_buffer_32_1 f958(.wen(f958_wen), .wdata(f958_wdata), .clk(f958_clk), .rst(f958_rst), .rdata(f958_rdata));
  assign f958_clk = clk;
  assign f958_rst = rst;
  // Bindings to f958

  // f960
  logic [0:0] f960_wen;
  logic [31:0] f960_wdata;
  logic [0:0] f960_clk;
  logic [0:0] f960_rst;
  logic [31:0] f960_rdata;
  sr_buffer_32_1 f960(.wen(f960_wen), .wdata(f960_wdata), .clk(f960_clk), .rst(f960_rst), .rdata(f960_rdata));
  assign f960_clk = clk;
  assign f960_rst = rst;
  // Bindings to f960

  // f980
  logic [0:0] f980_wen;
  logic [31:0] f980_wdata;
  logic [0:0] f980_clk;
  logic [0:0] f980_rst;
  logic [31:0] f980_rdata;
  sr_buffer_32_1 f980(.wen(f980_wen), .wdata(f980_wdata), .clk(f980_clk), .rst(f980_rst), .rdata(f980_rdata));
  assign f980_clk = clk;
  assign f980_rst = rst;
  // Bindings to f980



endmodule


module dark_gauss_blur_1_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module dark_gauss_blur_1_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1265;
    end
  end

endmodule


module in_wire_dark_update_0_write_wen(output [0:0] dark_update_0_write_wen);

endmodule


module dark_gauss_blur_1_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2527;
    end
  end

endmodule


module dark_gauss_blur_1_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1264;
    end
  end

endmodule


module dark_gauss_blur_1_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module dark_gauss_blur_1_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_weights_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_gauss_blur_1_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (1259 - d0 >= 0) ? (2526) : (-1260 + d0 == 0) ? (2526) : 0;
    end
  end

endmodule


module dark_gauss_blur_1_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (1259 - d0 >= 0) ? (1263) : (-1260 + d0 == 0) ? (1263) : 0;
    end
  end

endmodule


module in_wire_dark_update_0_write_wdata(output [31:0] dark_update_0_write_wdata);

endmodule


module dark(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_update_0_write_wen, input [31:0] dark_weights_update_0_read_dummy, input [31:0] dark_update_0_write_wdata, input [287:0] dark_gauss_blur_1_update_0_read_dummy, output [287:0] dark_gauss_blur_1_update_0_read_rdata, input [31:0] dark_laplace_diff_0_update_0_read_dummy, output [31:0] dark_laplace_diff_0_update_0_read_rdata, output [31:0] dark_weights_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;
  logic [31:0] rd_6;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;
  reg [31:0] rd_6_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;
      rd_6_stage_1 <= rd_6;


    end

  end


  // Data processing units...
  // dark_dark_update_0_write0_merged_banks_10
  logic [0:0] dark_dark_update_0_write0_merged_banks_10_clk;
  logic [0:0] dark_dark_update_0_write0_merged_banks_10_rst;
  logic [0:0] dark_dark_update_0_write0_merged_banks_10_start;
  logic [0:0] dark_dark_update_0_write0_merged_banks_10_done;
  dark_dark_update_0_write0_merged_banks_10 dark_dark_update_0_write0_merged_banks_10(.clk(dark_dark_update_0_write0_merged_banks_10_clk), .rst(dark_dark_update_0_write0_merged_banks_10_rst), .start(dark_dark_update_0_write0_merged_banks_10_start), .done(dark_dark_update_0_write0_merged_banks_10_done));
  assign dark_dark_update_0_write0_merged_banks_10_clk = clk;
  assign dark_dark_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to dark_dark_update_0_write0_merged_banks_10

  // Bindings to dark_update_0_write_wen
    // rd_0
  assign rd_0 = dark_update_0_write_wen;

  // Bindings to dark_weights_update_0_read_dummy
    // rd_6
  assign rd_6 = dark_weights_update_0_read_dummy;

  // dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0
  logic [0:0] dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_clk;
  logic [0:0] dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_rst;
  logic [0:0] dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_start;
  logic [0:0] dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_done;
  dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0 dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0(.clk(dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_clk), .rst(dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_rst), .start(dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_start), .done(dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_done));
  assign dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_clk = clk;
  assign dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0_rst = rst;
  // Bindings to dark_dark_update_0_write0_to_dark_laplace_diff_0_rd0

  // selector_dark_gauss_blur_1_rd0_select
  logic [0:0] selector_dark_gauss_blur_1_rd0_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd0_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd0_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd0_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd0_select_out;
  dark_gauss_blur_1_rd0_select selector_dark_gauss_blur_1_rd0_select(.clk(selector_dark_gauss_blur_1_rd0_select_clk), .rst(selector_dark_gauss_blur_1_rd0_select_rst), .d0(selector_dark_gauss_blur_1_rd0_select_d0), .d1(selector_dark_gauss_blur_1_rd0_select_d1), .out(selector_dark_gauss_blur_1_rd0_select_out));
  assign selector_dark_gauss_blur_1_rd0_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd0_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd0_select

  // selector_dark_gauss_blur_1_rd1_select
  logic [0:0] selector_dark_gauss_blur_1_rd1_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd1_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd1_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd1_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd1_select_out;
  dark_gauss_blur_1_rd1_select selector_dark_gauss_blur_1_rd1_select(.clk(selector_dark_gauss_blur_1_rd1_select_clk), .rst(selector_dark_gauss_blur_1_rd1_select_rst), .d0(selector_dark_gauss_blur_1_rd1_select_d0), .d1(selector_dark_gauss_blur_1_rd1_select_d1), .out(selector_dark_gauss_blur_1_rd1_select_out));
  assign selector_dark_gauss_blur_1_rd1_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd1_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd1_select

  // selector_dark_gauss_blur_1_rd2_select
  logic [0:0] selector_dark_gauss_blur_1_rd2_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd2_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd2_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd2_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd2_select_out;
  dark_gauss_blur_1_rd2_select selector_dark_gauss_blur_1_rd2_select(.clk(selector_dark_gauss_blur_1_rd2_select_clk), .rst(selector_dark_gauss_blur_1_rd2_select_rst), .d0(selector_dark_gauss_blur_1_rd2_select_d0), .d1(selector_dark_gauss_blur_1_rd2_select_d1), .out(selector_dark_gauss_blur_1_rd2_select_out));
  assign selector_dark_gauss_blur_1_rd2_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd2_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd2_select

  // selector_dark_gauss_blur_1_rd3_select
  logic [0:0] selector_dark_gauss_blur_1_rd3_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd3_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd3_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd3_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd3_select_out;
  dark_gauss_blur_1_rd3_select selector_dark_gauss_blur_1_rd3_select(.clk(selector_dark_gauss_blur_1_rd3_select_clk), .rst(selector_dark_gauss_blur_1_rd3_select_rst), .d0(selector_dark_gauss_blur_1_rd3_select_d0), .d1(selector_dark_gauss_blur_1_rd3_select_d1), .out(selector_dark_gauss_blur_1_rd3_select_out));
  assign selector_dark_gauss_blur_1_rd3_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd3_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd3_select

  // selector_dark_gauss_blur_1_rd4_select
  logic [0:0] selector_dark_gauss_blur_1_rd4_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd4_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd4_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd4_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd4_select_out;
  dark_gauss_blur_1_rd4_select selector_dark_gauss_blur_1_rd4_select(.clk(selector_dark_gauss_blur_1_rd4_select_clk), .rst(selector_dark_gauss_blur_1_rd4_select_rst), .d0(selector_dark_gauss_blur_1_rd4_select_d0), .d1(selector_dark_gauss_blur_1_rd4_select_d1), .out(selector_dark_gauss_blur_1_rd4_select_out));
  assign selector_dark_gauss_blur_1_rd4_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd4_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd4_select

  // selector_dark_gauss_blur_1_rd5_select
  logic [0:0] selector_dark_gauss_blur_1_rd5_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd5_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd5_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd5_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd5_select_out;
  dark_gauss_blur_1_rd5_select selector_dark_gauss_blur_1_rd5_select(.clk(selector_dark_gauss_blur_1_rd5_select_clk), .rst(selector_dark_gauss_blur_1_rd5_select_rst), .d0(selector_dark_gauss_blur_1_rd5_select_d0), .d1(selector_dark_gauss_blur_1_rd5_select_d1), .out(selector_dark_gauss_blur_1_rd5_select_out));
  assign selector_dark_gauss_blur_1_rd5_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd5_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd5_select

  // selector_dark_gauss_blur_1_rd6_select
  logic [0:0] selector_dark_gauss_blur_1_rd6_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd6_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd6_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd6_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd6_select_out;
  dark_gauss_blur_1_rd6_select selector_dark_gauss_blur_1_rd6_select(.clk(selector_dark_gauss_blur_1_rd6_select_clk), .rst(selector_dark_gauss_blur_1_rd6_select_rst), .d0(selector_dark_gauss_blur_1_rd6_select_d0), .d1(selector_dark_gauss_blur_1_rd6_select_d1), .out(selector_dark_gauss_blur_1_rd6_select_out));
  assign selector_dark_gauss_blur_1_rd6_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd6_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd6_select

  // selector_dark_gauss_blur_1_rd7_select
  logic [0:0] selector_dark_gauss_blur_1_rd7_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd7_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd7_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd7_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd7_select_out;
  dark_gauss_blur_1_rd7_select selector_dark_gauss_blur_1_rd7_select(.clk(selector_dark_gauss_blur_1_rd7_select_clk), .rst(selector_dark_gauss_blur_1_rd7_select_rst), .d0(selector_dark_gauss_blur_1_rd7_select_d0), .d1(selector_dark_gauss_blur_1_rd7_select_d1), .out(selector_dark_gauss_blur_1_rd7_select_out));
  assign selector_dark_gauss_blur_1_rd7_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd7_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd7_select

  // selector_dark_gauss_blur_1_rd8_select
  logic [0:0] selector_dark_gauss_blur_1_rd8_select_clk;
  logic [0:0] selector_dark_gauss_blur_1_rd8_select_rst;
  logic [31:0] selector_dark_gauss_blur_1_rd8_select_d0;
  logic [31:0] selector_dark_gauss_blur_1_rd8_select_d1;
  logic [31:0] selector_dark_gauss_blur_1_rd8_select_out;
  dark_gauss_blur_1_rd8_select selector_dark_gauss_blur_1_rd8_select(.clk(selector_dark_gauss_blur_1_rd8_select_clk), .rst(selector_dark_gauss_blur_1_rd8_select_rst), .d0(selector_dark_gauss_blur_1_rd8_select_d0), .d1(selector_dark_gauss_blur_1_rd8_select_d1), .out(selector_dark_gauss_blur_1_rd8_select_out));
  assign selector_dark_gauss_blur_1_rd8_select_clk = clk;
  assign selector_dark_gauss_blur_1_rd8_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_1_rd8_select

  // Bindings to dark_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_update_0_write_wdata;

  // selector_dark_laplace_diff_0_rd0_select
  logic [0:0] selector_dark_laplace_diff_0_rd0_select_clk;
  logic [0:0] selector_dark_laplace_diff_0_rd0_select_rst;
  logic [31:0] selector_dark_laplace_diff_0_rd0_select_d0;
  logic [31:0] selector_dark_laplace_diff_0_rd0_select_d1;
  logic [31:0] selector_dark_laplace_diff_0_rd0_select_out;
  dark_laplace_diff_0_rd0_select selector_dark_laplace_diff_0_rd0_select(.clk(selector_dark_laplace_diff_0_rd0_select_clk), .rst(selector_dark_laplace_diff_0_rd0_select_rst), .d0(selector_dark_laplace_diff_0_rd0_select_d0), .d1(selector_dark_laplace_diff_0_rd0_select_d1), .out(selector_dark_laplace_diff_0_rd0_select_out));
  assign selector_dark_laplace_diff_0_rd0_select_clk = clk;
  assign selector_dark_laplace_diff_0_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_diff_0_rd0_select

  // selector_dark_weights_rd0_select
  logic [0:0] selector_dark_weights_rd0_select_clk;
  logic [0:0] selector_dark_weights_rd0_select_rst;
  logic [31:0] selector_dark_weights_rd0_select_d0;
  logic [31:0] selector_dark_weights_rd0_select_d1;
  logic [31:0] selector_dark_weights_rd0_select_out;
  dark_weights_rd0_select selector_dark_weights_rd0_select(.clk(selector_dark_weights_rd0_select_clk), .rst(selector_dark_weights_rd0_select_rst), .d0(selector_dark_weights_rd0_select_d0), .d1(selector_dark_weights_rd0_select_d1), .out(selector_dark_weights_rd0_select_out));
  assign selector_dark_weights_rd0_select_clk = clk;
  assign selector_dark_weights_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_rd0_select

  // Bindings to dark_gauss_blur_1_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_gauss_blur_1_update_0_read_dummy;

  // Bindings to dark_gauss_blur_1_update_0_read_rdata
    // wr_3
  assign dark_gauss_blur_1_update_0_read_rdata = rd_2;

  // Bindings to dark_laplace_diff_0_update_0_read_dummy
    // rd_4
  assign rd_4 = dark_laplace_diff_0_update_0_read_dummy;

  // Bindings to dark_laplace_diff_0_update_0_read_rdata
    // wr_5
  assign dark_laplace_diff_0_update_0_read_rdata = rd_4;

  // Bindings to dark_weights_update_0_read_rdata
    // wr_7
  assign dark_weights_update_0_read_rdata = rd_6;



endmodule


module in_wire_dark_gauss_blur_1_update_0_read_dummy(output [287:0] dark_gauss_blur_1_update_0_read_dummy);

endmodule


module out_wire_dark_gauss_blur_1_update_0_read_rdata(input [287:0] dark_gauss_blur_1_update_0_read_rdata);

endmodule


module in_wire_dark_laplace_diff_0_update_0_read_dummy(output [31:0] dark_laplace_diff_0_update_0_read_dummy);

endmodule


module out_wire_dark_laplace_diff_0_update_0_read_rdata(input [31:0] dark_laplace_diff_0_update_0_read_rdata);

endmodule


module in_wire_dark_weights_update_0_read_dummy(output [31:0] dark_weights_update_0_read_dummy);

endmodule


module out_wire_dark_weights_update_0_read_rdata(input [31:0] dark_weights_update_0_read_rdata);

endmodule


module dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_gauss_blur_1_update_0_write_wen(output [0:0] dark_gauss_blur_1_update_0_write_wen);

endmodule


module dark_gauss_ds_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_gauss_blur_1_update_0_write_wdata(output [31:0] dark_gauss_blur_1_update_0_write_wdata);

endmodule


module in_wire_dark_gauss_ds_1_update_0_read_dummy(output [31:0] dark_gauss_ds_1_update_0_read_dummy);

endmodule


module out_wire_dark_gauss_ds_1_update_0_read_rdata(input [31:0] dark_gauss_ds_1_update_0_read_rdata);

endmodule


module dark_gauss_blur_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_gauss_blur_1_update_0_write_wen, input [31:0] dark_gauss_ds_1_update_0_read_dummy, input [31:0] dark_gauss_blur_1_update_0_write_wdata, output [31:0] dark_gauss_ds_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_gauss_blur_1_update_0_write_wen
    // rd_0
  assign rd_0 = dark_gauss_blur_1_update_0_write_wen;

  // dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1
  logic [0:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_done;
  dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1 dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1(.clk(dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_clk), .rst(dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_rst), .start(dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_start), .done(dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_done));
  assign dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_clk = clk;
  assign dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_gauss_blur_1_dark_gauss_blur_1_update_0_write0_merged_banks_1

  // Bindings to dark_gauss_ds_1_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_gauss_ds_1_update_0_read_dummy;

  // selector_dark_gauss_ds_1_rd0_select
  logic [0:0] selector_dark_gauss_ds_1_rd0_select_clk;
  logic [0:0] selector_dark_gauss_ds_1_rd0_select_rst;
  logic [31:0] selector_dark_gauss_ds_1_rd0_select_d0;
  logic [31:0] selector_dark_gauss_ds_1_rd0_select_d1;
  logic [31:0] selector_dark_gauss_ds_1_rd0_select_out;
  dark_gauss_ds_1_rd0_select selector_dark_gauss_ds_1_rd0_select(.clk(selector_dark_gauss_ds_1_rd0_select_clk), .rst(selector_dark_gauss_ds_1_rd0_select_rst), .d0(selector_dark_gauss_ds_1_rd0_select_d0), .d1(selector_dark_gauss_ds_1_rd0_select_d1), .out(selector_dark_gauss_ds_1_rd0_select_out));
  assign selector_dark_gauss_ds_1_rd0_select_clk = clk;
  assign selector_dark_gauss_ds_1_rd0_select_rst = rst;
  // Bindings to selector_dark_gauss_ds_1_rd0_select

  // Bindings to dark_gauss_blur_1_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_gauss_blur_1_update_0_write_wdata;

  // Bindings to dark_gauss_ds_1_update_0_read_rdata
    // wr_3
  assign dark_gauss_ds_1_update_0_read_rdata = rd_2;



endmodule


module dark_gauss_ds_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] dark_laplace_us_0_update_0_read_rdata, output [31:0] dark_laplace_diff_1_update_0_read_rdata, input [287:0] dark_gauss_blur_2_update_0_read_dummy, input [31:0] dark_laplace_us_0_update_0_read_dummy, input [31:0] dark_laplace_diff_1_update_0_read_dummy, output [287:0] dark_gauss_blur_2_update_0_read_rdata, input [0:0] dark_gauss_ds_1_update_0_write_wen, input [31:0] dark_gauss_ds_1_update_0_write_wdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;
  logic [31:0] rd_6;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;
  reg [31:0] rd_6_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;
      rd_6_stage_1 <= rd_6;


    end

  end


  // Data processing units...
  // Bindings to dark_laplace_us_0_update_0_read_rdata
    // wr_7
  assign dark_laplace_us_0_update_0_read_rdata = rd_6;

  // Bindings to dark_laplace_diff_1_update_0_read_rdata
    // wr_5
  assign dark_laplace_diff_1_update_0_read_rdata = rd_4;

  // dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_clk;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_rst;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_start;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_done;
  dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0 dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0(.clk(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_clk), .rst(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_rst), .start(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_start), .done(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_done));
  assign dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_clk = clk;
  assign dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0_rst = rst;
  // Bindings to dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_to_dark_laplace_us_0_rd0

  // Bindings to dark_gauss_blur_2_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_gauss_blur_2_update_0_read_dummy;

  // Bindings to dark_laplace_us_0_update_0_read_dummy
    // rd_6
  assign rd_6 = dark_laplace_us_0_update_0_read_dummy;

  // Bindings to dark_laplace_diff_1_update_0_read_dummy
    // rd_4
  assign rd_4 = dark_laplace_diff_1_update_0_read_dummy;

  // Bindings to dark_gauss_blur_2_update_0_read_rdata
    // wr_3
  assign dark_gauss_blur_2_update_0_read_rdata = rd_2;

  // dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10_clk;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10_rst;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10_start;
  logic [0:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10_done;
  dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10 dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10(.clk(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10_clk), .rst(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10_rst), .start(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10_start), .done(dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10_done));
  assign dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10_clk = clk;
  assign dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10

  // Bindings to dark_gauss_ds_1_update_0_write_wen
    // rd_0
  assign rd_0 = dark_gauss_ds_1_update_0_write_wen;

  // Bindings to dark_gauss_ds_1_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_gauss_ds_1_update_0_write_wdata;

  // selector_dark_laplace_diff_1_rd0_select
  logic [0:0] selector_dark_laplace_diff_1_rd0_select_clk;
  logic [0:0] selector_dark_laplace_diff_1_rd0_select_rst;
  logic [31:0] selector_dark_laplace_diff_1_rd0_select_d0;
  logic [31:0] selector_dark_laplace_diff_1_rd0_select_d1;
  logic [31:0] selector_dark_laplace_diff_1_rd0_select_out;
  dark_laplace_diff_1_rd0_select selector_dark_laplace_diff_1_rd0_select(.clk(selector_dark_laplace_diff_1_rd0_select_clk), .rst(selector_dark_laplace_diff_1_rd0_select_rst), .d0(selector_dark_laplace_diff_1_rd0_select_d0), .d1(selector_dark_laplace_diff_1_rd0_select_d1), .out(selector_dark_laplace_diff_1_rd0_select_out));
  assign selector_dark_laplace_diff_1_rd0_select_clk = clk;
  assign selector_dark_laplace_diff_1_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_diff_1_rd0_select

  // selector_dark_laplace_us_0_rd0_select
  logic [0:0] selector_dark_laplace_us_0_rd0_select_clk;
  logic [0:0] selector_dark_laplace_us_0_rd0_select_rst;
  logic [31:0] selector_dark_laplace_us_0_rd0_select_d0;
  logic [31:0] selector_dark_laplace_us_0_rd0_select_d1;
  logic [31:0] selector_dark_laplace_us_0_rd0_select_out;
  dark_laplace_us_0_rd0_select selector_dark_laplace_us_0_rd0_select(.clk(selector_dark_laplace_us_0_rd0_select_clk), .rst(selector_dark_laplace_us_0_rd0_select_rst), .d0(selector_dark_laplace_us_0_rd0_select_d0), .d1(selector_dark_laplace_us_0_rd0_select_d1), .out(selector_dark_laplace_us_0_rd0_select_out));
  assign selector_dark_laplace_us_0_rd0_select_clk = clk;
  assign selector_dark_laplace_us_0_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_us_0_rd0_select

  // selector_dark_gauss_blur_2_rd8_select
  logic [0:0] selector_dark_gauss_blur_2_rd8_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd8_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd8_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd8_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd8_select_out;
  dark_gauss_blur_2_rd8_select selector_dark_gauss_blur_2_rd8_select(.clk(selector_dark_gauss_blur_2_rd8_select_clk), .rst(selector_dark_gauss_blur_2_rd8_select_rst), .d0(selector_dark_gauss_blur_2_rd8_select_d0), .d1(selector_dark_gauss_blur_2_rd8_select_d1), .out(selector_dark_gauss_blur_2_rd8_select_out));
  assign selector_dark_gauss_blur_2_rd8_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd8_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd8_select

  // selector_dark_gauss_blur_2_rd7_select
  logic [0:0] selector_dark_gauss_blur_2_rd7_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd7_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd7_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd7_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd7_select_out;
  dark_gauss_blur_2_rd7_select selector_dark_gauss_blur_2_rd7_select(.clk(selector_dark_gauss_blur_2_rd7_select_clk), .rst(selector_dark_gauss_blur_2_rd7_select_rst), .d0(selector_dark_gauss_blur_2_rd7_select_d0), .d1(selector_dark_gauss_blur_2_rd7_select_d1), .out(selector_dark_gauss_blur_2_rd7_select_out));
  assign selector_dark_gauss_blur_2_rd7_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd7_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd7_select

  // selector_dark_gauss_blur_2_rd6_select
  logic [0:0] selector_dark_gauss_blur_2_rd6_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd6_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd6_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd6_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd6_select_out;
  dark_gauss_blur_2_rd6_select selector_dark_gauss_blur_2_rd6_select(.clk(selector_dark_gauss_blur_2_rd6_select_clk), .rst(selector_dark_gauss_blur_2_rd6_select_rst), .d0(selector_dark_gauss_blur_2_rd6_select_d0), .d1(selector_dark_gauss_blur_2_rd6_select_d1), .out(selector_dark_gauss_blur_2_rd6_select_out));
  assign selector_dark_gauss_blur_2_rd6_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd6_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd6_select

  // selector_dark_gauss_blur_2_rd5_select
  logic [0:0] selector_dark_gauss_blur_2_rd5_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd5_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd5_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd5_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd5_select_out;
  dark_gauss_blur_2_rd5_select selector_dark_gauss_blur_2_rd5_select(.clk(selector_dark_gauss_blur_2_rd5_select_clk), .rst(selector_dark_gauss_blur_2_rd5_select_rst), .d0(selector_dark_gauss_blur_2_rd5_select_d0), .d1(selector_dark_gauss_blur_2_rd5_select_d1), .out(selector_dark_gauss_blur_2_rd5_select_out));
  assign selector_dark_gauss_blur_2_rd5_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd5_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd5_select

  // selector_dark_gauss_blur_2_rd3_select
  logic [0:0] selector_dark_gauss_blur_2_rd3_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd3_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd3_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd3_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd3_select_out;
  dark_gauss_blur_2_rd3_select selector_dark_gauss_blur_2_rd3_select(.clk(selector_dark_gauss_blur_2_rd3_select_clk), .rst(selector_dark_gauss_blur_2_rd3_select_rst), .d0(selector_dark_gauss_blur_2_rd3_select_d0), .d1(selector_dark_gauss_blur_2_rd3_select_d1), .out(selector_dark_gauss_blur_2_rd3_select_out));
  assign selector_dark_gauss_blur_2_rd3_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd3_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd3_select

  // selector_dark_gauss_blur_2_rd4_select
  logic [0:0] selector_dark_gauss_blur_2_rd4_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd4_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd4_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd4_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd4_select_out;
  dark_gauss_blur_2_rd4_select selector_dark_gauss_blur_2_rd4_select(.clk(selector_dark_gauss_blur_2_rd4_select_clk), .rst(selector_dark_gauss_blur_2_rd4_select_rst), .d0(selector_dark_gauss_blur_2_rd4_select_d0), .d1(selector_dark_gauss_blur_2_rd4_select_d1), .out(selector_dark_gauss_blur_2_rd4_select_out));
  assign selector_dark_gauss_blur_2_rd4_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd4_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd4_select

  // selector_dark_gauss_blur_2_rd2_select
  logic [0:0] selector_dark_gauss_blur_2_rd2_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd2_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd2_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd2_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd2_select_out;
  dark_gauss_blur_2_rd2_select selector_dark_gauss_blur_2_rd2_select(.clk(selector_dark_gauss_blur_2_rd2_select_clk), .rst(selector_dark_gauss_blur_2_rd2_select_rst), .d0(selector_dark_gauss_blur_2_rd2_select_d0), .d1(selector_dark_gauss_blur_2_rd2_select_d1), .out(selector_dark_gauss_blur_2_rd2_select_out));
  assign selector_dark_gauss_blur_2_rd2_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd2_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd2_select

  // selector_dark_gauss_blur_2_rd0_select
  logic [0:0] selector_dark_gauss_blur_2_rd0_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd0_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd0_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd0_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd0_select_out;
  dark_gauss_blur_2_rd0_select selector_dark_gauss_blur_2_rd0_select(.clk(selector_dark_gauss_blur_2_rd0_select_clk), .rst(selector_dark_gauss_blur_2_rd0_select_rst), .d0(selector_dark_gauss_blur_2_rd0_select_d0), .d1(selector_dark_gauss_blur_2_rd0_select_d1), .out(selector_dark_gauss_blur_2_rd0_select_out));
  assign selector_dark_gauss_blur_2_rd0_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd0_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd0_select

  // selector_dark_gauss_blur_2_rd1_select
  logic [0:0] selector_dark_gauss_blur_2_rd1_select_clk;
  logic [0:0] selector_dark_gauss_blur_2_rd1_select_rst;
  logic [31:0] selector_dark_gauss_blur_2_rd1_select_d0;
  logic [31:0] selector_dark_gauss_blur_2_rd1_select_d1;
  logic [31:0] selector_dark_gauss_blur_2_rd1_select_out;
  dark_gauss_blur_2_rd1_select selector_dark_gauss_blur_2_rd1_select(.clk(selector_dark_gauss_blur_2_rd1_select_clk), .rst(selector_dark_gauss_blur_2_rd1_select_rst), .d0(selector_dark_gauss_blur_2_rd1_select_d0), .d1(selector_dark_gauss_blur_2_rd1_select_d1), .out(selector_dark_gauss_blur_2_rd1_select_out));
  assign selector_dark_gauss_blur_2_rd1_select_clk = clk;
  assign selector_dark_gauss_blur_2_rd1_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_2_rd1_select



endmodule


module dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236



endmodule


module in_wire_dark_gauss_ds_3_update_0_write_wen(output [0:0] dark_gauss_ds_3_update_0_write_wen);

endmodule


module dark_laplace_us_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = ((-1 - d1) % 2 == 0 && 311 - d0 >= 0) ? ((156 - floord(2*d0, 4))) : 0;
    end
  end

endmodule


module in_wire_dark_gauss_ds_3_update_0_write_wdata(output [31:0] dark_gauss_ds_3_update_0_write_wdata);

endmodule


module in_wire_dark_laplace_us_2_update_0_read_dummy(output [31:0] dark_laplace_us_2_update_0_read_dummy);

endmodule


module out_wire_dark_laplace_us_2_update_0_read_rdata(input [31:0] dark_laplace_us_2_update_0_read_rdata);

endmodule


module dark_gauss_ds_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_gauss_ds_3_update_0_write_wen, input [31:0] dark_gauss_ds_3_update_0_write_wdata, input [31:0] dark_laplace_us_2_update_0_read_dummy, output [31:0] dark_laplace_us_2_update_0_read_rdata, input [31:0] fused_level_3_update_0_read_dummy, output [31:0] fused_level_3_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // Bindings to dark_gauss_ds_3_update_0_write_wen
    // rd_0
  assign rd_0 = dark_gauss_ds_3_update_0_write_wen;

  // dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_clk;
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_rst;
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_start;
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_done;
  dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0 dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0(.clk(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_clk), .rst(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_rst), .start(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_start), .done(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_done));
  assign dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_clk = clk;
  assign dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0_rst = rst;
  // Bindings to dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_to_dark_laplace_us_2_rd0

  // selector_fused_level_3_rd0_select
  logic [0:0] selector_fused_level_3_rd0_select_clk;
  logic [0:0] selector_fused_level_3_rd0_select_rst;
  logic [31:0] selector_fused_level_3_rd0_select_d0;
  logic [31:0] selector_fused_level_3_rd0_select_d1;
  logic [31:0] selector_fused_level_3_rd0_select_out;
  fused_level_3_rd0_select selector_fused_level_3_rd0_select(.clk(selector_fused_level_3_rd0_select_clk), .rst(selector_fused_level_3_rd0_select_rst), .d0(selector_fused_level_3_rd0_select_d0), .d1(selector_fused_level_3_rd0_select_d1), .out(selector_fused_level_3_rd0_select_out));
  assign selector_fused_level_3_rd0_select_clk = clk;
  assign selector_fused_level_3_rd0_select_rst = rst;
  // Bindings to selector_fused_level_3_rd0_select

  // selector_dark_laplace_us_2_rd0_select
  logic [0:0] selector_dark_laplace_us_2_rd0_select_clk;
  logic [0:0] selector_dark_laplace_us_2_rd0_select_rst;
  logic [31:0] selector_dark_laplace_us_2_rd0_select_d0;
  logic [31:0] selector_dark_laplace_us_2_rd0_select_d1;
  logic [31:0] selector_dark_laplace_us_2_rd0_select_out;
  dark_laplace_us_2_rd0_select selector_dark_laplace_us_2_rd0_select(.clk(selector_dark_laplace_us_2_rd0_select_clk), .rst(selector_dark_laplace_us_2_rd0_select_rst), .d0(selector_dark_laplace_us_2_rd0_select_d0), .d1(selector_dark_laplace_us_2_rd0_select_d1), .out(selector_dark_laplace_us_2_rd0_select_out));
  assign selector_dark_laplace_us_2_rd0_select_clk = clk;
  assign selector_dark_laplace_us_2_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_us_2_rd0_select

  // dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_done;
  dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1 dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1(.clk(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_clk), .rst(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_rst), .start(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_start), .done(dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_done));
  assign dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_clk = clk;
  assign dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_gauss_ds_3_dark_gauss_ds_3_update_0_write0_merged_banks_1

  // Bindings to dark_gauss_ds_3_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_gauss_ds_3_update_0_write_wdata;

  // Bindings to dark_laplace_us_2_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_laplace_us_2_update_0_read_dummy;

  // Bindings to dark_laplace_us_2_update_0_read_rdata
    // wr_3
  assign dark_laplace_us_2_update_0_read_rdata = rd_2;

  // Bindings to fused_level_3_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_3_update_0_read_dummy;

  // Bindings to fused_level_3_update_0_read_rdata
    // wr_5
  assign fused_level_3_update_0_read_rdata = rd_4;



endmodule


module dark_weights_normed_gauss_blur_1_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (1259 - d0 >= 0) ? (2526) : (-1260 + d0 == 0) ? (2526) : 0;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2528;
    end
  end

endmodule


module dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1454
  logic [0:0] f1454_wen;
  logic [31:0] f1454_wdata;
  logic [0:0] f1454_clk;
  logic [0:0] f1454_rst;
  logic [31:0] f1454_rdata;
  sr_buffer_32_1 f1454(.wen(f1454_wen), .wdata(f1454_wdata), .clk(f1454_clk), .rst(f1454_rst), .rdata(f1454_rdata));
  assign f1454_clk = clk;
  assign f1454_rst = rst;
  // Bindings to f1454

  // f1456
  logic [0:0] f1456_wen;
  logic [31:0] f1456_wdata;
  logic [0:0] f1456_clk;
  logic [0:0] f1456_rst;
  logic [31:0] f1456_rdata;
  sr_buffer_32_1 f1456(.wen(f1456_wen), .wdata(f1456_wdata), .clk(f1456_clk), .rst(f1456_rst), .rdata(f1456_rdata));
  assign f1456_clk = clk;
  assign f1456_rst = rst;
  // Bindings to f1456

  // f1458
  logic [0:0] f1458_wen;
  logic [31:0] f1458_wdata;
  logic [0:0] f1458_clk;
  logic [0:0] f1458_rst;
  logic [31:0] f1458_rdata;
  sr_buffer_32_1 f1458(.wen(f1458_wen), .wdata(f1458_wdata), .clk(f1458_clk), .rst(f1458_rst), .rdata(f1458_rdata));
  assign f1458_clk = clk;
  assign f1458_rst = rst;
  // Bindings to f1458

  // f1460
  logic [0:0] f1460_wen;
  logic [31:0] f1460_wdata;
  logic [0:0] f1460_clk;
  logic [0:0] f1460_rst;
  logic [31:0] f1460_rdata;
  sr_buffer_32_1 f1460(.wen(f1460_wen), .wdata(f1460_wdata), .clk(f1460_clk), .rst(f1460_rst), .rdata(f1460_rdata));
  assign f1460_clk = clk;
  assign f1460_rst = rst;
  // Bindings to f1460

  // f1462
  logic [0:0] f1462_wen;
  logic [31:0] f1462_wdata;
  logic [0:0] f1462_clk;
  logic [0:0] f1462_rst;
  logic [31:0] f1462_rdata;
  sr_buffer_32_1 f1462(.wen(f1462_wen), .wdata(f1462_wdata), .clk(f1462_clk), .rst(f1462_rst), .rdata(f1462_rdata));
  assign f1462_clk = clk;
  assign f1462_rst = rst;
  // Bindings to f1462

  // f1464
  logic [0:0] f1464_wen;
  logic [31:0] f1464_wdata;
  logic [0:0] f1464_clk;
  logic [0:0] f1464_rst;
  logic [31:0] f1464_rdata;
  sr_buffer_32_1 f1464(.wen(f1464_wen), .wdata(f1464_wdata), .clk(f1464_clk), .rst(f1464_rst), .rdata(f1464_rdata));
  assign f1464_clk = clk;
  assign f1464_rst = rst;
  // Bindings to f1464

  // f1466
  logic [0:0] f1466_wen;
  logic [31:0] f1466_wdata;
  logic [0:0] f1466_clk;
  logic [0:0] f1466_rst;
  logic [31:0] f1466_rdata;
  sr_buffer_32_1 f1466(.wen(f1466_wen), .wdata(f1466_wdata), .clk(f1466_clk), .rst(f1466_rst), .rdata(f1466_rdata));
  assign f1466_clk = clk;
  assign f1466_rst = rst;
  // Bindings to f1466

  // f1468
  logic [0:0] f1468_wen;
  logic [31:0] f1468_wdata;
  logic [0:0] f1468_clk;
  logic [0:0] f1468_rst;
  logic [31:0] f1468_rdata;
  sr_buffer_32_1 f1468(.wen(f1468_wen), .wdata(f1468_wdata), .clk(f1468_clk), .rst(f1468_rst), .rdata(f1468_rdata));
  assign f1468_clk = clk;
  assign f1468_rst = rst;
  // Bindings to f1468

  // f1470
  logic [0:0] f1470_wen;
  logic [31:0] f1470_wdata;
  logic [0:0] f1470_clk;
  logic [0:0] f1470_rst;
  logic [31:0] f1470_rdata;
  sr_buffer_32_1 f1470(.wen(f1470_wen), .wdata(f1470_wdata), .clk(f1470_clk), .rst(f1470_rst), .rdata(f1470_rdata));
  assign f1470_clk = clk;
  assign f1470_rst = rst;
  // Bindings to f1470

  // f1472
  logic [0:0] f1472_wen;
  logic [31:0] f1472_wdata;
  logic [0:0] f1472_clk;
  logic [0:0] f1472_rst;
  logic [31:0] f1472_rdata;
  sr_buffer_32_1 f1472(.wen(f1472_wen), .wdata(f1472_wdata), .clk(f1472_clk), .rst(f1472_rst), .rdata(f1472_rdata));
  assign f1472_clk = clk;
  assign f1472_rst = rst;
  // Bindings to f1472

  // f1474
  logic [0:0] f1474_wen;
  logic [31:0] f1474_wdata;
  logic [0:0] f1474_clk;
  logic [0:0] f1474_rst;
  logic [31:0] f1474_rdata;
  sr_buffer_32_1 f1474(.wen(f1474_wen), .wdata(f1474_wdata), .clk(f1474_clk), .rst(f1474_rst), .rdata(f1474_rdata));
  assign f1474_clk = clk;
  assign f1474_rst = rst;
  // Bindings to f1474

  // f1476
  logic [0:0] f1476_wen;
  logic [31:0] f1476_wdata;
  logic [0:0] f1476_clk;
  logic [0:0] f1476_rst;
  logic [31:0] f1476_rdata;
  sr_buffer_32_1 f1476(.wen(f1476_wen), .wdata(f1476_wdata), .clk(f1476_clk), .rst(f1476_rst), .rdata(f1476_rdata));
  assign f1476_clk = clk;
  assign f1476_rst = rst;
  // Bindings to f1476

  // f1478
  logic [0:0] f1478_wen;
  logic [31:0] f1478_wdata;
  logic [0:0] f1478_clk;
  logic [0:0] f1478_rst;
  logic [31:0] f1478_rdata;
  sr_buffer_32_1 f1478(.wen(f1478_wen), .wdata(f1478_wdata), .clk(f1478_clk), .rst(f1478_rst), .rdata(f1478_rdata));
  assign f1478_clk = clk;
  assign f1478_rst = rst;
  // Bindings to f1478

  // f1480
  logic [0:0] f1480_wen;
  logic [31:0] f1480_wdata;
  logic [0:0] f1480_clk;
  logic [0:0] f1480_rst;
  logic [31:0] f1480_rdata;
  sr_buffer_32_1 f1480(.wen(f1480_wen), .wdata(f1480_wdata), .clk(f1480_clk), .rst(f1480_rst), .rdata(f1480_rdata));
  assign f1480_clk = clk;
  assign f1480_rst = rst;
  // Bindings to f1480

  // f1482
  logic [0:0] f1482_wen;
  logic [31:0] f1482_wdata;
  logic [0:0] f1482_clk;
  logic [0:0] f1482_rst;
  logic [31:0] f1482_rdata;
  sr_buffer_32_1 f1482(.wen(f1482_wen), .wdata(f1482_wdata), .clk(f1482_clk), .rst(f1482_rst), .rdata(f1482_rdata));
  assign f1482_clk = clk;
  assign f1482_rst = rst;
  // Bindings to f1482

  // f1484
  logic [0:0] f1484_wen;
  logic [31:0] f1484_wdata;
  logic [0:0] f1484_clk;
  logic [0:0] f1484_rst;
  logic [31:0] f1484_rdata;
  sr_buffer_32_1 f1484(.wen(f1484_wen), .wdata(f1484_wdata), .clk(f1484_clk), .rst(f1484_rst), .rdata(f1484_rdata));
  assign f1484_clk = clk;
  assign f1484_rst = rst;
  // Bindings to f1484

  // f1486
  logic [0:0] f1486_wen;
  logic [31:0] f1486_wdata;
  logic [0:0] f1486_clk;
  logic [0:0] f1486_rst;
  logic [31:0] f1486_rdata;
  sr_buffer_32_1 f1486(.wen(f1486_wen), .wdata(f1486_wdata), .clk(f1486_clk), .rst(f1486_rst), .rdata(f1486_rdata));
  assign f1486_clk = clk;
  assign f1486_rst = rst;
  // Bindings to f1486

  // f1488
  logic [0:0] f1488_wen;
  logic [31:0] f1488_wdata;
  logic [0:0] f1488_clk;
  logic [0:0] f1488_rst;
  logic [31:0] f1488_rdata;
  sr_buffer_32_1 f1488(.wen(f1488_wen), .wdata(f1488_wdata), .clk(f1488_clk), .rst(f1488_rst), .rdata(f1488_rdata));
  assign f1488_clk = clk;
  assign f1488_rst = rst;
  // Bindings to f1488

  // f1490
  logic [0:0] f1490_wen;
  logic [31:0] f1490_wdata;
  logic [0:0] f1490_clk;
  logic [0:0] f1490_rst;
  logic [31:0] f1490_rdata;
  sr_buffer_32_1 f1490(.wen(f1490_wen), .wdata(f1490_wdata), .clk(f1490_clk), .rst(f1490_rst), .rdata(f1490_rdata));
  assign f1490_clk = clk;
  assign f1490_rst = rst;
  // Bindings to f1490

  // f1492
  logic [0:0] f1492_wen;
  logic [31:0] f1492_wdata;
  logic [0:0] f1492_clk;
  logic [0:0] f1492_rst;
  logic [31:0] f1492_rdata;
  sr_buffer_32_1 f1492(.wen(f1492_wen), .wdata(f1492_wdata), .clk(f1492_clk), .rst(f1492_rst), .rdata(f1492_rdata));
  assign f1492_clk = clk;
  assign f1492_rst = rst;
  // Bindings to f1492

  // f1494
  logic [0:0] f1494_wen;
  logic [31:0] f1494_wdata;
  logic [0:0] f1494_clk;
  logic [0:0] f1494_rst;
  logic [31:0] f1494_rdata;
  sr_buffer_32_1 f1494(.wen(f1494_wen), .wdata(f1494_wdata), .clk(f1494_clk), .rst(f1494_rst), .rdata(f1494_rdata));
  assign f1494_clk = clk;
  assign f1494_rst = rst;
  // Bindings to f1494

  // f1496
  logic [0:0] f1496_wen;
  logic [31:0] f1496_wdata;
  logic [0:0] f1496_clk;
  logic [0:0] f1496_rst;
  logic [31:0] f1496_rdata;
  sr_buffer_32_1 f1496(.wen(f1496_wen), .wdata(f1496_wdata), .clk(f1496_clk), .rst(f1496_rst), .rdata(f1496_rdata));
  assign f1496_clk = clk;
  assign f1496_rst = rst;
  // Bindings to f1496

  // f1498
  logic [0:0] f1498_wen;
  logic [31:0] f1498_wdata;
  logic [0:0] f1498_clk;
  logic [0:0] f1498_rst;
  logic [31:0] f1498_rdata;
  sr_buffer_32_1 f1498(.wen(f1498_wen), .wdata(f1498_wdata), .clk(f1498_clk), .rst(f1498_rst), .rdata(f1498_rdata));
  assign f1498_clk = clk;
  assign f1498_rst = rst;
  // Bindings to f1498

  // f1500
  logic [0:0] f1500_wen;
  logic [31:0] f1500_wdata;
  logic [0:0] f1500_clk;
  logic [0:0] f1500_rst;
  logic [31:0] f1500_rdata;
  sr_buffer_32_1 f1500(.wen(f1500_wen), .wdata(f1500_wdata), .clk(f1500_clk), .rst(f1500_rst), .rdata(f1500_rdata));
  assign f1500_clk = clk;
  assign f1500_rst = rst;
  // Bindings to f1500

  // f1502
  logic [0:0] f1502_wen;
  logic [31:0] f1502_wdata;
  logic [0:0] f1502_clk;
  logic [0:0] f1502_rst;
  logic [31:0] f1502_rdata;
  sr_buffer_32_1 f1502(.wen(f1502_wen), .wdata(f1502_wdata), .clk(f1502_clk), .rst(f1502_rst), .rdata(f1502_rdata));
  assign f1502_clk = clk;
  assign f1502_rst = rst;
  // Bindings to f1502

  // f1504
  logic [0:0] f1504_wen;
  logic [31:0] f1504_wdata;
  logic [0:0] f1504_clk;
  logic [0:0] f1504_rst;
  logic [31:0] f1504_rdata;
  sr_buffer_32_1 f1504(.wen(f1504_wen), .wdata(f1504_wdata), .clk(f1504_clk), .rst(f1504_rst), .rdata(f1504_rdata));
  assign f1504_clk = clk;
  assign f1504_rst = rst;
  // Bindings to f1504

  // f1506
  logic [0:0] f1506_wen;
  logic [31:0] f1506_wdata;
  logic [0:0] f1506_clk;
  logic [0:0] f1506_rst;
  logic [31:0] f1506_rdata;
  sr_buffer_32_1 f1506(.wen(f1506_wen), .wdata(f1506_wdata), .clk(f1506_clk), .rst(f1506_rst), .rdata(f1506_rdata));
  assign f1506_clk = clk;
  assign f1506_rst = rst;
  // Bindings to f1506

  // f1508
  logic [0:0] f1508_wen;
  logic [31:0] f1508_wdata;
  logic [0:0] f1508_clk;
  logic [0:0] f1508_rst;
  logic [31:0] f1508_rdata;
  sr_buffer_32_1 f1508(.wen(f1508_wen), .wdata(f1508_wdata), .clk(f1508_clk), .rst(f1508_rst), .rdata(f1508_rdata));
  assign f1508_clk = clk;
  assign f1508_rst = rst;
  // Bindings to f1508

  // f1510
  logic [0:0] f1510_wen;
  logic [31:0] f1510_wdata;
  logic [0:0] f1510_clk;
  logic [0:0] f1510_rst;
  logic [31:0] f1510_rdata;
  sr_buffer_32_1 f1510(.wen(f1510_wen), .wdata(f1510_wdata), .clk(f1510_clk), .rst(f1510_rst), .rdata(f1510_rdata));
  assign f1510_clk = clk;
  assign f1510_rst = rst;
  // Bindings to f1510

  // f1512
  logic [0:0] f1512_wen;
  logic [31:0] f1512_wdata;
  logic [0:0] f1512_clk;
  logic [0:0] f1512_rst;
  logic [31:0] f1512_rdata;
  sr_buffer_32_1 f1512(.wen(f1512_wen), .wdata(f1512_wdata), .clk(f1512_clk), .rst(f1512_rst), .rdata(f1512_rdata));
  assign f1512_clk = clk;
  assign f1512_rst = rst;
  // Bindings to f1512

  // f1514
  logic [0:0] f1514_wen;
  logic [31:0] f1514_wdata;
  logic [0:0] f1514_clk;
  logic [0:0] f1514_rst;
  logic [31:0] f1514_rdata;
  sr_buffer_32_1 f1514(.wen(f1514_wen), .wdata(f1514_wdata), .clk(f1514_clk), .rst(f1514_rst), .rdata(f1514_rdata));
  assign f1514_clk = clk;
  assign f1514_rst = rst;
  // Bindings to f1514

  // f1516
  logic [0:0] f1516_wen;
  logic [31:0] f1516_wdata;
  logic [0:0] f1516_clk;
  logic [0:0] f1516_rst;
  logic [31:0] f1516_rdata;
  sr_buffer_32_1 f1516(.wen(f1516_wen), .wdata(f1516_wdata), .clk(f1516_clk), .rst(f1516_rst), .rdata(f1516_rdata));
  assign f1516_clk = clk;
  assign f1516_rst = rst;
  // Bindings to f1516

  // f1518
  logic [0:0] f1518_wen;
  logic [31:0] f1518_wdata;
  logic [0:0] f1518_clk;
  logic [0:0] f1518_rst;
  logic [31:0] f1518_rdata;
  sr_buffer_32_1 f1518(.wen(f1518_wen), .wdata(f1518_wdata), .clk(f1518_clk), .rst(f1518_rst), .rdata(f1518_rdata));
  assign f1518_clk = clk;
  assign f1518_rst = rst;
  // Bindings to f1518

  // f1520
  logic [0:0] f1520_wen;
  logic [31:0] f1520_wdata;
  logic [0:0] f1520_clk;
  logic [0:0] f1520_rst;
  logic [31:0] f1520_rdata;
  sr_buffer_32_1 f1520(.wen(f1520_wen), .wdata(f1520_wdata), .clk(f1520_clk), .rst(f1520_rst), .rdata(f1520_rdata));
  assign f1520_clk = clk;
  assign f1520_rst = rst;
  // Bindings to f1520

  // f1522
  logic [0:0] f1522_wen;
  logic [31:0] f1522_wdata;
  logic [0:0] f1522_clk;
  logic [0:0] f1522_rst;
  logic [31:0] f1522_rdata;
  sr_buffer_32_1 f1522(.wen(f1522_wen), .wdata(f1522_wdata), .clk(f1522_clk), .rst(f1522_rst), .rdata(f1522_rdata));
  assign f1522_clk = clk;
  assign f1522_rst = rst;
  // Bindings to f1522

  // f1524
  logic [0:0] f1524_wen;
  logic [31:0] f1524_wdata;
  logic [0:0] f1524_clk;
  logic [0:0] f1524_rst;
  logic [31:0] f1524_rdata;
  sr_buffer_32_1 f1524(.wen(f1524_wen), .wdata(f1524_wdata), .clk(f1524_clk), .rst(f1524_rst), .rdata(f1524_rdata));
  assign f1524_clk = clk;
  assign f1524_rst = rst;
  // Bindings to f1524

  // f1526
  logic [0:0] f1526_wen;
  logic [31:0] f1526_wdata;
  logic [0:0] f1526_clk;
  logic [0:0] f1526_rst;
  logic [31:0] f1526_rdata;
  sr_buffer_32_1 f1526(.wen(f1526_wen), .wdata(f1526_wdata), .clk(f1526_clk), .rst(f1526_rst), .rdata(f1526_rdata));
  assign f1526_clk = clk;
  assign f1526_rst = rst;
  // Bindings to f1526

  // f1528
  logic [0:0] f1528_wen;
  logic [31:0] f1528_wdata;
  logic [0:0] f1528_clk;
  logic [0:0] f1528_rst;
  logic [31:0] f1528_rdata;
  sr_buffer_32_1 f1528(.wen(f1528_wen), .wdata(f1528_wdata), .clk(f1528_clk), .rst(f1528_rst), .rdata(f1528_rdata));
  assign f1528_clk = clk;
  assign f1528_rst = rst;
  // Bindings to f1528

  // f1530
  logic [0:0] f1530_wen;
  logic [31:0] f1530_wdata;
  logic [0:0] f1530_clk;
  logic [0:0] f1530_rst;
  logic [31:0] f1530_rdata;
  sr_buffer_32_1 f1530(.wen(f1530_wen), .wdata(f1530_wdata), .clk(f1530_clk), .rst(f1530_rst), .rdata(f1530_rdata));
  assign f1530_clk = clk;
  assign f1530_rst = rst;
  // Bindings to f1530

  // f1532
  logic [0:0] f1532_wen;
  logic [31:0] f1532_wdata;
  logic [0:0] f1532_clk;
  logic [0:0] f1532_rst;
  logic [31:0] f1532_rdata;
  sr_buffer_32_1 f1532(.wen(f1532_wen), .wdata(f1532_wdata), .clk(f1532_clk), .rst(f1532_rst), .rdata(f1532_rdata));
  assign f1532_clk = clk;
  assign f1532_rst = rst;
  // Bindings to f1532

  // f1534
  logic [0:0] f1534_wen;
  logic [31:0] f1534_wdata;
  logic [0:0] f1534_clk;
  logic [0:0] f1534_rst;
  logic [31:0] f1534_rdata;
  sr_buffer_32_1 f1534(.wen(f1534_wen), .wdata(f1534_wdata), .clk(f1534_clk), .rst(f1534_rst), .rdata(f1534_rdata));
  assign f1534_clk = clk;
  assign f1534_rst = rst;
  // Bindings to f1534

  // f1536
  logic [0:0] f1536_wen;
  logic [31:0] f1536_wdata;
  logic [0:0] f1536_clk;
  logic [0:0] f1536_rst;
  logic [31:0] f1536_rdata;
  sr_buffer_32_1 f1536(.wen(f1536_wen), .wdata(f1536_wdata), .clk(f1536_clk), .rst(f1536_rst), .rdata(f1536_rdata));
  assign f1536_clk = clk;
  assign f1536_rst = rst;
  // Bindings to f1536

  // f1538
  logic [0:0] f1538_wen;
  logic [31:0] f1538_wdata;
  logic [0:0] f1538_clk;
  logic [0:0] f1538_rst;
  logic [31:0] f1538_rdata;
  sr_buffer_32_1 f1538(.wen(f1538_wen), .wdata(f1538_wdata), .clk(f1538_clk), .rst(f1538_rst), .rdata(f1538_rdata));
  assign f1538_clk = clk;
  assign f1538_rst = rst;
  // Bindings to f1538

  // f1540
  logic [0:0] f1540_wen;
  logic [31:0] f1540_wdata;
  logic [0:0] f1540_clk;
  logic [0:0] f1540_rst;
  logic [31:0] f1540_rdata;
  sr_buffer_32_1 f1540(.wen(f1540_wen), .wdata(f1540_wdata), .clk(f1540_clk), .rst(f1540_rst), .rdata(f1540_rdata));
  assign f1540_clk = clk;
  assign f1540_rst = rst;
  // Bindings to f1540

  // f1542
  logic [0:0] f1542_wen;
  logic [31:0] f1542_wdata;
  logic [0:0] f1542_clk;
  logic [0:0] f1542_rst;
  logic [31:0] f1542_rdata;
  sr_buffer_32_1 f1542(.wen(f1542_wen), .wdata(f1542_wdata), .clk(f1542_clk), .rst(f1542_rst), .rdata(f1542_rdata));
  assign f1542_clk = clk;
  assign f1542_rst = rst;
  // Bindings to f1542

  // f1544
  logic [0:0] f1544_wen;
  logic [31:0] f1544_wdata;
  logic [0:0] f1544_clk;
  logic [0:0] f1544_rst;
  logic [31:0] f1544_rdata;
  sr_buffer_32_1 f1544(.wen(f1544_wen), .wdata(f1544_wdata), .clk(f1544_clk), .rst(f1544_rst), .rdata(f1544_rdata));
  assign f1544_clk = clk;
  assign f1544_rst = rst;
  // Bindings to f1544

  // f1546
  logic [0:0] f1546_wen;
  logic [31:0] f1546_wdata;
  logic [0:0] f1546_clk;
  logic [0:0] f1546_rst;
  logic [31:0] f1546_rdata;
  sr_buffer_32_1 f1546(.wen(f1546_wen), .wdata(f1546_wdata), .clk(f1546_clk), .rst(f1546_rst), .rdata(f1546_rdata));
  assign f1546_clk = clk;
  assign f1546_rst = rst;
  // Bindings to f1546

  // f1548
  logic [0:0] f1548_wen;
  logic [31:0] f1548_wdata;
  logic [0:0] f1548_clk;
  logic [0:0] f1548_rst;
  logic [31:0] f1548_rdata;
  sr_buffer_32_1 f1548(.wen(f1548_wen), .wdata(f1548_wdata), .clk(f1548_clk), .rst(f1548_rst), .rdata(f1548_rdata));
  assign f1548_clk = clk;
  assign f1548_rst = rst;
  // Bindings to f1548

  // f1550
  logic [0:0] f1550_wen;
  logic [31:0] f1550_wdata;
  logic [0:0] f1550_clk;
  logic [0:0] f1550_rst;
  logic [31:0] f1550_rdata;
  sr_buffer_32_1 f1550(.wen(f1550_wen), .wdata(f1550_wdata), .clk(f1550_clk), .rst(f1550_rst), .rdata(f1550_rdata));
  assign f1550_clk = clk;
  assign f1550_rst = rst;
  // Bindings to f1550

  // f1552
  logic [0:0] f1552_wen;
  logic [31:0] f1552_wdata;
  logic [0:0] f1552_clk;
  logic [0:0] f1552_rst;
  logic [31:0] f1552_rdata;
  sr_buffer_32_1 f1552(.wen(f1552_wen), .wdata(f1552_wdata), .clk(f1552_clk), .rst(f1552_rst), .rdata(f1552_rdata));
  assign f1552_clk = clk;
  assign f1552_rst = rst;
  // Bindings to f1552

  // f1554
  logic [0:0] f1554_wen;
  logic [31:0] f1554_wdata;
  logic [0:0] f1554_clk;
  logic [0:0] f1554_rst;
  logic [31:0] f1554_rdata;
  sr_buffer_32_1 f1554(.wen(f1554_wen), .wdata(f1554_wdata), .clk(f1554_clk), .rst(f1554_rst), .rdata(f1554_rdata));
  assign f1554_clk = clk;
  assign f1554_rst = rst;
  // Bindings to f1554

  // f1556
  logic [0:0] f1556_wen;
  logic [31:0] f1556_wdata;
  logic [0:0] f1556_clk;
  logic [0:0] f1556_rst;
  logic [31:0] f1556_rdata;
  sr_buffer_32_1 f1556(.wen(f1556_wen), .wdata(f1556_wdata), .clk(f1556_clk), .rst(f1556_rst), .rdata(f1556_rdata));
  assign f1556_clk = clk;
  assign f1556_rst = rst;
  // Bindings to f1556

  // f1558
  logic [0:0] f1558_wen;
  logic [31:0] f1558_wdata;
  logic [0:0] f1558_clk;
  logic [0:0] f1558_rst;
  logic [31:0] f1558_rdata;
  sr_buffer_32_1 f1558(.wen(f1558_wen), .wdata(f1558_wdata), .clk(f1558_clk), .rst(f1558_rst), .rdata(f1558_rdata));
  assign f1558_clk = clk;
  assign f1558_rst = rst;
  // Bindings to f1558

  // f1560
  logic [0:0] f1560_wen;
  logic [31:0] f1560_wdata;
  logic [0:0] f1560_clk;
  logic [0:0] f1560_rst;
  logic [31:0] f1560_rdata;
  sr_buffer_32_1 f1560(.wen(f1560_wen), .wdata(f1560_wdata), .clk(f1560_clk), .rst(f1560_rst), .rdata(f1560_rdata));
  assign f1560_clk = clk;
  assign f1560_rst = rst;
  // Bindings to f1560

  // f1562
  logic [0:0] f1562_wen;
  logic [31:0] f1562_wdata;
  logic [0:0] f1562_clk;
  logic [0:0] f1562_rst;
  logic [31:0] f1562_rdata;
  sr_buffer_32_1 f1562(.wen(f1562_wen), .wdata(f1562_wdata), .clk(f1562_clk), .rst(f1562_rst), .rdata(f1562_rdata));
  assign f1562_clk = clk;
  assign f1562_rst = rst;
  // Bindings to f1562

  // f1564
  logic [0:0] f1564_wen;
  logic [31:0] f1564_wdata;
  logic [0:0] f1564_clk;
  logic [0:0] f1564_rst;
  logic [31:0] f1564_rdata;
  sr_buffer_32_1 f1564(.wen(f1564_wen), .wdata(f1564_wdata), .clk(f1564_clk), .rst(f1564_rst), .rdata(f1564_rdata));
  assign f1564_clk = clk;
  assign f1564_rst = rst;
  // Bindings to f1564

  // f1566
  logic [0:0] f1566_wen;
  logic [31:0] f1566_wdata;
  logic [0:0] f1566_clk;
  logic [0:0] f1566_rst;
  logic [31:0] f1566_rdata;
  sr_buffer_32_1 f1566(.wen(f1566_wen), .wdata(f1566_wdata), .clk(f1566_clk), .rst(f1566_rst), .rdata(f1566_rdata));
  assign f1566_clk = clk;
  assign f1566_rst = rst;
  // Bindings to f1566

  // f1568
  logic [0:0] f1568_wen;
  logic [31:0] f1568_wdata;
  logic [0:0] f1568_clk;
  logic [0:0] f1568_rst;
  logic [31:0] f1568_rdata;
  sr_buffer_32_1 f1568(.wen(f1568_wen), .wdata(f1568_wdata), .clk(f1568_clk), .rst(f1568_rst), .rdata(f1568_rdata));
  assign f1568_clk = clk;
  assign f1568_rst = rst;
  // Bindings to f1568

  // f1570
  logic [0:0] f1570_wen;
  logic [31:0] f1570_wdata;
  logic [0:0] f1570_clk;
  logic [0:0] f1570_rst;
  logic [31:0] f1570_rdata;
  sr_buffer_32_1 f1570(.wen(f1570_wen), .wdata(f1570_wdata), .clk(f1570_clk), .rst(f1570_rst), .rdata(f1570_rdata));
  assign f1570_clk = clk;
  assign f1570_rst = rst;
  // Bindings to f1570

  // f1572
  logic [0:0] f1572_wen;
  logic [31:0] f1572_wdata;
  logic [0:0] f1572_clk;
  logic [0:0] f1572_rst;
  logic [31:0] f1572_rdata;
  sr_buffer_32_1 f1572(.wen(f1572_wen), .wdata(f1572_wdata), .clk(f1572_clk), .rst(f1572_rst), .rdata(f1572_rdata));
  assign f1572_clk = clk;
  assign f1572_rst = rst;
  // Bindings to f1572

  // f1574
  logic [0:0] f1574_wen;
  logic [31:0] f1574_wdata;
  logic [0:0] f1574_clk;
  logic [0:0] f1574_rst;
  logic [31:0] f1574_rdata;
  sr_buffer_32_1 f1574(.wen(f1574_wen), .wdata(f1574_wdata), .clk(f1574_clk), .rst(f1574_rst), .rdata(f1574_rdata));
  assign f1574_clk = clk;
  assign f1574_rst = rst;
  // Bindings to f1574

  // f1576
  logic [0:0] f1576_wen;
  logic [31:0] f1576_wdata;
  logic [0:0] f1576_clk;
  logic [0:0] f1576_rst;
  logic [31:0] f1576_rdata;
  sr_buffer_32_1 f1576(.wen(f1576_wen), .wdata(f1576_wdata), .clk(f1576_clk), .rst(f1576_rst), .rdata(f1576_rdata));
  assign f1576_clk = clk;
  assign f1576_rst = rst;
  // Bindings to f1576

  // f1578
  logic [0:0] f1578_wen;
  logic [31:0] f1578_wdata;
  logic [0:0] f1578_clk;
  logic [0:0] f1578_rst;
  logic [31:0] f1578_rdata;
  sr_buffer_32_1 f1578(.wen(f1578_wen), .wdata(f1578_wdata), .clk(f1578_clk), .rst(f1578_rst), .rdata(f1578_rdata));
  assign f1578_clk = clk;
  assign f1578_rst = rst;
  // Bindings to f1578

  // f1580
  logic [0:0] f1580_wen;
  logic [31:0] f1580_wdata;
  logic [0:0] f1580_clk;
  logic [0:0] f1580_rst;
  logic [31:0] f1580_rdata;
  sr_buffer_32_1 f1580(.wen(f1580_wen), .wdata(f1580_wdata), .clk(f1580_clk), .rst(f1580_rst), .rdata(f1580_rdata));
  assign f1580_clk = clk;
  assign f1580_rst = rst;
  // Bindings to f1580

  // f1582
  logic [0:0] f1582_wen;
  logic [31:0] f1582_wdata;
  logic [0:0] f1582_clk;
  logic [0:0] f1582_rst;
  logic [31:0] f1582_rdata;
  sr_buffer_32_1 f1582(.wen(f1582_wen), .wdata(f1582_wdata), .clk(f1582_clk), .rst(f1582_rst), .rdata(f1582_rdata));
  assign f1582_clk = clk;
  assign f1582_rst = rst;
  // Bindings to f1582

  // f1584
  logic [0:0] f1584_wen;
  logic [31:0] f1584_wdata;
  logic [0:0] f1584_clk;
  logic [0:0] f1584_rst;
  logic [31:0] f1584_rdata;
  sr_buffer_32_1 f1584(.wen(f1584_wen), .wdata(f1584_wdata), .clk(f1584_clk), .rst(f1584_rst), .rdata(f1584_rdata));
  assign f1584_clk = clk;
  assign f1584_rst = rst;
  // Bindings to f1584

  // f1586
  logic [0:0] f1586_wen;
  logic [31:0] f1586_wdata;
  logic [0:0] f1586_clk;
  logic [0:0] f1586_rst;
  logic [31:0] f1586_rdata;
  sr_buffer_32_1 f1586(.wen(f1586_wen), .wdata(f1586_wdata), .clk(f1586_clk), .rst(f1586_rst), .rdata(f1586_rdata));
  assign f1586_clk = clk;
  assign f1586_rst = rst;
  // Bindings to f1586

  // f1588
  logic [0:0] f1588_wen;
  logic [31:0] f1588_wdata;
  logic [0:0] f1588_clk;
  logic [0:0] f1588_rst;
  logic [31:0] f1588_rdata;
  sr_buffer_32_1 f1588(.wen(f1588_wen), .wdata(f1588_wdata), .clk(f1588_clk), .rst(f1588_rst), .rdata(f1588_rdata));
  assign f1588_clk = clk;
  assign f1588_rst = rst;
  // Bindings to f1588

  // f1590
  logic [0:0] f1590_wen;
  logic [31:0] f1590_wdata;
  logic [0:0] f1590_clk;
  logic [0:0] f1590_rst;
  logic [31:0] f1590_rdata;
  sr_buffer_32_1 f1590(.wen(f1590_wen), .wdata(f1590_wdata), .clk(f1590_clk), .rst(f1590_rst), .rdata(f1590_rdata));
  assign f1590_clk = clk;
  assign f1590_rst = rst;
  // Bindings to f1590

  // f1592
  logic [0:0] f1592_wen;
  logic [31:0] f1592_wdata;
  logic [0:0] f1592_clk;
  logic [0:0] f1592_rst;
  logic [31:0] f1592_rdata;
  sr_buffer_32_1 f1592(.wen(f1592_wen), .wdata(f1592_wdata), .clk(f1592_clk), .rst(f1592_rst), .rdata(f1592_rdata));
  assign f1592_clk = clk;
  assign f1592_rst = rst;
  // Bindings to f1592

  // f1594
  logic [0:0] f1594_wen;
  logic [31:0] f1594_wdata;
  logic [0:0] f1594_clk;
  logic [0:0] f1594_rst;
  logic [31:0] f1594_rdata;
  sr_buffer_32_1 f1594(.wen(f1594_wen), .wdata(f1594_wdata), .clk(f1594_clk), .rst(f1594_rst), .rdata(f1594_rdata));
  assign f1594_clk = clk;
  assign f1594_rst = rst;
  // Bindings to f1594

  // f1596
  logic [0:0] f1596_wen;
  logic [31:0] f1596_wdata;
  logic [0:0] f1596_clk;
  logic [0:0] f1596_rst;
  logic [31:0] f1596_rdata;
  sr_buffer_32_1 f1596(.wen(f1596_wen), .wdata(f1596_wdata), .clk(f1596_clk), .rst(f1596_rst), .rdata(f1596_rdata));
  assign f1596_clk = clk;
  assign f1596_rst = rst;
  // Bindings to f1596

  // f1598
  logic [0:0] f1598_wen;
  logic [31:0] f1598_wdata;
  logic [0:0] f1598_clk;
  logic [0:0] f1598_rst;
  logic [31:0] f1598_rdata;
  sr_buffer_32_1 f1598(.wen(f1598_wen), .wdata(f1598_wdata), .clk(f1598_clk), .rst(f1598_rst), .rdata(f1598_rdata));
  assign f1598_clk = clk;
  assign f1598_rst = rst;
  // Bindings to f1598

  // f1600
  logic [0:0] f1600_wen;
  logic [31:0] f1600_wdata;
  logic [0:0] f1600_clk;
  logic [0:0] f1600_rst;
  logic [31:0] f1600_rdata;
  sr_buffer_32_1 f1600(.wen(f1600_wen), .wdata(f1600_wdata), .clk(f1600_clk), .rst(f1600_rst), .rdata(f1600_rdata));
  assign f1600_clk = clk;
  assign f1600_rst = rst;
  // Bindings to f1600

  // f1602
  logic [0:0] f1602_wen;
  logic [31:0] f1602_wdata;
  logic [0:0] f1602_clk;
  logic [0:0] f1602_rst;
  logic [31:0] f1602_rdata;
  sr_buffer_32_1 f1602(.wen(f1602_wen), .wdata(f1602_wdata), .clk(f1602_clk), .rst(f1602_rst), .rdata(f1602_rdata));
  assign f1602_clk = clk;
  assign f1602_rst = rst;
  // Bindings to f1602

  // f1604
  logic [0:0] f1604_wen;
  logic [31:0] f1604_wdata;
  logic [0:0] f1604_clk;
  logic [0:0] f1604_rst;
  logic [31:0] f1604_rdata;
  sr_buffer_32_1 f1604(.wen(f1604_wen), .wdata(f1604_wdata), .clk(f1604_clk), .rst(f1604_rst), .rdata(f1604_rdata));
  assign f1604_clk = clk;
  assign f1604_rst = rst;
  // Bindings to f1604

  // f1606
  logic [0:0] f1606_wen;
  logic [31:0] f1606_wdata;
  logic [0:0] f1606_clk;
  logic [0:0] f1606_rst;
  logic [31:0] f1606_rdata;
  sr_buffer_32_1 f1606(.wen(f1606_wen), .wdata(f1606_wdata), .clk(f1606_clk), .rst(f1606_rst), .rdata(f1606_rdata));
  assign f1606_clk = clk;
  assign f1606_rst = rst;
  // Bindings to f1606

  // f1608
  logic [0:0] f1608_wen;
  logic [31:0] f1608_wdata;
  logic [0:0] f1608_clk;
  logic [0:0] f1608_rst;
  logic [31:0] f1608_rdata;
  sr_buffer_32_1 f1608(.wen(f1608_wen), .wdata(f1608_wdata), .clk(f1608_clk), .rst(f1608_rst), .rdata(f1608_rdata));
  assign f1608_clk = clk;
  assign f1608_rst = rst;
  // Bindings to f1608

  // f1610
  logic [0:0] f1610_wen;
  logic [31:0] f1610_wdata;
  logic [0:0] f1610_clk;
  logic [0:0] f1610_rst;
  logic [31:0] f1610_rdata;
  sr_buffer_32_1 f1610(.wen(f1610_wen), .wdata(f1610_wdata), .clk(f1610_clk), .rst(f1610_rst), .rdata(f1610_rdata));
  assign f1610_clk = clk;
  assign f1610_rst = rst;
  // Bindings to f1610

  // f1612
  logic [0:0] f1612_wen;
  logic [31:0] f1612_wdata;
  logic [0:0] f1612_clk;
  logic [0:0] f1612_rst;
  logic [31:0] f1612_rdata;
  sr_buffer_32_1 f1612(.wen(f1612_wen), .wdata(f1612_wdata), .clk(f1612_clk), .rst(f1612_rst), .rdata(f1612_rdata));
  assign f1612_clk = clk;
  assign f1612_rst = rst;
  // Bindings to f1612

  // f1614
  logic [0:0] f1614_wen;
  logic [31:0] f1614_wdata;
  logic [0:0] f1614_clk;
  logic [0:0] f1614_rst;
  logic [31:0] f1614_rdata;
  sr_buffer_32_1 f1614(.wen(f1614_wen), .wdata(f1614_wdata), .clk(f1614_clk), .rst(f1614_rst), .rdata(f1614_rdata));
  assign f1614_clk = clk;
  assign f1614_rst = rst;
  // Bindings to f1614

  // f1616
  logic [0:0] f1616_wen;
  logic [31:0] f1616_wdata;
  logic [0:0] f1616_clk;
  logic [0:0] f1616_rst;
  logic [31:0] f1616_rdata;
  sr_buffer_32_1 f1616(.wen(f1616_wen), .wdata(f1616_wdata), .clk(f1616_clk), .rst(f1616_rst), .rdata(f1616_rdata));
  assign f1616_clk = clk;
  assign f1616_rst = rst;
  // Bindings to f1616

  // f1618
  logic [0:0] f1618_wen;
  logic [31:0] f1618_wdata;
  logic [0:0] f1618_clk;
  logic [0:0] f1618_rst;
  logic [31:0] f1618_rdata;
  sr_buffer_32_1 f1618(.wen(f1618_wen), .wdata(f1618_wdata), .clk(f1618_clk), .rst(f1618_rst), .rdata(f1618_rdata));
  assign f1618_clk = clk;
  assign f1618_rst = rst;
  // Bindings to f1618

  // f1620
  logic [0:0] f1620_wen;
  logic [31:0] f1620_wdata;
  logic [0:0] f1620_clk;
  logic [0:0] f1620_rst;
  logic [31:0] f1620_rdata;
  sr_buffer_32_1 f1620(.wen(f1620_wen), .wdata(f1620_wdata), .clk(f1620_clk), .rst(f1620_rst), .rdata(f1620_rdata));
  assign f1620_clk = clk;
  assign f1620_rst = rst;
  // Bindings to f1620

  // f1622
  logic [0:0] f1622_wen;
  logic [31:0] f1622_wdata;
  logic [0:0] f1622_clk;
  logic [0:0] f1622_rst;
  logic [31:0] f1622_rdata;
  sr_buffer_32_1 f1622(.wen(f1622_wen), .wdata(f1622_wdata), .clk(f1622_clk), .rst(f1622_rst), .rdata(f1622_rdata));
  assign f1622_clk = clk;
  assign f1622_rst = rst;
  // Bindings to f1622

  // f1624
  logic [0:0] f1624_wen;
  logic [31:0] f1624_wdata;
  logic [0:0] f1624_clk;
  logic [0:0] f1624_rst;
  logic [31:0] f1624_rdata;
  sr_buffer_32_1 f1624(.wen(f1624_wen), .wdata(f1624_wdata), .clk(f1624_clk), .rst(f1624_rst), .rdata(f1624_rdata));
  assign f1624_clk = clk;
  assign f1624_rst = rst;
  // Bindings to f1624

  // f1626
  logic [0:0] f1626_wen;
  logic [31:0] f1626_wdata;
  logic [0:0] f1626_clk;
  logic [0:0] f1626_rst;
  logic [31:0] f1626_rdata;
  sr_buffer_32_1 f1626(.wen(f1626_wen), .wdata(f1626_wdata), .clk(f1626_clk), .rst(f1626_rst), .rdata(f1626_rdata));
  assign f1626_clk = clk;
  assign f1626_rst = rst;
  // Bindings to f1626

  // f1628
  logic [0:0] f1628_wen;
  logic [31:0] f1628_wdata;
  logic [0:0] f1628_clk;
  logic [0:0] f1628_rst;
  logic [31:0] f1628_rdata;
  sr_buffer_32_1 f1628(.wen(f1628_wen), .wdata(f1628_wdata), .clk(f1628_clk), .rst(f1628_rst), .rdata(f1628_rdata));
  assign f1628_clk = clk;
  assign f1628_rst = rst;
  // Bindings to f1628

  // f1630
  logic [0:0] f1630_wen;
  logic [31:0] f1630_wdata;
  logic [0:0] f1630_clk;
  logic [0:0] f1630_rst;
  logic [31:0] f1630_rdata;
  sr_buffer_32_1 f1630(.wen(f1630_wen), .wdata(f1630_wdata), .clk(f1630_clk), .rst(f1630_rst), .rdata(f1630_rdata));
  assign f1630_clk = clk;
  assign f1630_rst = rst;
  // Bindings to f1630

  // f1632
  logic [0:0] f1632_wen;
  logic [31:0] f1632_wdata;
  logic [0:0] f1632_clk;
  logic [0:0] f1632_rst;
  logic [31:0] f1632_rdata;
  sr_buffer_32_1 f1632(.wen(f1632_wen), .wdata(f1632_wdata), .clk(f1632_clk), .rst(f1632_rst), .rdata(f1632_rdata));
  assign f1632_clk = clk;
  assign f1632_rst = rst;
  // Bindings to f1632

  // f1634
  logic [0:0] f1634_wen;
  logic [31:0] f1634_wdata;
  logic [0:0] f1634_clk;
  logic [0:0] f1634_rst;
  logic [31:0] f1634_rdata;
  sr_buffer_32_1 f1634(.wen(f1634_wen), .wdata(f1634_wdata), .clk(f1634_clk), .rst(f1634_rst), .rdata(f1634_rdata));
  assign f1634_clk = clk;
  assign f1634_rst = rst;
  // Bindings to f1634

  // f1636
  logic [0:0] f1636_wen;
  logic [31:0] f1636_wdata;
  logic [0:0] f1636_clk;
  logic [0:0] f1636_rst;
  logic [31:0] f1636_rdata;
  sr_buffer_32_1 f1636(.wen(f1636_wen), .wdata(f1636_wdata), .clk(f1636_clk), .rst(f1636_rst), .rdata(f1636_rdata));
  assign f1636_clk = clk;
  assign f1636_rst = rst;
  // Bindings to f1636

  // f1638
  logic [0:0] f1638_wen;
  logic [31:0] f1638_wdata;
  logic [0:0] f1638_clk;
  logic [0:0] f1638_rst;
  logic [31:0] f1638_rdata;
  sr_buffer_32_1 f1638(.wen(f1638_wen), .wdata(f1638_wdata), .clk(f1638_clk), .rst(f1638_rst), .rdata(f1638_rdata));
  assign f1638_clk = clk;
  assign f1638_rst = rst;
  // Bindings to f1638

  // f1640
  logic [0:0] f1640_wen;
  logic [31:0] f1640_wdata;
  logic [0:0] f1640_clk;
  logic [0:0] f1640_rst;
  logic [31:0] f1640_rdata;
  sr_buffer_32_1 f1640(.wen(f1640_wen), .wdata(f1640_wdata), .clk(f1640_clk), .rst(f1640_rst), .rdata(f1640_rdata));
  assign f1640_clk = clk;
  assign f1640_rst = rst;
  // Bindings to f1640

  // f1642
  logic [0:0] f1642_wen;
  logic [31:0] f1642_wdata;
  logic [0:0] f1642_clk;
  logic [0:0] f1642_rst;
  logic [31:0] f1642_rdata;
  sr_buffer_32_1 f1642(.wen(f1642_wen), .wdata(f1642_wdata), .clk(f1642_clk), .rst(f1642_rst), .rdata(f1642_rdata));
  assign f1642_clk = clk;
  assign f1642_rst = rst;
  // Bindings to f1642

  // f1644
  logic [0:0] f1644_wen;
  logic [31:0] f1644_wdata;
  logic [0:0] f1644_clk;
  logic [0:0] f1644_rst;
  logic [31:0] f1644_rdata;
  sr_buffer_32_1 f1644(.wen(f1644_wen), .wdata(f1644_wdata), .clk(f1644_clk), .rst(f1644_rst), .rdata(f1644_rdata));
  assign f1644_clk = clk;
  assign f1644_rst = rst;
  // Bindings to f1644

  // f1646
  logic [0:0] f1646_wen;
  logic [31:0] f1646_wdata;
  logic [0:0] f1646_clk;
  logic [0:0] f1646_rst;
  logic [31:0] f1646_rdata;
  sr_buffer_32_1 f1646(.wen(f1646_wen), .wdata(f1646_wdata), .clk(f1646_clk), .rst(f1646_rst), .rdata(f1646_rdata));
  assign f1646_clk = clk;
  assign f1646_rst = rst;
  // Bindings to f1646

  // f1648
  logic [0:0] f1648_wen;
  logic [31:0] f1648_wdata;
  logic [0:0] f1648_clk;
  logic [0:0] f1648_rst;
  logic [31:0] f1648_rdata;
  sr_buffer_32_1 f1648(.wen(f1648_wen), .wdata(f1648_wdata), .clk(f1648_clk), .rst(f1648_rst), .rdata(f1648_rdata));
  assign f1648_clk = clk;
  assign f1648_rst = rst;
  // Bindings to f1648

  // f1650
  logic [0:0] f1650_wen;
  logic [31:0] f1650_wdata;
  logic [0:0] f1650_clk;
  logic [0:0] f1650_rst;
  logic [31:0] f1650_rdata;
  sr_buffer_32_1 f1650(.wen(f1650_wen), .wdata(f1650_wdata), .clk(f1650_clk), .rst(f1650_rst), .rdata(f1650_rdata));
  assign f1650_clk = clk;
  assign f1650_rst = rst;
  // Bindings to f1650

  // f1652
  logic [0:0] f1652_wen;
  logic [31:0] f1652_wdata;
  logic [0:0] f1652_clk;
  logic [0:0] f1652_rst;
  logic [31:0] f1652_rdata;
  sr_buffer_32_1 f1652(.wen(f1652_wen), .wdata(f1652_wdata), .clk(f1652_clk), .rst(f1652_rst), .rdata(f1652_rdata));
  assign f1652_clk = clk;
  assign f1652_rst = rst;
  // Bindings to f1652

  // f1654
  logic [0:0] f1654_wen;
  logic [31:0] f1654_wdata;
  logic [0:0] f1654_clk;
  logic [0:0] f1654_rst;
  logic [31:0] f1654_rdata;
  sr_buffer_32_1 f1654(.wen(f1654_wen), .wdata(f1654_wdata), .clk(f1654_clk), .rst(f1654_rst), .rdata(f1654_rdata));
  assign f1654_clk = clk;
  assign f1654_rst = rst;
  // Bindings to f1654

  // f1656
  logic [0:0] f1656_wen;
  logic [31:0] f1656_wdata;
  logic [0:0] f1656_clk;
  logic [0:0] f1656_rst;
  logic [31:0] f1656_rdata;
  sr_buffer_32_1 f1656(.wen(f1656_wen), .wdata(f1656_wdata), .clk(f1656_clk), .rst(f1656_rst), .rdata(f1656_rdata));
  assign f1656_clk = clk;
  assign f1656_rst = rst;
  // Bindings to f1656

  // f1658
  logic [0:0] f1658_wen;
  logic [31:0] f1658_wdata;
  logic [0:0] f1658_clk;
  logic [0:0] f1658_rst;
  logic [31:0] f1658_rdata;
  sr_buffer_32_1 f1658(.wen(f1658_wen), .wdata(f1658_wdata), .clk(f1658_clk), .rst(f1658_rst), .rdata(f1658_rdata));
  assign f1658_clk = clk;
  assign f1658_rst = rst;
  // Bindings to f1658

  // f1660
  logic [0:0] f1660_wen;
  logic [31:0] f1660_wdata;
  logic [0:0] f1660_clk;
  logic [0:0] f1660_rst;
  logic [31:0] f1660_rdata;
  sr_buffer_32_1 f1660(.wen(f1660_wen), .wdata(f1660_wdata), .clk(f1660_clk), .rst(f1660_rst), .rdata(f1660_rdata));
  assign f1660_clk = clk;
  assign f1660_rst = rst;
  // Bindings to f1660

  // f1662
  logic [0:0] f1662_wen;
  logic [31:0] f1662_wdata;
  logic [0:0] f1662_clk;
  logic [0:0] f1662_rst;
  logic [31:0] f1662_rdata;
  sr_buffer_32_1 f1662(.wen(f1662_wen), .wdata(f1662_wdata), .clk(f1662_clk), .rst(f1662_rst), .rdata(f1662_rdata));
  assign f1662_clk = clk;
  assign f1662_rst = rst;
  // Bindings to f1662

  // f1664
  logic [0:0] f1664_wen;
  logic [31:0] f1664_wdata;
  logic [0:0] f1664_clk;
  logic [0:0] f1664_rst;
  logic [31:0] f1664_rdata;
  sr_buffer_32_1 f1664(.wen(f1664_wen), .wdata(f1664_wdata), .clk(f1664_clk), .rst(f1664_rst), .rdata(f1664_rdata));
  assign f1664_clk = clk;
  assign f1664_rst = rst;
  // Bindings to f1664

  // f1666
  logic [0:0] f1666_wen;
  logic [31:0] f1666_wdata;
  logic [0:0] f1666_clk;
  logic [0:0] f1666_rst;
  logic [31:0] f1666_rdata;
  sr_buffer_32_1 f1666(.wen(f1666_wen), .wdata(f1666_wdata), .clk(f1666_clk), .rst(f1666_rst), .rdata(f1666_rdata));
  assign f1666_clk = clk;
  assign f1666_rst = rst;
  // Bindings to f1666

  // f1668
  logic [0:0] f1668_wen;
  logic [31:0] f1668_wdata;
  logic [0:0] f1668_clk;
  logic [0:0] f1668_rst;
  logic [31:0] f1668_rdata;
  sr_buffer_32_1 f1668(.wen(f1668_wen), .wdata(f1668_wdata), .clk(f1668_clk), .rst(f1668_rst), .rdata(f1668_rdata));
  assign f1668_clk = clk;
  assign f1668_rst = rst;
  // Bindings to f1668

  // f1670
  logic [0:0] f1670_wen;
  logic [31:0] f1670_wdata;
  logic [0:0] f1670_clk;
  logic [0:0] f1670_rst;
  logic [31:0] f1670_rdata;
  sr_buffer_32_1 f1670(.wen(f1670_wen), .wdata(f1670_wdata), .clk(f1670_clk), .rst(f1670_rst), .rdata(f1670_rdata));
  assign f1670_clk = clk;
  assign f1670_rst = rst;
  // Bindings to f1670

  // f1672
  logic [0:0] f1672_wen;
  logic [31:0] f1672_wdata;
  logic [0:0] f1672_clk;
  logic [0:0] f1672_rst;
  logic [31:0] f1672_rdata;
  sr_buffer_32_1 f1672(.wen(f1672_wen), .wdata(f1672_wdata), .clk(f1672_clk), .rst(f1672_rst), .rdata(f1672_rdata));
  assign f1672_clk = clk;
  assign f1672_rst = rst;
  // Bindings to f1672

  // f1674
  logic [0:0] f1674_wen;
  logic [31:0] f1674_wdata;
  logic [0:0] f1674_clk;
  logic [0:0] f1674_rst;
  logic [31:0] f1674_rdata;
  sr_buffer_32_1 f1674(.wen(f1674_wen), .wdata(f1674_wdata), .clk(f1674_clk), .rst(f1674_rst), .rdata(f1674_rdata));
  assign f1674_clk = clk;
  assign f1674_rst = rst;
  // Bindings to f1674

  // f1676
  logic [0:0] f1676_wen;
  logic [31:0] f1676_wdata;
  logic [0:0] f1676_clk;
  logic [0:0] f1676_rst;
  logic [31:0] f1676_rdata;
  sr_buffer_32_1 f1676(.wen(f1676_wen), .wdata(f1676_wdata), .clk(f1676_clk), .rst(f1676_rst), .rdata(f1676_rdata));
  assign f1676_clk = clk;
  assign f1676_rst = rst;
  // Bindings to f1676

  // f1678
  logic [0:0] f1678_wen;
  logic [31:0] f1678_wdata;
  logic [0:0] f1678_clk;
  logic [0:0] f1678_rst;
  logic [31:0] f1678_rdata;
  sr_buffer_32_1 f1678(.wen(f1678_wen), .wdata(f1678_wdata), .clk(f1678_clk), .rst(f1678_rst), .rdata(f1678_rdata));
  assign f1678_clk = clk;
  assign f1678_rst = rst;
  // Bindings to f1678

  // f1680
  logic [0:0] f1680_wen;
  logic [31:0] f1680_wdata;
  logic [0:0] f1680_clk;
  logic [0:0] f1680_rst;
  logic [31:0] f1680_rdata;
  sr_buffer_32_1 f1680(.wen(f1680_wen), .wdata(f1680_wdata), .clk(f1680_clk), .rst(f1680_rst), .rdata(f1680_rdata));
  assign f1680_clk = clk;
  assign f1680_rst = rst;
  // Bindings to f1680

  // f1682
  logic [0:0] f1682_wen;
  logic [31:0] f1682_wdata;
  logic [0:0] f1682_clk;
  logic [0:0] f1682_rst;
  logic [31:0] f1682_rdata;
  sr_buffer_32_1 f1682(.wen(f1682_wen), .wdata(f1682_wdata), .clk(f1682_clk), .rst(f1682_rst), .rdata(f1682_rdata));
  assign f1682_clk = clk;
  assign f1682_rst = rst;
  // Bindings to f1682

  // f1684
  logic [0:0] f1684_wen;
  logic [31:0] f1684_wdata;
  logic [0:0] f1684_clk;
  logic [0:0] f1684_rst;
  logic [31:0] f1684_rdata;
  sr_buffer_32_1 f1684(.wen(f1684_wen), .wdata(f1684_wdata), .clk(f1684_clk), .rst(f1684_rst), .rdata(f1684_rdata));
  assign f1684_clk = clk;
  assign f1684_rst = rst;
  // Bindings to f1684

  // f1686
  logic [0:0] f1686_wen;
  logic [31:0] f1686_wdata;
  logic [0:0] f1686_clk;
  logic [0:0] f1686_rst;
  logic [31:0] f1686_rdata;
  sr_buffer_32_1 f1686(.wen(f1686_wen), .wdata(f1686_wdata), .clk(f1686_clk), .rst(f1686_rst), .rdata(f1686_rdata));
  assign f1686_clk = clk;
  assign f1686_rst = rst;
  // Bindings to f1686

  // f1688
  logic [0:0] f1688_wen;
  logic [31:0] f1688_wdata;
  logic [0:0] f1688_clk;
  logic [0:0] f1688_rst;
  logic [31:0] f1688_rdata;
  sr_buffer_32_1 f1688(.wen(f1688_wen), .wdata(f1688_wdata), .clk(f1688_clk), .rst(f1688_rst), .rdata(f1688_rdata));
  assign f1688_clk = clk;
  assign f1688_rst = rst;
  // Bindings to f1688

  // f1690
  logic [0:0] f1690_wen;
  logic [31:0] f1690_wdata;
  logic [0:0] f1690_clk;
  logic [0:0] f1690_rst;
  logic [31:0] f1690_rdata;
  sr_buffer_32_1 f1690(.wen(f1690_wen), .wdata(f1690_wdata), .clk(f1690_clk), .rst(f1690_rst), .rdata(f1690_rdata));
  assign f1690_clk = clk;
  assign f1690_rst = rst;
  // Bindings to f1690

  // f1692
  logic [0:0] f1692_wen;
  logic [31:0] f1692_wdata;
  logic [0:0] f1692_clk;
  logic [0:0] f1692_rst;
  logic [31:0] f1692_rdata;
  sr_buffer_32_1 f1692(.wen(f1692_wen), .wdata(f1692_wdata), .clk(f1692_clk), .rst(f1692_rst), .rdata(f1692_rdata));
  assign f1692_clk = clk;
  assign f1692_rst = rst;
  // Bindings to f1692

  // f1694
  logic [0:0] f1694_wen;
  logic [31:0] f1694_wdata;
  logic [0:0] f1694_clk;
  logic [0:0] f1694_rst;
  logic [31:0] f1694_rdata;
  sr_buffer_32_1 f1694(.wen(f1694_wen), .wdata(f1694_wdata), .clk(f1694_clk), .rst(f1694_rst), .rdata(f1694_rdata));
  assign f1694_clk = clk;
  assign f1694_rst = rst;
  // Bindings to f1694

  // f1696
  logic [0:0] f1696_wen;
  logic [31:0] f1696_wdata;
  logic [0:0] f1696_clk;
  logic [0:0] f1696_rst;
  logic [31:0] f1696_rdata;
  sr_buffer_32_1 f1696(.wen(f1696_wen), .wdata(f1696_wdata), .clk(f1696_clk), .rst(f1696_rst), .rdata(f1696_rdata));
  assign f1696_clk = clk;
  assign f1696_rst = rst;
  // Bindings to f1696

  // f1698
  logic [0:0] f1698_wen;
  logic [31:0] f1698_wdata;
  logic [0:0] f1698_clk;
  logic [0:0] f1698_rst;
  logic [31:0] f1698_rdata;
  sr_buffer_32_1 f1698(.wen(f1698_wen), .wdata(f1698_wdata), .clk(f1698_clk), .rst(f1698_rst), .rdata(f1698_rdata));
  assign f1698_clk = clk;
  assign f1698_rst = rst;
  // Bindings to f1698

  // f1700
  logic [0:0] f1700_wen;
  logic [31:0] f1700_wdata;
  logic [0:0] f1700_clk;
  logic [0:0] f1700_rst;
  logic [31:0] f1700_rdata;
  sr_buffer_32_1 f1700(.wen(f1700_wen), .wdata(f1700_wdata), .clk(f1700_clk), .rst(f1700_rst), .rdata(f1700_rdata));
  assign f1700_clk = clk;
  assign f1700_rst = rst;
  // Bindings to f1700

  // f1702
  logic [0:0] f1702_wen;
  logic [31:0] f1702_wdata;
  logic [0:0] f1702_clk;
  logic [0:0] f1702_rst;
  logic [31:0] f1702_rdata;
  sr_buffer_32_1 f1702(.wen(f1702_wen), .wdata(f1702_wdata), .clk(f1702_clk), .rst(f1702_rst), .rdata(f1702_rdata));
  assign f1702_clk = clk;
  assign f1702_rst = rst;
  // Bindings to f1702

  // f1704
  logic [0:0] f1704_wen;
  logic [31:0] f1704_wdata;
  logic [0:0] f1704_clk;
  logic [0:0] f1704_rst;
  logic [31:0] f1704_rdata;
  sr_buffer_32_1 f1704(.wen(f1704_wen), .wdata(f1704_wdata), .clk(f1704_clk), .rst(f1704_rst), .rdata(f1704_rdata));
  assign f1704_clk = clk;
  assign f1704_rst = rst;
  // Bindings to f1704

  // f1706
  logic [0:0] f1706_wen;
  logic [31:0] f1706_wdata;
  logic [0:0] f1706_clk;
  logic [0:0] f1706_rst;
  logic [31:0] f1706_rdata;
  sr_buffer_32_1 f1706(.wen(f1706_wen), .wdata(f1706_wdata), .clk(f1706_clk), .rst(f1706_rst), .rdata(f1706_rdata));
  assign f1706_clk = clk;
  assign f1706_rst = rst;
  // Bindings to f1706

  // f1708
  logic [0:0] f1708_wen;
  logic [31:0] f1708_wdata;
  logic [0:0] f1708_clk;
  logic [0:0] f1708_rst;
  logic [31:0] f1708_rdata;
  sr_buffer_32_1 f1708(.wen(f1708_wen), .wdata(f1708_wdata), .clk(f1708_clk), .rst(f1708_rst), .rdata(f1708_rdata));
  assign f1708_clk = clk;
  assign f1708_rst = rst;
  // Bindings to f1708

  // f1710
  logic [0:0] f1710_wen;
  logic [31:0] f1710_wdata;
  logic [0:0] f1710_clk;
  logic [0:0] f1710_rst;
  logic [31:0] f1710_rdata;
  sr_buffer_32_1 f1710(.wen(f1710_wen), .wdata(f1710_wdata), .clk(f1710_clk), .rst(f1710_rst), .rdata(f1710_rdata));
  assign f1710_clk = clk;
  assign f1710_rst = rst;
  // Bindings to f1710

  // f1712
  logic [0:0] f1712_wen;
  logic [31:0] f1712_wdata;
  logic [0:0] f1712_clk;
  logic [0:0] f1712_rst;
  logic [31:0] f1712_rdata;
  sr_buffer_32_1 f1712(.wen(f1712_wen), .wdata(f1712_wdata), .clk(f1712_clk), .rst(f1712_rst), .rdata(f1712_rdata));
  assign f1712_clk = clk;
  assign f1712_rst = rst;
  // Bindings to f1712

  // f1714
  logic [0:0] f1714_wen;
  logic [31:0] f1714_wdata;
  logic [0:0] f1714_clk;
  logic [0:0] f1714_rst;
  logic [31:0] f1714_rdata;
  sr_buffer_32_1 f1714(.wen(f1714_wen), .wdata(f1714_wdata), .clk(f1714_clk), .rst(f1714_rst), .rdata(f1714_rdata));
  assign f1714_clk = clk;
  assign f1714_rst = rst;
  // Bindings to f1714

  // f1716
  logic [0:0] f1716_wen;
  logic [31:0] f1716_wdata;
  logic [0:0] f1716_clk;
  logic [0:0] f1716_rst;
  logic [31:0] f1716_rdata;
  sr_buffer_32_1 f1716(.wen(f1716_wen), .wdata(f1716_wdata), .clk(f1716_clk), .rst(f1716_rst), .rdata(f1716_rdata));
  assign f1716_clk = clk;
  assign f1716_rst = rst;
  // Bindings to f1716

  // f1718
  logic [0:0] f1718_wen;
  logic [31:0] f1718_wdata;
  logic [0:0] f1718_clk;
  logic [0:0] f1718_rst;
  logic [31:0] f1718_rdata;
  sr_buffer_32_1 f1718(.wen(f1718_wen), .wdata(f1718_wdata), .clk(f1718_clk), .rst(f1718_rst), .rdata(f1718_rdata));
  assign f1718_clk = clk;
  assign f1718_rst = rst;
  // Bindings to f1718

  // f1720
  logic [0:0] f1720_wen;
  logic [31:0] f1720_wdata;
  logic [0:0] f1720_clk;
  logic [0:0] f1720_rst;
  logic [31:0] f1720_rdata;
  sr_buffer_32_1 f1720(.wen(f1720_wen), .wdata(f1720_wdata), .clk(f1720_clk), .rst(f1720_rst), .rdata(f1720_rdata));
  assign f1720_clk = clk;
  assign f1720_rst = rst;
  // Bindings to f1720

  // f1722
  logic [0:0] f1722_wen;
  logic [31:0] f1722_wdata;
  logic [0:0] f1722_clk;
  logic [0:0] f1722_rst;
  logic [31:0] f1722_rdata;
  sr_buffer_32_1 f1722(.wen(f1722_wen), .wdata(f1722_wdata), .clk(f1722_clk), .rst(f1722_rst), .rdata(f1722_rdata));
  assign f1722_clk = clk;
  assign f1722_rst = rst;
  // Bindings to f1722

  // f1724
  logic [0:0] f1724_wen;
  logic [31:0] f1724_wdata;
  logic [0:0] f1724_clk;
  logic [0:0] f1724_rst;
  logic [31:0] f1724_rdata;
  sr_buffer_32_1 f1724(.wen(f1724_wen), .wdata(f1724_wdata), .clk(f1724_clk), .rst(f1724_rst), .rdata(f1724_rdata));
  assign f1724_clk = clk;
  assign f1724_rst = rst;
  // Bindings to f1724

  // f1726
  logic [0:0] f1726_wen;
  logic [31:0] f1726_wdata;
  logic [0:0] f1726_clk;
  logic [0:0] f1726_rst;
  logic [31:0] f1726_rdata;
  sr_buffer_32_1 f1726(.wen(f1726_wen), .wdata(f1726_wdata), .clk(f1726_clk), .rst(f1726_rst), .rdata(f1726_rdata));
  assign f1726_clk = clk;
  assign f1726_rst = rst;
  // Bindings to f1726

  // f1728
  logic [0:0] f1728_wen;
  logic [31:0] f1728_wdata;
  logic [0:0] f1728_clk;
  logic [0:0] f1728_rst;
  logic [31:0] f1728_rdata;
  sr_buffer_32_1 f1728(.wen(f1728_wen), .wdata(f1728_wdata), .clk(f1728_clk), .rst(f1728_rst), .rdata(f1728_rdata));
  assign f1728_clk = clk;
  assign f1728_rst = rst;
  // Bindings to f1728

  // f1730
  logic [0:0] f1730_wen;
  logic [31:0] f1730_wdata;
  logic [0:0] f1730_clk;
  logic [0:0] f1730_rst;
  logic [31:0] f1730_rdata;
  sr_buffer_32_1 f1730(.wen(f1730_wen), .wdata(f1730_wdata), .clk(f1730_clk), .rst(f1730_rst), .rdata(f1730_rdata));
  assign f1730_clk = clk;
  assign f1730_rst = rst;
  // Bindings to f1730

  // f1732
  logic [0:0] f1732_wen;
  logic [31:0] f1732_wdata;
  logic [0:0] f1732_clk;
  logic [0:0] f1732_rst;
  logic [31:0] f1732_rdata;
  sr_buffer_32_1 f1732(.wen(f1732_wen), .wdata(f1732_wdata), .clk(f1732_clk), .rst(f1732_rst), .rdata(f1732_rdata));
  assign f1732_clk = clk;
  assign f1732_rst = rst;
  // Bindings to f1732

  // f1734
  logic [0:0] f1734_wen;
  logic [31:0] f1734_wdata;
  logic [0:0] f1734_clk;
  logic [0:0] f1734_rst;
  logic [31:0] f1734_rdata;
  sr_buffer_32_1 f1734(.wen(f1734_wen), .wdata(f1734_wdata), .clk(f1734_clk), .rst(f1734_rst), .rdata(f1734_rdata));
  assign f1734_clk = clk;
  assign f1734_rst = rst;
  // Bindings to f1734

  // f1736
  logic [0:0] f1736_wen;
  logic [31:0] f1736_wdata;
  logic [0:0] f1736_clk;
  logic [0:0] f1736_rst;
  logic [31:0] f1736_rdata;
  sr_buffer_32_1 f1736(.wen(f1736_wen), .wdata(f1736_wdata), .clk(f1736_clk), .rst(f1736_rst), .rdata(f1736_rdata));
  assign f1736_clk = clk;
  assign f1736_rst = rst;
  // Bindings to f1736

  // f1738
  logic [0:0] f1738_wen;
  logic [31:0] f1738_wdata;
  logic [0:0] f1738_clk;
  logic [0:0] f1738_rst;
  logic [31:0] f1738_rdata;
  sr_buffer_32_1 f1738(.wen(f1738_wen), .wdata(f1738_wdata), .clk(f1738_clk), .rst(f1738_rst), .rdata(f1738_rdata));
  assign f1738_clk = clk;
  assign f1738_rst = rst;
  // Bindings to f1738

  // f1740
  logic [0:0] f1740_wen;
  logic [31:0] f1740_wdata;
  logic [0:0] f1740_clk;
  logic [0:0] f1740_rst;
  logic [31:0] f1740_rdata;
  sr_buffer_32_1 f1740(.wen(f1740_wen), .wdata(f1740_wdata), .clk(f1740_clk), .rst(f1740_rst), .rdata(f1740_rdata));
  assign f1740_clk = clk;
  assign f1740_rst = rst;
  // Bindings to f1740

  // f1742
  logic [0:0] f1742_wen;
  logic [31:0] f1742_wdata;
  logic [0:0] f1742_clk;
  logic [0:0] f1742_rst;
  logic [31:0] f1742_rdata;
  sr_buffer_32_1 f1742(.wen(f1742_wen), .wdata(f1742_wdata), .clk(f1742_clk), .rst(f1742_rst), .rdata(f1742_rdata));
  assign f1742_clk = clk;
  assign f1742_rst = rst;
  // Bindings to f1742

  // f1744
  logic [0:0] f1744_wen;
  logic [31:0] f1744_wdata;
  logic [0:0] f1744_clk;
  logic [0:0] f1744_rst;
  logic [31:0] f1744_rdata;
  sr_buffer_32_1 f1744(.wen(f1744_wen), .wdata(f1744_wdata), .clk(f1744_clk), .rst(f1744_rst), .rdata(f1744_rdata));
  assign f1744_clk = clk;
  assign f1744_rst = rst;
  // Bindings to f1744

  // f1746
  logic [0:0] f1746_wen;
  logic [31:0] f1746_wdata;
  logic [0:0] f1746_clk;
  logic [0:0] f1746_rst;
  logic [31:0] f1746_rdata;
  sr_buffer_32_1 f1746(.wen(f1746_wen), .wdata(f1746_wdata), .clk(f1746_clk), .rst(f1746_rst), .rdata(f1746_rdata));
  assign f1746_clk = clk;
  assign f1746_rst = rst;
  // Bindings to f1746

  // f1748
  logic [0:0] f1748_wen;
  logic [31:0] f1748_wdata;
  logic [0:0] f1748_clk;
  logic [0:0] f1748_rst;
  logic [31:0] f1748_rdata;
  sr_buffer_32_1 f1748(.wen(f1748_wen), .wdata(f1748_wdata), .clk(f1748_clk), .rst(f1748_rst), .rdata(f1748_rdata));
  assign f1748_clk = clk;
  assign f1748_rst = rst;
  // Bindings to f1748

  // f1750
  logic [0:0] f1750_wen;
  logic [31:0] f1750_wdata;
  logic [0:0] f1750_clk;
  logic [0:0] f1750_rst;
  logic [31:0] f1750_rdata;
  sr_buffer_32_1 f1750(.wen(f1750_wen), .wdata(f1750_wdata), .clk(f1750_clk), .rst(f1750_rst), .rdata(f1750_rdata));
  assign f1750_clk = clk;
  assign f1750_rst = rst;
  // Bindings to f1750

  // f1752
  logic [0:0] f1752_wen;
  logic [31:0] f1752_wdata;
  logic [0:0] f1752_clk;
  logic [0:0] f1752_rst;
  logic [31:0] f1752_rdata;
  sr_buffer_32_1 f1752(.wen(f1752_wen), .wdata(f1752_wdata), .clk(f1752_clk), .rst(f1752_rst), .rdata(f1752_rdata));
  assign f1752_clk = clk;
  assign f1752_rst = rst;
  // Bindings to f1752

  // f1754
  logic [0:0] f1754_wen;
  logic [31:0] f1754_wdata;
  logic [0:0] f1754_clk;
  logic [0:0] f1754_rst;
  logic [31:0] f1754_rdata;
  sr_buffer_32_1 f1754(.wen(f1754_wen), .wdata(f1754_wdata), .clk(f1754_clk), .rst(f1754_rst), .rdata(f1754_rdata));
  assign f1754_clk = clk;
  assign f1754_rst = rst;
  // Bindings to f1754

  // f1756
  logic [0:0] f1756_wen;
  logic [31:0] f1756_wdata;
  logic [0:0] f1756_clk;
  logic [0:0] f1756_rst;
  logic [31:0] f1756_rdata;
  sr_buffer_32_1 f1756(.wen(f1756_wen), .wdata(f1756_wdata), .clk(f1756_clk), .rst(f1756_rst), .rdata(f1756_rdata));
  assign f1756_clk = clk;
  assign f1756_rst = rst;
  // Bindings to f1756

  // f1758
  logic [0:0] f1758_wen;
  logic [31:0] f1758_wdata;
  logic [0:0] f1758_clk;
  logic [0:0] f1758_rst;
  logic [31:0] f1758_rdata;
  sr_buffer_32_1 f1758(.wen(f1758_wen), .wdata(f1758_wdata), .clk(f1758_clk), .rst(f1758_rst), .rdata(f1758_rdata));
  assign f1758_clk = clk;
  assign f1758_rst = rst;
  // Bindings to f1758

  // f1760
  logic [0:0] f1760_wen;
  logic [31:0] f1760_wdata;
  logic [0:0] f1760_clk;
  logic [0:0] f1760_rst;
  logic [31:0] f1760_rdata;
  sr_buffer_32_1 f1760(.wen(f1760_wen), .wdata(f1760_wdata), .clk(f1760_clk), .rst(f1760_rst), .rdata(f1760_rdata));
  assign f1760_clk = clk;
  assign f1760_rst = rst;
  // Bindings to f1760

  // f1762
  logic [0:0] f1762_wen;
  logic [31:0] f1762_wdata;
  logic [0:0] f1762_clk;
  logic [0:0] f1762_rst;
  logic [31:0] f1762_rdata;
  sr_buffer_32_1 f1762(.wen(f1762_wen), .wdata(f1762_wdata), .clk(f1762_clk), .rst(f1762_rst), .rdata(f1762_rdata));
  assign f1762_clk = clk;
  assign f1762_rst = rst;
  // Bindings to f1762

  // f1764
  logic [0:0] f1764_wen;
  logic [31:0] f1764_wdata;
  logic [0:0] f1764_clk;
  logic [0:0] f1764_rst;
  logic [31:0] f1764_rdata;
  sr_buffer_32_1 f1764(.wen(f1764_wen), .wdata(f1764_wdata), .clk(f1764_clk), .rst(f1764_rst), .rdata(f1764_rdata));
  assign f1764_clk = clk;
  assign f1764_rst = rst;
  // Bindings to f1764

  // f1766
  logic [0:0] f1766_wen;
  logic [31:0] f1766_wdata;
  logic [0:0] f1766_clk;
  logic [0:0] f1766_rst;
  logic [31:0] f1766_rdata;
  sr_buffer_32_1 f1766(.wen(f1766_wen), .wdata(f1766_wdata), .clk(f1766_clk), .rst(f1766_rst), .rdata(f1766_rdata));
  assign f1766_clk = clk;
  assign f1766_rst = rst;
  // Bindings to f1766

  // f1768
  logic [0:0] f1768_wen;
  logic [31:0] f1768_wdata;
  logic [0:0] f1768_clk;
  logic [0:0] f1768_rst;
  logic [31:0] f1768_rdata;
  sr_buffer_32_1 f1768(.wen(f1768_wen), .wdata(f1768_wdata), .clk(f1768_clk), .rst(f1768_rst), .rdata(f1768_rdata));
  assign f1768_clk = clk;
  assign f1768_rst = rst;
  // Bindings to f1768

  // f1770
  logic [0:0] f1770_wen;
  logic [31:0] f1770_wdata;
  logic [0:0] f1770_clk;
  logic [0:0] f1770_rst;
  logic [31:0] f1770_rdata;
  sr_buffer_32_1 f1770(.wen(f1770_wen), .wdata(f1770_wdata), .clk(f1770_clk), .rst(f1770_rst), .rdata(f1770_rdata));
  assign f1770_clk = clk;
  assign f1770_rst = rst;
  // Bindings to f1770

  // f1772
  logic [0:0] f1772_wen;
  logic [31:0] f1772_wdata;
  logic [0:0] f1772_clk;
  logic [0:0] f1772_rst;
  logic [31:0] f1772_rdata;
  sr_buffer_32_1 f1772(.wen(f1772_wen), .wdata(f1772_wdata), .clk(f1772_clk), .rst(f1772_rst), .rdata(f1772_rdata));
  assign f1772_clk = clk;
  assign f1772_rst = rst;
  // Bindings to f1772

  // f1774
  logic [0:0] f1774_wen;
  logic [31:0] f1774_wdata;
  logic [0:0] f1774_clk;
  logic [0:0] f1774_rst;
  logic [31:0] f1774_rdata;
  sr_buffer_32_1 f1774(.wen(f1774_wen), .wdata(f1774_wdata), .clk(f1774_clk), .rst(f1774_rst), .rdata(f1774_rdata));
  assign f1774_clk = clk;
  assign f1774_rst = rst;
  // Bindings to f1774

  // f1776
  logic [0:0] f1776_wen;
  logic [31:0] f1776_wdata;
  logic [0:0] f1776_clk;
  logic [0:0] f1776_rst;
  logic [31:0] f1776_rdata;
  sr_buffer_32_1 f1776(.wen(f1776_wen), .wdata(f1776_wdata), .clk(f1776_clk), .rst(f1776_rst), .rdata(f1776_rdata));
  assign f1776_clk = clk;
  assign f1776_rst = rst;
  // Bindings to f1776

  // f1778
  logic [0:0] f1778_wen;
  logic [31:0] f1778_wdata;
  logic [0:0] f1778_clk;
  logic [0:0] f1778_rst;
  logic [31:0] f1778_rdata;
  sr_buffer_32_1 f1778(.wen(f1778_wen), .wdata(f1778_wdata), .clk(f1778_clk), .rst(f1778_rst), .rdata(f1778_rdata));
  assign f1778_clk = clk;
  assign f1778_rst = rst;
  // Bindings to f1778

  // f1780
  logic [0:0] f1780_wen;
  logic [31:0] f1780_wdata;
  logic [0:0] f1780_clk;
  logic [0:0] f1780_rst;
  logic [31:0] f1780_rdata;
  sr_buffer_32_1 f1780(.wen(f1780_wen), .wdata(f1780_wdata), .clk(f1780_clk), .rst(f1780_rst), .rdata(f1780_rdata));
  assign f1780_clk = clk;
  assign f1780_rst = rst;
  // Bindings to f1780

  // f1782
  logic [0:0] f1782_wen;
  logic [31:0] f1782_wdata;
  logic [0:0] f1782_clk;
  logic [0:0] f1782_rst;
  logic [31:0] f1782_rdata;
  sr_buffer_32_1 f1782(.wen(f1782_wen), .wdata(f1782_wdata), .clk(f1782_clk), .rst(f1782_rst), .rdata(f1782_rdata));
  assign f1782_clk = clk;
  assign f1782_rst = rst;
  // Bindings to f1782

  // f1784
  logic [0:0] f1784_wen;
  logic [31:0] f1784_wdata;
  logic [0:0] f1784_clk;
  logic [0:0] f1784_rst;
  logic [31:0] f1784_rdata;
  sr_buffer_32_1 f1784(.wen(f1784_wen), .wdata(f1784_wdata), .clk(f1784_clk), .rst(f1784_rst), .rdata(f1784_rdata));
  assign f1784_clk = clk;
  assign f1784_rst = rst;
  // Bindings to f1784

  // f1786
  logic [0:0] f1786_wen;
  logic [31:0] f1786_wdata;
  logic [0:0] f1786_clk;
  logic [0:0] f1786_rst;
  logic [31:0] f1786_rdata;
  sr_buffer_32_1 f1786(.wen(f1786_wen), .wdata(f1786_wdata), .clk(f1786_clk), .rst(f1786_rst), .rdata(f1786_rdata));
  assign f1786_clk = clk;
  assign f1786_rst = rst;
  // Bindings to f1786

  // f1788
  logic [0:0] f1788_wen;
  logic [31:0] f1788_wdata;
  logic [0:0] f1788_clk;
  logic [0:0] f1788_rst;
  logic [31:0] f1788_rdata;
  sr_buffer_32_1 f1788(.wen(f1788_wen), .wdata(f1788_wdata), .clk(f1788_clk), .rst(f1788_rst), .rdata(f1788_rdata));
  assign f1788_clk = clk;
  assign f1788_rst = rst;
  // Bindings to f1788

  // f1790
  logic [0:0] f1790_wen;
  logic [31:0] f1790_wdata;
  logic [0:0] f1790_clk;
  logic [0:0] f1790_rst;
  logic [31:0] f1790_rdata;
  sr_buffer_32_1 f1790(.wen(f1790_wen), .wdata(f1790_wdata), .clk(f1790_clk), .rst(f1790_rst), .rdata(f1790_rdata));
  assign f1790_clk = clk;
  assign f1790_rst = rst;
  // Bindings to f1790

  // f1792
  logic [0:0] f1792_wen;
  logic [31:0] f1792_wdata;
  logic [0:0] f1792_clk;
  logic [0:0] f1792_rst;
  logic [31:0] f1792_rdata;
  sr_buffer_32_1 f1792(.wen(f1792_wen), .wdata(f1792_wdata), .clk(f1792_clk), .rst(f1792_rst), .rdata(f1792_rdata));
  assign f1792_clk = clk;
  assign f1792_rst = rst;
  // Bindings to f1792

  // f1794
  logic [0:0] f1794_wen;
  logic [31:0] f1794_wdata;
  logic [0:0] f1794_clk;
  logic [0:0] f1794_rst;
  logic [31:0] f1794_rdata;
  sr_buffer_32_1 f1794(.wen(f1794_wen), .wdata(f1794_wdata), .clk(f1794_clk), .rst(f1794_rst), .rdata(f1794_rdata));
  assign f1794_clk = clk;
  assign f1794_rst = rst;
  // Bindings to f1794

  // f1796
  logic [0:0] f1796_wen;
  logic [31:0] f1796_wdata;
  logic [0:0] f1796_clk;
  logic [0:0] f1796_rst;
  logic [31:0] f1796_rdata;
  sr_buffer_32_1 f1796(.wen(f1796_wen), .wdata(f1796_wdata), .clk(f1796_clk), .rst(f1796_rst), .rdata(f1796_rdata));
  assign f1796_clk = clk;
  assign f1796_rst = rst;
  // Bindings to f1796

  // f1798
  logic [0:0] f1798_wen;
  logic [31:0] f1798_wdata;
  logic [0:0] f1798_clk;
  logic [0:0] f1798_rst;
  logic [31:0] f1798_rdata;
  sr_buffer_32_1 f1798(.wen(f1798_wen), .wdata(f1798_wdata), .clk(f1798_clk), .rst(f1798_rst), .rdata(f1798_rdata));
  assign f1798_clk = clk;
  assign f1798_rst = rst;
  // Bindings to f1798

  // f1800
  logic [0:0] f1800_wen;
  logic [31:0] f1800_wdata;
  logic [0:0] f1800_clk;
  logic [0:0] f1800_rst;
  logic [31:0] f1800_rdata;
  sr_buffer_32_1 f1800(.wen(f1800_wen), .wdata(f1800_wdata), .clk(f1800_clk), .rst(f1800_rst), .rdata(f1800_rdata));
  assign f1800_clk = clk;
  assign f1800_rst = rst;
  // Bindings to f1800

  // f1802
  logic [0:0] f1802_wen;
  logic [31:0] f1802_wdata;
  logic [0:0] f1802_clk;
  logic [0:0] f1802_rst;
  logic [31:0] f1802_rdata;
  sr_buffer_32_1 f1802(.wen(f1802_wen), .wdata(f1802_wdata), .clk(f1802_clk), .rst(f1802_rst), .rdata(f1802_rdata));
  assign f1802_clk = clk;
  assign f1802_rst = rst;
  // Bindings to f1802

  // f1804
  logic [0:0] f1804_wen;
  logic [31:0] f1804_wdata;
  logic [0:0] f1804_clk;
  logic [0:0] f1804_rst;
  logic [31:0] f1804_rdata;
  sr_buffer_32_1 f1804(.wen(f1804_wen), .wdata(f1804_wdata), .clk(f1804_clk), .rst(f1804_rst), .rdata(f1804_rdata));
  assign f1804_clk = clk;
  assign f1804_rst = rst;
  // Bindings to f1804

  // f1806
  logic [0:0] f1806_wen;
  logic [31:0] f1806_wdata;
  logic [0:0] f1806_clk;
  logic [0:0] f1806_rst;
  logic [31:0] f1806_rdata;
  sr_buffer_32_1 f1806(.wen(f1806_wen), .wdata(f1806_wdata), .clk(f1806_clk), .rst(f1806_rst), .rdata(f1806_rdata));
  assign f1806_clk = clk;
  assign f1806_rst = rst;
  // Bindings to f1806

  // f1808
  logic [0:0] f1808_wen;
  logic [31:0] f1808_wdata;
  logic [0:0] f1808_clk;
  logic [0:0] f1808_rst;
  logic [31:0] f1808_rdata;
  sr_buffer_32_1 f1808(.wen(f1808_wen), .wdata(f1808_wdata), .clk(f1808_clk), .rst(f1808_rst), .rdata(f1808_rdata));
  assign f1808_clk = clk;
  assign f1808_rst = rst;
  // Bindings to f1808

  // f1810
  logic [0:0] f1810_wen;
  logic [31:0] f1810_wdata;
  logic [0:0] f1810_clk;
  logic [0:0] f1810_rst;
  logic [31:0] f1810_rdata;
  sr_buffer_32_1 f1810(.wen(f1810_wen), .wdata(f1810_wdata), .clk(f1810_clk), .rst(f1810_rst), .rdata(f1810_rdata));
  assign f1810_clk = clk;
  assign f1810_rst = rst;
  // Bindings to f1810

  // f1812
  logic [0:0] f1812_wen;
  logic [31:0] f1812_wdata;
  logic [0:0] f1812_clk;
  logic [0:0] f1812_rst;
  logic [31:0] f1812_rdata;
  sr_buffer_32_1 f1812(.wen(f1812_wen), .wdata(f1812_wdata), .clk(f1812_clk), .rst(f1812_rst), .rdata(f1812_rdata));
  assign f1812_clk = clk;
  assign f1812_rst = rst;
  // Bindings to f1812

  // f1814
  logic [0:0] f1814_wen;
  logic [31:0] f1814_wdata;
  logic [0:0] f1814_clk;
  logic [0:0] f1814_rst;
  logic [31:0] f1814_rdata;
  sr_buffer_32_1 f1814(.wen(f1814_wen), .wdata(f1814_wdata), .clk(f1814_clk), .rst(f1814_rst), .rdata(f1814_rdata));
  assign f1814_clk = clk;
  assign f1814_rst = rst;
  // Bindings to f1814

  // f1816
  logic [0:0] f1816_wen;
  logic [31:0] f1816_wdata;
  logic [0:0] f1816_clk;
  logic [0:0] f1816_rst;
  logic [31:0] f1816_rdata;
  sr_buffer_32_1 f1816(.wen(f1816_wen), .wdata(f1816_wdata), .clk(f1816_clk), .rst(f1816_rst), .rdata(f1816_rdata));
  assign f1816_clk = clk;
  assign f1816_rst = rst;
  // Bindings to f1816

  // f1818
  logic [0:0] f1818_wen;
  logic [31:0] f1818_wdata;
  logic [0:0] f1818_clk;
  logic [0:0] f1818_rst;
  logic [31:0] f1818_rdata;
  sr_buffer_32_1 f1818(.wen(f1818_wen), .wdata(f1818_wdata), .clk(f1818_clk), .rst(f1818_rst), .rdata(f1818_rdata));
  assign f1818_clk = clk;
  assign f1818_rst = rst;
  // Bindings to f1818

  // f1820
  logic [0:0] f1820_wen;
  logic [31:0] f1820_wdata;
  logic [0:0] f1820_clk;
  logic [0:0] f1820_rst;
  logic [31:0] f1820_rdata;
  sr_buffer_32_1 f1820(.wen(f1820_wen), .wdata(f1820_wdata), .clk(f1820_clk), .rst(f1820_rst), .rdata(f1820_rdata));
  assign f1820_clk = clk;
  assign f1820_rst = rst;
  // Bindings to f1820

  // f1822
  logic [0:0] f1822_wen;
  logic [31:0] f1822_wdata;
  logic [0:0] f1822_clk;
  logic [0:0] f1822_rst;
  logic [31:0] f1822_rdata;
  sr_buffer_32_1 f1822(.wen(f1822_wen), .wdata(f1822_wdata), .clk(f1822_clk), .rst(f1822_rst), .rdata(f1822_rdata));
  assign f1822_clk = clk;
  assign f1822_rst = rst;
  // Bindings to f1822

  // f1824
  logic [0:0] f1824_wen;
  logic [31:0] f1824_wdata;
  logic [0:0] f1824_clk;
  logic [0:0] f1824_rst;
  logic [31:0] f1824_rdata;
  sr_buffer_32_1 f1824(.wen(f1824_wen), .wdata(f1824_wdata), .clk(f1824_clk), .rst(f1824_rst), .rdata(f1824_rdata));
  assign f1824_clk = clk;
  assign f1824_rst = rst;
  // Bindings to f1824

  // f1826
  logic [0:0] f1826_wen;
  logic [31:0] f1826_wdata;
  logic [0:0] f1826_clk;
  logic [0:0] f1826_rst;
  logic [31:0] f1826_rdata;
  sr_buffer_32_1 f1826(.wen(f1826_wen), .wdata(f1826_wdata), .clk(f1826_clk), .rst(f1826_rst), .rdata(f1826_rdata));
  assign f1826_clk = clk;
  assign f1826_rst = rst;
  // Bindings to f1826

  // f1828
  logic [0:0] f1828_wen;
  logic [31:0] f1828_wdata;
  logic [0:0] f1828_clk;
  logic [0:0] f1828_rst;
  logic [31:0] f1828_rdata;
  sr_buffer_32_1 f1828(.wen(f1828_wen), .wdata(f1828_wdata), .clk(f1828_clk), .rst(f1828_rst), .rdata(f1828_rdata));
  assign f1828_clk = clk;
  assign f1828_rst = rst;
  // Bindings to f1828

  // f1830
  logic [0:0] f1830_wen;
  logic [31:0] f1830_wdata;
  logic [0:0] f1830_clk;
  logic [0:0] f1830_rst;
  logic [31:0] f1830_rdata;
  sr_buffer_32_1 f1830(.wen(f1830_wen), .wdata(f1830_wdata), .clk(f1830_clk), .rst(f1830_rst), .rdata(f1830_rdata));
  assign f1830_clk = clk;
  assign f1830_rst = rst;
  // Bindings to f1830

  // f1832
  logic [0:0] f1832_wen;
  logic [31:0] f1832_wdata;
  logic [0:0] f1832_clk;
  logic [0:0] f1832_rst;
  logic [31:0] f1832_rdata;
  sr_buffer_32_1 f1832(.wen(f1832_wen), .wdata(f1832_wdata), .clk(f1832_clk), .rst(f1832_rst), .rdata(f1832_rdata));
  assign f1832_clk = clk;
  assign f1832_rst = rst;
  // Bindings to f1832

  // f1834
  logic [0:0] f1834_wen;
  logic [31:0] f1834_wdata;
  logic [0:0] f1834_clk;
  logic [0:0] f1834_rst;
  logic [31:0] f1834_rdata;
  sr_buffer_32_1 f1834(.wen(f1834_wen), .wdata(f1834_wdata), .clk(f1834_clk), .rst(f1834_rst), .rdata(f1834_rdata));
  assign f1834_clk = clk;
  assign f1834_rst = rst;
  // Bindings to f1834

  // f1836
  logic [0:0] f1836_wen;
  logic [31:0] f1836_wdata;
  logic [0:0] f1836_clk;
  logic [0:0] f1836_rst;
  logic [31:0] f1836_rdata;
  sr_buffer_32_1 f1836(.wen(f1836_wen), .wdata(f1836_wdata), .clk(f1836_clk), .rst(f1836_rst), .rdata(f1836_rdata));
  assign f1836_clk = clk;
  assign f1836_rst = rst;
  // Bindings to f1836

  // f1838
  logic [0:0] f1838_wen;
  logic [31:0] f1838_wdata;
  logic [0:0] f1838_clk;
  logic [0:0] f1838_rst;
  logic [31:0] f1838_rdata;
  sr_buffer_32_1 f1838(.wen(f1838_wen), .wdata(f1838_wdata), .clk(f1838_clk), .rst(f1838_rst), .rdata(f1838_rdata));
  assign f1838_clk = clk;
  assign f1838_rst = rst;
  // Bindings to f1838

  // f1840
  logic [0:0] f1840_wen;
  logic [31:0] f1840_wdata;
  logic [0:0] f1840_clk;
  logic [0:0] f1840_rst;
  logic [31:0] f1840_rdata;
  sr_buffer_32_1 f1840(.wen(f1840_wen), .wdata(f1840_wdata), .clk(f1840_clk), .rst(f1840_rst), .rdata(f1840_rdata));
  assign f1840_clk = clk;
  assign f1840_rst = rst;
  // Bindings to f1840

  // f1842
  logic [0:0] f1842_wen;
  logic [31:0] f1842_wdata;
  logic [0:0] f1842_clk;
  logic [0:0] f1842_rst;
  logic [31:0] f1842_rdata;
  sr_buffer_32_1 f1842(.wen(f1842_wen), .wdata(f1842_wdata), .clk(f1842_clk), .rst(f1842_rst), .rdata(f1842_rdata));
  assign f1842_clk = clk;
  assign f1842_rst = rst;
  // Bindings to f1842

  // f1844
  logic [0:0] f1844_wen;
  logic [31:0] f1844_wdata;
  logic [0:0] f1844_clk;
  logic [0:0] f1844_rst;
  logic [31:0] f1844_rdata;
  sr_buffer_32_1 f1844(.wen(f1844_wen), .wdata(f1844_wdata), .clk(f1844_clk), .rst(f1844_rst), .rdata(f1844_rdata));
  assign f1844_clk = clk;
  assign f1844_rst = rst;
  // Bindings to f1844

  // f1846
  logic [0:0] f1846_wen;
  logic [31:0] f1846_wdata;
  logic [0:0] f1846_clk;
  logic [0:0] f1846_rst;
  logic [31:0] f1846_rdata;
  sr_buffer_32_1 f1846(.wen(f1846_wen), .wdata(f1846_wdata), .clk(f1846_clk), .rst(f1846_rst), .rdata(f1846_rdata));
  assign f1846_clk = clk;
  assign f1846_rst = rst;
  // Bindings to f1846

  // f1848
  logic [0:0] f1848_wen;
  logic [31:0] f1848_wdata;
  logic [0:0] f1848_clk;
  logic [0:0] f1848_rst;
  logic [31:0] f1848_rdata;
  sr_buffer_32_1 f1848(.wen(f1848_wen), .wdata(f1848_wdata), .clk(f1848_clk), .rst(f1848_rst), .rdata(f1848_rdata));
  assign f1848_clk = clk;
  assign f1848_rst = rst;
  // Bindings to f1848

  // f1850
  logic [0:0] f1850_wen;
  logic [31:0] f1850_wdata;
  logic [0:0] f1850_clk;
  logic [0:0] f1850_rst;
  logic [31:0] f1850_rdata;
  sr_buffer_32_1 f1850(.wen(f1850_wen), .wdata(f1850_wdata), .clk(f1850_clk), .rst(f1850_rst), .rdata(f1850_rdata));
  assign f1850_clk = clk;
  assign f1850_rst = rst;
  // Bindings to f1850

  // f1852
  logic [0:0] f1852_wen;
  logic [31:0] f1852_wdata;
  logic [0:0] f1852_clk;
  logic [0:0] f1852_rst;
  logic [31:0] f1852_rdata;
  sr_buffer_32_1 f1852(.wen(f1852_wen), .wdata(f1852_wdata), .clk(f1852_clk), .rst(f1852_rst), .rdata(f1852_rdata));
  assign f1852_clk = clk;
  assign f1852_rst = rst;
  // Bindings to f1852

  // f1854
  logic [0:0] f1854_wen;
  logic [31:0] f1854_wdata;
  logic [0:0] f1854_clk;
  logic [0:0] f1854_rst;
  logic [31:0] f1854_rdata;
  sr_buffer_32_1 f1854(.wen(f1854_wen), .wdata(f1854_wdata), .clk(f1854_clk), .rst(f1854_rst), .rdata(f1854_rdata));
  assign f1854_clk = clk;
  assign f1854_rst = rst;
  // Bindings to f1854

  // f1856
  logic [0:0] f1856_wen;
  logic [31:0] f1856_wdata;
  logic [0:0] f1856_clk;
  logic [0:0] f1856_rst;
  logic [31:0] f1856_rdata;
  sr_buffer_32_1 f1856(.wen(f1856_wen), .wdata(f1856_wdata), .clk(f1856_clk), .rst(f1856_rst), .rdata(f1856_rdata));
  assign f1856_clk = clk;
  assign f1856_rst = rst;
  // Bindings to f1856

  // f1858
  logic [0:0] f1858_wen;
  logic [31:0] f1858_wdata;
  logic [0:0] f1858_clk;
  logic [0:0] f1858_rst;
  logic [31:0] f1858_rdata;
  sr_buffer_32_1 f1858(.wen(f1858_wen), .wdata(f1858_wdata), .clk(f1858_clk), .rst(f1858_rst), .rdata(f1858_rdata));
  assign f1858_clk = clk;
  assign f1858_rst = rst;
  // Bindings to f1858

  // f1860
  logic [0:0] f1860_wen;
  logic [31:0] f1860_wdata;
  logic [0:0] f1860_clk;
  logic [0:0] f1860_rst;
  logic [31:0] f1860_rdata;
  sr_buffer_32_1 f1860(.wen(f1860_wen), .wdata(f1860_wdata), .clk(f1860_clk), .rst(f1860_rst), .rdata(f1860_rdata));
  assign f1860_clk = clk;
  assign f1860_rst = rst;
  // Bindings to f1860

  // f1862
  logic [0:0] f1862_wen;
  logic [31:0] f1862_wdata;
  logic [0:0] f1862_clk;
  logic [0:0] f1862_rst;
  logic [31:0] f1862_rdata;
  sr_buffer_32_1 f1862(.wen(f1862_wen), .wdata(f1862_wdata), .clk(f1862_clk), .rst(f1862_rst), .rdata(f1862_rdata));
  assign f1862_clk = clk;
  assign f1862_rst = rst;
  // Bindings to f1862

  // f1864
  logic [0:0] f1864_wen;
  logic [31:0] f1864_wdata;
  logic [0:0] f1864_clk;
  logic [0:0] f1864_rst;
  logic [31:0] f1864_rdata;
  sr_buffer_32_1 f1864(.wen(f1864_wen), .wdata(f1864_wdata), .clk(f1864_clk), .rst(f1864_rst), .rdata(f1864_rdata));
  assign f1864_clk = clk;
  assign f1864_rst = rst;
  // Bindings to f1864

  // f1866
  logic [0:0] f1866_wen;
  logic [31:0] f1866_wdata;
  logic [0:0] f1866_clk;
  logic [0:0] f1866_rst;
  logic [31:0] f1866_rdata;
  sr_buffer_32_1 f1866(.wen(f1866_wen), .wdata(f1866_wdata), .clk(f1866_clk), .rst(f1866_rst), .rdata(f1866_rdata));
  assign f1866_clk = clk;
  assign f1866_rst = rst;
  // Bindings to f1866

  // f1868
  logic [0:0] f1868_wen;
  logic [31:0] f1868_wdata;
  logic [0:0] f1868_clk;
  logic [0:0] f1868_rst;
  logic [31:0] f1868_rdata;
  sr_buffer_32_1 f1868(.wen(f1868_wen), .wdata(f1868_wdata), .clk(f1868_clk), .rst(f1868_rst), .rdata(f1868_rdata));
  assign f1868_clk = clk;
  assign f1868_rst = rst;
  // Bindings to f1868

  // f1870
  logic [0:0] f1870_wen;
  logic [31:0] f1870_wdata;
  logic [0:0] f1870_clk;
  logic [0:0] f1870_rst;
  logic [31:0] f1870_rdata;
  sr_buffer_32_1 f1870(.wen(f1870_wen), .wdata(f1870_wdata), .clk(f1870_clk), .rst(f1870_rst), .rdata(f1870_rdata));
  assign f1870_clk = clk;
  assign f1870_rst = rst;
  // Bindings to f1870

  // f1872
  logic [0:0] f1872_wen;
  logic [31:0] f1872_wdata;
  logic [0:0] f1872_clk;
  logic [0:0] f1872_rst;
  logic [31:0] f1872_rdata;
  sr_buffer_32_1 f1872(.wen(f1872_wen), .wdata(f1872_wdata), .clk(f1872_clk), .rst(f1872_rst), .rdata(f1872_rdata));
  assign f1872_clk = clk;
  assign f1872_rst = rst;
  // Bindings to f1872

  // f1874
  logic [0:0] f1874_wen;
  logic [31:0] f1874_wdata;
  logic [0:0] f1874_clk;
  logic [0:0] f1874_rst;
  logic [31:0] f1874_rdata;
  sr_buffer_32_1 f1874(.wen(f1874_wen), .wdata(f1874_wdata), .clk(f1874_clk), .rst(f1874_rst), .rdata(f1874_rdata));
  assign f1874_clk = clk;
  assign f1874_rst = rst;
  // Bindings to f1874

  // f1876
  logic [0:0] f1876_wen;
  logic [31:0] f1876_wdata;
  logic [0:0] f1876_clk;
  logic [0:0] f1876_rst;
  logic [31:0] f1876_rdata;
  sr_buffer_32_1 f1876(.wen(f1876_wen), .wdata(f1876_wdata), .clk(f1876_clk), .rst(f1876_rst), .rdata(f1876_rdata));
  assign f1876_clk = clk;
  assign f1876_rst = rst;
  // Bindings to f1876

  // f1878
  logic [0:0] f1878_wen;
  logic [31:0] f1878_wdata;
  logic [0:0] f1878_clk;
  logic [0:0] f1878_rst;
  logic [31:0] f1878_rdata;
  sr_buffer_32_1 f1878(.wen(f1878_wen), .wdata(f1878_wdata), .clk(f1878_clk), .rst(f1878_rst), .rdata(f1878_rdata));
  assign f1878_clk = clk;
  assign f1878_rst = rst;
  // Bindings to f1878

  // f1880
  logic [0:0] f1880_wen;
  logic [31:0] f1880_wdata;
  logic [0:0] f1880_clk;
  logic [0:0] f1880_rst;
  logic [31:0] f1880_rdata;
  sr_buffer_32_1 f1880(.wen(f1880_wen), .wdata(f1880_wdata), .clk(f1880_clk), .rst(f1880_rst), .rdata(f1880_rdata));
  assign f1880_clk = clk;
  assign f1880_rst = rst;
  // Bindings to f1880

  // f1882
  logic [0:0] f1882_wen;
  logic [31:0] f1882_wdata;
  logic [0:0] f1882_clk;
  logic [0:0] f1882_rst;
  logic [31:0] f1882_rdata;
  sr_buffer_32_1 f1882(.wen(f1882_wen), .wdata(f1882_wdata), .clk(f1882_clk), .rst(f1882_rst), .rdata(f1882_rdata));
  assign f1882_clk = clk;
  assign f1882_rst = rst;
  // Bindings to f1882

  // f1884
  logic [0:0] f1884_wen;
  logic [31:0] f1884_wdata;
  logic [0:0] f1884_clk;
  logic [0:0] f1884_rst;
  logic [31:0] f1884_rdata;
  sr_buffer_32_1 f1884(.wen(f1884_wen), .wdata(f1884_wdata), .clk(f1884_clk), .rst(f1884_rst), .rdata(f1884_rdata));
  assign f1884_clk = clk;
  assign f1884_rst = rst;
  // Bindings to f1884

  // f1886
  logic [0:0] f1886_wen;
  logic [31:0] f1886_wdata;
  logic [0:0] f1886_clk;
  logic [0:0] f1886_rst;
  logic [31:0] f1886_rdata;
  sr_buffer_32_1 f1886(.wen(f1886_wen), .wdata(f1886_wdata), .clk(f1886_clk), .rst(f1886_rst), .rdata(f1886_rdata));
  assign f1886_clk = clk;
  assign f1886_rst = rst;
  // Bindings to f1886

  // f1888
  logic [0:0] f1888_wen;
  logic [31:0] f1888_wdata;
  logic [0:0] f1888_clk;
  logic [0:0] f1888_rst;
  logic [31:0] f1888_rdata;
  sr_buffer_32_1 f1888(.wen(f1888_wen), .wdata(f1888_wdata), .clk(f1888_clk), .rst(f1888_rst), .rdata(f1888_rdata));
  assign f1888_clk = clk;
  assign f1888_rst = rst;
  // Bindings to f1888

  // f1890
  logic [0:0] f1890_wen;
  logic [31:0] f1890_wdata;
  logic [0:0] f1890_clk;
  logic [0:0] f1890_rst;
  logic [31:0] f1890_rdata;
  sr_buffer_32_1 f1890(.wen(f1890_wen), .wdata(f1890_wdata), .clk(f1890_clk), .rst(f1890_rst), .rdata(f1890_rdata));
  assign f1890_clk = clk;
  assign f1890_rst = rst;
  // Bindings to f1890

  // f1892
  logic [0:0] f1892_wen;
  logic [31:0] f1892_wdata;
  logic [0:0] f1892_clk;
  logic [0:0] f1892_rst;
  logic [31:0] f1892_rdata;
  sr_buffer_32_1 f1892(.wen(f1892_wen), .wdata(f1892_wdata), .clk(f1892_clk), .rst(f1892_rst), .rdata(f1892_rdata));
  assign f1892_clk = clk;
  assign f1892_rst = rst;
  // Bindings to f1892

  // f1894
  logic [0:0] f1894_wen;
  logic [31:0] f1894_wdata;
  logic [0:0] f1894_clk;
  logic [0:0] f1894_rst;
  logic [31:0] f1894_rdata;
  sr_buffer_32_1 f1894(.wen(f1894_wen), .wdata(f1894_wdata), .clk(f1894_clk), .rst(f1894_rst), .rdata(f1894_rdata));
  assign f1894_clk = clk;
  assign f1894_rst = rst;
  // Bindings to f1894

  // f1896
  logic [0:0] f1896_wen;
  logic [31:0] f1896_wdata;
  logic [0:0] f1896_clk;
  logic [0:0] f1896_rst;
  logic [31:0] f1896_rdata;
  sr_buffer_32_1 f1896(.wen(f1896_wen), .wdata(f1896_wdata), .clk(f1896_clk), .rst(f1896_rst), .rdata(f1896_rdata));
  assign f1896_clk = clk;
  assign f1896_rst = rst;
  // Bindings to f1896

  // f1898
  logic [0:0] f1898_wen;
  logic [31:0] f1898_wdata;
  logic [0:0] f1898_clk;
  logic [0:0] f1898_rst;
  logic [31:0] f1898_rdata;
  sr_buffer_32_1 f1898(.wen(f1898_wen), .wdata(f1898_wdata), .clk(f1898_clk), .rst(f1898_rst), .rdata(f1898_rdata));
  assign f1898_clk = clk;
  assign f1898_rst = rst;
  // Bindings to f1898

  // f1900
  logic [0:0] f1900_wen;
  logic [31:0] f1900_wdata;
  logic [0:0] f1900_clk;
  logic [0:0] f1900_rst;
  logic [31:0] f1900_rdata;
  sr_buffer_32_1 f1900(.wen(f1900_wen), .wdata(f1900_wdata), .clk(f1900_clk), .rst(f1900_rst), .rdata(f1900_rdata));
  assign f1900_clk = clk;
  assign f1900_rst = rst;
  // Bindings to f1900

  // f1902
  logic [0:0] f1902_wen;
  logic [31:0] f1902_wdata;
  logic [0:0] f1902_clk;
  logic [0:0] f1902_rst;
  logic [31:0] f1902_rdata;
  sr_buffer_32_1 f1902(.wen(f1902_wen), .wdata(f1902_wdata), .clk(f1902_clk), .rst(f1902_rst), .rdata(f1902_rdata));
  assign f1902_clk = clk;
  assign f1902_rst = rst;
  // Bindings to f1902

  // f1904
  logic [0:0] f1904_wen;
  logic [31:0] f1904_wdata;
  logic [0:0] f1904_clk;
  logic [0:0] f1904_rst;
  logic [31:0] f1904_rdata;
  sr_buffer_32_1 f1904(.wen(f1904_wen), .wdata(f1904_wdata), .clk(f1904_clk), .rst(f1904_rst), .rdata(f1904_rdata));
  assign f1904_clk = clk;
  assign f1904_rst = rst;
  // Bindings to f1904

  // f1906
  logic [0:0] f1906_wen;
  logic [31:0] f1906_wdata;
  logic [0:0] f1906_clk;
  logic [0:0] f1906_rst;
  logic [31:0] f1906_rdata;
  sr_buffer_32_1 f1906(.wen(f1906_wen), .wdata(f1906_wdata), .clk(f1906_clk), .rst(f1906_rst), .rdata(f1906_rdata));
  assign f1906_clk = clk;
  assign f1906_rst = rst;
  // Bindings to f1906

  // f1908
  logic [0:0] f1908_wen;
  logic [31:0] f1908_wdata;
  logic [0:0] f1908_clk;
  logic [0:0] f1908_rst;
  logic [31:0] f1908_rdata;
  sr_buffer_32_1 f1908(.wen(f1908_wen), .wdata(f1908_wdata), .clk(f1908_clk), .rst(f1908_rst), .rdata(f1908_rdata));
  assign f1908_clk = clk;
  assign f1908_rst = rst;
  // Bindings to f1908

  // f1910
  logic [0:0] f1910_wen;
  logic [31:0] f1910_wdata;
  logic [0:0] f1910_clk;
  logic [0:0] f1910_rst;
  logic [31:0] f1910_rdata;
  sr_buffer_32_1 f1910(.wen(f1910_wen), .wdata(f1910_wdata), .clk(f1910_clk), .rst(f1910_rst), .rdata(f1910_rdata));
  assign f1910_clk = clk;
  assign f1910_rst = rst;
  // Bindings to f1910

  // f1912
  logic [0:0] f1912_wen;
  logic [31:0] f1912_wdata;
  logic [0:0] f1912_clk;
  logic [0:0] f1912_rst;
  logic [31:0] f1912_rdata;
  sr_buffer_32_1 f1912(.wen(f1912_wen), .wdata(f1912_wdata), .clk(f1912_clk), .rst(f1912_rst), .rdata(f1912_rdata));
  assign f1912_clk = clk;
  assign f1912_rst = rst;
  // Bindings to f1912

  // f1914
  logic [0:0] f1914_wen;
  logic [31:0] f1914_wdata;
  logic [0:0] f1914_clk;
  logic [0:0] f1914_rst;
  logic [31:0] f1914_rdata;
  sr_buffer_32_1 f1914(.wen(f1914_wen), .wdata(f1914_wdata), .clk(f1914_clk), .rst(f1914_rst), .rdata(f1914_rdata));
  assign f1914_clk = clk;
  assign f1914_rst = rst;
  // Bindings to f1914

  // f1916
  logic [0:0] f1916_wen;
  logic [31:0] f1916_wdata;
  logic [0:0] f1916_clk;
  logic [0:0] f1916_rst;
  logic [31:0] f1916_rdata;
  sr_buffer_32_1 f1916(.wen(f1916_wen), .wdata(f1916_wdata), .clk(f1916_clk), .rst(f1916_rst), .rdata(f1916_rdata));
  assign f1916_clk = clk;
  assign f1916_rst = rst;
  // Bindings to f1916

  // f1918
  logic [0:0] f1918_wen;
  logic [31:0] f1918_wdata;
  logic [0:0] f1918_clk;
  logic [0:0] f1918_rst;
  logic [31:0] f1918_rdata;
  sr_buffer_32_1 f1918(.wen(f1918_wen), .wdata(f1918_wdata), .clk(f1918_clk), .rst(f1918_rst), .rdata(f1918_rdata));
  assign f1918_clk = clk;
  assign f1918_rst = rst;
  // Bindings to f1918

  // f1920
  logic [0:0] f1920_wen;
  logic [31:0] f1920_wdata;
  logic [0:0] f1920_clk;
  logic [0:0] f1920_rst;
  logic [31:0] f1920_rdata;
  sr_buffer_32_1 f1920(.wen(f1920_wen), .wdata(f1920_wdata), .clk(f1920_clk), .rst(f1920_rst), .rdata(f1920_rdata));
  assign f1920_clk = clk;
  assign f1920_rst = rst;
  // Bindings to f1920

  // f1922
  logic [0:0] f1922_wen;
  logic [31:0] f1922_wdata;
  logic [0:0] f1922_clk;
  logic [0:0] f1922_rst;
  logic [31:0] f1922_rdata;
  sr_buffer_32_1 f1922(.wen(f1922_wen), .wdata(f1922_wdata), .clk(f1922_clk), .rst(f1922_rst), .rdata(f1922_rdata));
  assign f1922_clk = clk;
  assign f1922_rst = rst;
  // Bindings to f1922

  // f1924
  logic [0:0] f1924_wen;
  logic [31:0] f1924_wdata;
  logic [0:0] f1924_clk;
  logic [0:0] f1924_rst;
  logic [31:0] f1924_rdata;
  sr_buffer_32_1 f1924(.wen(f1924_wen), .wdata(f1924_wdata), .clk(f1924_clk), .rst(f1924_rst), .rdata(f1924_rdata));
  assign f1924_clk = clk;
  assign f1924_rst = rst;
  // Bindings to f1924

  // f1926
  logic [0:0] f1926_wen;
  logic [31:0] f1926_wdata;
  logic [0:0] f1926_clk;
  logic [0:0] f1926_rst;
  logic [31:0] f1926_rdata;
  sr_buffer_32_1 f1926(.wen(f1926_wen), .wdata(f1926_wdata), .clk(f1926_clk), .rst(f1926_rst), .rdata(f1926_rdata));
  assign f1926_clk = clk;
  assign f1926_rst = rst;
  // Bindings to f1926

  // f1928
  logic [0:0] f1928_wen;
  logic [31:0] f1928_wdata;
  logic [0:0] f1928_clk;
  logic [0:0] f1928_rst;
  logic [31:0] f1928_rdata;
  sr_buffer_32_1 f1928(.wen(f1928_wen), .wdata(f1928_wdata), .clk(f1928_clk), .rst(f1928_rst), .rdata(f1928_rdata));
  assign f1928_clk = clk;
  assign f1928_rst = rst;
  // Bindings to f1928

  // f1930
  logic [0:0] f1930_wen;
  logic [31:0] f1930_wdata;
  logic [0:0] f1930_clk;
  logic [0:0] f1930_rst;
  logic [31:0] f1930_rdata;
  sr_buffer_32_1 f1930(.wen(f1930_wen), .wdata(f1930_wdata), .clk(f1930_clk), .rst(f1930_rst), .rdata(f1930_rdata));
  assign f1930_clk = clk;
  assign f1930_rst = rst;
  // Bindings to f1930

  // f1932
  logic [0:0] f1932_wen;
  logic [31:0] f1932_wdata;
  logic [0:0] f1932_clk;
  logic [0:0] f1932_rst;
  logic [31:0] f1932_rdata;
  sr_buffer_32_1 f1932(.wen(f1932_wen), .wdata(f1932_wdata), .clk(f1932_clk), .rst(f1932_rst), .rdata(f1932_rdata));
  assign f1932_clk = clk;
  assign f1932_rst = rst;
  // Bindings to f1932

  // f1934
  logic [0:0] f1934_wen;
  logic [31:0] f1934_wdata;
  logic [0:0] f1934_clk;
  logic [0:0] f1934_rst;
  logic [31:0] f1934_rdata;
  sr_buffer_32_1 f1934(.wen(f1934_wen), .wdata(f1934_wdata), .clk(f1934_clk), .rst(f1934_rst), .rdata(f1934_rdata));
  assign f1934_clk = clk;
  assign f1934_rst = rst;
  // Bindings to f1934

  // f1936
  logic [0:0] f1936_wen;
  logic [31:0] f1936_wdata;
  logic [0:0] f1936_clk;
  logic [0:0] f1936_rst;
  logic [31:0] f1936_rdata;
  sr_buffer_32_1 f1936(.wen(f1936_wen), .wdata(f1936_wdata), .clk(f1936_clk), .rst(f1936_rst), .rdata(f1936_rdata));
  assign f1936_clk = clk;
  assign f1936_rst = rst;
  // Bindings to f1936

  // f1938
  logic [0:0] f1938_wen;
  logic [31:0] f1938_wdata;
  logic [0:0] f1938_clk;
  logic [0:0] f1938_rst;
  logic [31:0] f1938_rdata;
  sr_buffer_32_1 f1938(.wen(f1938_wen), .wdata(f1938_wdata), .clk(f1938_clk), .rst(f1938_rst), .rdata(f1938_rdata));
  assign f1938_clk = clk;
  assign f1938_rst = rst;
  // Bindings to f1938

  // f1940
  logic [0:0] f1940_wen;
  logic [31:0] f1940_wdata;
  logic [0:0] f1940_clk;
  logic [0:0] f1940_rst;
  logic [31:0] f1940_rdata;
  sr_buffer_32_1 f1940(.wen(f1940_wen), .wdata(f1940_wdata), .clk(f1940_clk), .rst(f1940_rst), .rdata(f1940_rdata));
  assign f1940_clk = clk;
  assign f1940_rst = rst;
  // Bindings to f1940

  // f1942
  logic [0:0] f1942_wen;
  logic [31:0] f1942_wdata;
  logic [0:0] f1942_clk;
  logic [0:0] f1942_rst;
  logic [31:0] f1942_rdata;
  sr_buffer_32_1 f1942(.wen(f1942_wen), .wdata(f1942_wdata), .clk(f1942_clk), .rst(f1942_rst), .rdata(f1942_rdata));
  assign f1942_clk = clk;
  assign f1942_rst = rst;
  // Bindings to f1942

  // f1944
  logic [0:0] f1944_wen;
  logic [31:0] f1944_wdata;
  logic [0:0] f1944_clk;
  logic [0:0] f1944_rst;
  logic [31:0] f1944_rdata;
  sr_buffer_32_1 f1944(.wen(f1944_wen), .wdata(f1944_wdata), .clk(f1944_clk), .rst(f1944_rst), .rdata(f1944_rdata));
  assign f1944_clk = clk;
  assign f1944_rst = rst;
  // Bindings to f1944

  // f1946
  logic [0:0] f1946_wen;
  logic [31:0] f1946_wdata;
  logic [0:0] f1946_clk;
  logic [0:0] f1946_rst;
  logic [31:0] f1946_rdata;
  sr_buffer_32_1 f1946(.wen(f1946_wen), .wdata(f1946_wdata), .clk(f1946_clk), .rst(f1946_rst), .rdata(f1946_rdata));
  assign f1946_clk = clk;
  assign f1946_rst = rst;
  // Bindings to f1946

  // f1948
  logic [0:0] f1948_wen;
  logic [31:0] f1948_wdata;
  logic [0:0] f1948_clk;
  logic [0:0] f1948_rst;
  logic [31:0] f1948_rdata;
  sr_buffer_32_1 f1948(.wen(f1948_wen), .wdata(f1948_wdata), .clk(f1948_clk), .rst(f1948_rst), .rdata(f1948_rdata));
  assign f1948_clk = clk;
  assign f1948_rst = rst;
  // Bindings to f1948

  // f1950
  logic [0:0] f1950_wen;
  logic [31:0] f1950_wdata;
  logic [0:0] f1950_clk;
  logic [0:0] f1950_rst;
  logic [31:0] f1950_rdata;
  sr_buffer_32_1 f1950(.wen(f1950_wen), .wdata(f1950_wdata), .clk(f1950_clk), .rst(f1950_rst), .rdata(f1950_rdata));
  assign f1950_clk = clk;
  assign f1950_rst = rst;
  // Bindings to f1950

  // f1952
  logic [0:0] f1952_wen;
  logic [31:0] f1952_wdata;
  logic [0:0] f1952_clk;
  logic [0:0] f1952_rst;
  logic [31:0] f1952_rdata;
  sr_buffer_32_1 f1952(.wen(f1952_wen), .wdata(f1952_wdata), .clk(f1952_clk), .rst(f1952_rst), .rdata(f1952_rdata));
  assign f1952_clk = clk;
  assign f1952_rst = rst;
  // Bindings to f1952

  // f1954
  logic [0:0] f1954_wen;
  logic [31:0] f1954_wdata;
  logic [0:0] f1954_clk;
  logic [0:0] f1954_rst;
  logic [31:0] f1954_rdata;
  sr_buffer_32_1 f1954(.wen(f1954_wen), .wdata(f1954_wdata), .clk(f1954_clk), .rst(f1954_rst), .rdata(f1954_rdata));
  assign f1954_clk = clk;
  assign f1954_rst = rst;
  // Bindings to f1954

  // f1956
  logic [0:0] f1956_wen;
  logic [31:0] f1956_wdata;
  logic [0:0] f1956_clk;
  logic [0:0] f1956_rst;
  logic [31:0] f1956_rdata;
  sr_buffer_32_1 f1956(.wen(f1956_wen), .wdata(f1956_wdata), .clk(f1956_clk), .rst(f1956_rst), .rdata(f1956_rdata));
  assign f1956_clk = clk;
  assign f1956_rst = rst;
  // Bindings to f1956

  // f1958
  logic [0:0] f1958_wen;
  logic [31:0] f1958_wdata;
  logic [0:0] f1958_clk;
  logic [0:0] f1958_rst;
  logic [31:0] f1958_rdata;
  sr_buffer_32_1 f1958(.wen(f1958_wen), .wdata(f1958_wdata), .clk(f1958_clk), .rst(f1958_rst), .rdata(f1958_rdata));
  assign f1958_clk = clk;
  assign f1958_rst = rst;
  // Bindings to f1958

  // f1960
  logic [0:0] f1960_wen;
  logic [31:0] f1960_wdata;
  logic [0:0] f1960_clk;
  logic [0:0] f1960_rst;
  logic [31:0] f1960_rdata;
  sr_buffer_32_1 f1960(.wen(f1960_wen), .wdata(f1960_wdata), .clk(f1960_clk), .rst(f1960_rst), .rdata(f1960_rdata));
  assign f1960_clk = clk;
  assign f1960_rst = rst;
  // Bindings to f1960

  // f1962
  logic [0:0] f1962_wen;
  logic [31:0] f1962_wdata;
  logic [0:0] f1962_clk;
  logic [0:0] f1962_rst;
  logic [31:0] f1962_rdata;
  sr_buffer_32_1 f1962(.wen(f1962_wen), .wdata(f1962_wdata), .clk(f1962_clk), .rst(f1962_rst), .rdata(f1962_rdata));
  assign f1962_clk = clk;
  assign f1962_rst = rst;
  // Bindings to f1962

  // f1964
  logic [0:0] f1964_wen;
  logic [31:0] f1964_wdata;
  logic [0:0] f1964_clk;
  logic [0:0] f1964_rst;
  logic [31:0] f1964_rdata;
  sr_buffer_32_1 f1964(.wen(f1964_wen), .wdata(f1964_wdata), .clk(f1964_clk), .rst(f1964_rst), .rdata(f1964_rdata));
  assign f1964_clk = clk;
  assign f1964_rst = rst;
  // Bindings to f1964

  // f1966
  logic [0:0] f1966_wen;
  logic [31:0] f1966_wdata;
  logic [0:0] f1966_clk;
  logic [0:0] f1966_rst;
  logic [31:0] f1966_rdata;
  sr_buffer_32_1 f1966(.wen(f1966_wen), .wdata(f1966_wdata), .clk(f1966_clk), .rst(f1966_rst), .rdata(f1966_rdata));
  assign f1966_clk = clk;
  assign f1966_rst = rst;
  // Bindings to f1966

  // f1968
  logic [0:0] f1968_wen;
  logic [31:0] f1968_wdata;
  logic [0:0] f1968_clk;
  logic [0:0] f1968_rst;
  logic [31:0] f1968_rdata;
  sr_buffer_32_1 f1968(.wen(f1968_wen), .wdata(f1968_wdata), .clk(f1968_clk), .rst(f1968_rst), .rdata(f1968_rdata));
  assign f1968_clk = clk;
  assign f1968_rst = rst;
  // Bindings to f1968

  // f1970
  logic [0:0] f1970_wen;
  logic [31:0] f1970_wdata;
  logic [0:0] f1970_clk;
  logic [0:0] f1970_rst;
  logic [31:0] f1970_rdata;
  sr_buffer_32_1 f1970(.wen(f1970_wen), .wdata(f1970_wdata), .clk(f1970_clk), .rst(f1970_rst), .rdata(f1970_rdata));
  assign f1970_clk = clk;
  assign f1970_rst = rst;
  // Bindings to f1970

  // f1972
  logic [0:0] f1972_wen;
  logic [31:0] f1972_wdata;
  logic [0:0] f1972_clk;
  logic [0:0] f1972_rst;
  logic [31:0] f1972_rdata;
  sr_buffer_32_1 f1972(.wen(f1972_wen), .wdata(f1972_wdata), .clk(f1972_clk), .rst(f1972_rst), .rdata(f1972_rdata));
  assign f1972_clk = clk;
  assign f1972_rst = rst;
  // Bindings to f1972

  // f1974
  logic [0:0] f1974_wen;
  logic [31:0] f1974_wdata;
  logic [0:0] f1974_clk;
  logic [0:0] f1974_rst;
  logic [31:0] f1974_rdata;
  sr_buffer_32_1 f1974(.wen(f1974_wen), .wdata(f1974_wdata), .clk(f1974_clk), .rst(f1974_rst), .rdata(f1974_rdata));
  assign f1974_clk = clk;
  assign f1974_rst = rst;
  // Bindings to f1974

  // f1976
  logic [0:0] f1976_wen;
  logic [31:0] f1976_wdata;
  logic [0:0] f1976_clk;
  logic [0:0] f1976_rst;
  logic [31:0] f1976_rdata;
  sr_buffer_32_1 f1976(.wen(f1976_wen), .wdata(f1976_wdata), .clk(f1976_clk), .rst(f1976_rst), .rdata(f1976_rdata));
  assign f1976_clk = clk;
  assign f1976_rst = rst;
  // Bindings to f1976

  // f1978
  logic [0:0] f1978_wen;
  logic [31:0] f1978_wdata;
  logic [0:0] f1978_clk;
  logic [0:0] f1978_rst;
  logic [31:0] f1978_rdata;
  sr_buffer_32_1 f1978(.wen(f1978_wen), .wdata(f1978_wdata), .clk(f1978_clk), .rst(f1978_rst), .rdata(f1978_rdata));
  assign f1978_clk = clk;
  assign f1978_rst = rst;
  // Bindings to f1978

  // f1980
  logic [0:0] f1980_wen;
  logic [31:0] f1980_wdata;
  logic [0:0] f1980_clk;
  logic [0:0] f1980_rst;
  logic [31:0] f1980_rdata;
  sr_buffer_32_1 f1980(.wen(f1980_wen), .wdata(f1980_wdata), .clk(f1980_clk), .rst(f1980_rst), .rdata(f1980_rdata));
  assign f1980_clk = clk;
  assign f1980_rst = rst;
  // Bindings to f1980

  // f1982
  logic [0:0] f1982_wen;
  logic [31:0] f1982_wdata;
  logic [0:0] f1982_clk;
  logic [0:0] f1982_rst;
  logic [31:0] f1982_rdata;
  sr_buffer_32_1 f1982(.wen(f1982_wen), .wdata(f1982_wdata), .clk(f1982_clk), .rst(f1982_rst), .rdata(f1982_rdata));
  assign f1982_clk = clk;
  assign f1982_rst = rst;
  // Bindings to f1982

  // f1984
  logic [0:0] f1984_wen;
  logic [31:0] f1984_wdata;
  logic [0:0] f1984_clk;
  logic [0:0] f1984_rst;
  logic [31:0] f1984_rdata;
  sr_buffer_32_1 f1984(.wen(f1984_wen), .wdata(f1984_wdata), .clk(f1984_clk), .rst(f1984_rst), .rdata(f1984_rdata));
  assign f1984_clk = clk;
  assign f1984_rst = rst;
  // Bindings to f1984

  // f1986
  logic [0:0] f1986_wen;
  logic [31:0] f1986_wdata;
  logic [0:0] f1986_clk;
  logic [0:0] f1986_rst;
  logic [31:0] f1986_rdata;
  sr_buffer_32_1 f1986(.wen(f1986_wen), .wdata(f1986_wdata), .clk(f1986_clk), .rst(f1986_rst), .rdata(f1986_rdata));
  assign f1986_clk = clk;
  assign f1986_rst = rst;
  // Bindings to f1986

  // f1988
  logic [0:0] f1988_wen;
  logic [31:0] f1988_wdata;
  logic [0:0] f1988_clk;
  logic [0:0] f1988_rst;
  logic [31:0] f1988_rdata;
  sr_buffer_32_1 f1988(.wen(f1988_wen), .wdata(f1988_wdata), .clk(f1988_clk), .rst(f1988_rst), .rdata(f1988_rdata));
  assign f1988_clk = clk;
  assign f1988_rst = rst;
  // Bindings to f1988

  // f1990
  logic [0:0] f1990_wen;
  logic [31:0] f1990_wdata;
  logic [0:0] f1990_clk;
  logic [0:0] f1990_rst;
  logic [31:0] f1990_rdata;
  sr_buffer_32_1 f1990(.wen(f1990_wen), .wdata(f1990_wdata), .clk(f1990_clk), .rst(f1990_rst), .rdata(f1990_rdata));
  assign f1990_clk = clk;
  assign f1990_rst = rst;
  // Bindings to f1990

  // f1992
  logic [0:0] f1992_wen;
  logic [31:0] f1992_wdata;
  logic [0:0] f1992_clk;
  logic [0:0] f1992_rst;
  logic [31:0] f1992_rdata;
  sr_buffer_32_1 f1992(.wen(f1992_wen), .wdata(f1992_wdata), .clk(f1992_clk), .rst(f1992_rst), .rdata(f1992_rdata));
  assign f1992_clk = clk;
  assign f1992_rst = rst;
  // Bindings to f1992

  // f1994
  logic [0:0] f1994_wen;
  logic [31:0] f1994_wdata;
  logic [0:0] f1994_clk;
  logic [0:0] f1994_rst;
  logic [31:0] f1994_rdata;
  sr_buffer_32_1 f1994(.wen(f1994_wen), .wdata(f1994_wdata), .clk(f1994_clk), .rst(f1994_rst), .rdata(f1994_rdata));
  assign f1994_clk = clk;
  assign f1994_rst = rst;
  // Bindings to f1994

  // f1996
  logic [0:0] f1996_wen;
  logic [31:0] f1996_wdata;
  logic [0:0] f1996_clk;
  logic [0:0] f1996_rst;
  logic [31:0] f1996_rdata;
  sr_buffer_32_1 f1996(.wen(f1996_wen), .wdata(f1996_wdata), .clk(f1996_clk), .rst(f1996_rst), .rdata(f1996_rdata));
  assign f1996_clk = clk;
  assign f1996_rst = rst;
  // Bindings to f1996

  // f1998
  logic [0:0] f1998_wen;
  logic [31:0] f1998_wdata;
  logic [0:0] f1998_clk;
  logic [0:0] f1998_rst;
  logic [31:0] f1998_rdata;
  sr_buffer_32_1 f1998(.wen(f1998_wen), .wdata(f1998_wdata), .clk(f1998_clk), .rst(f1998_rst), .rdata(f1998_rdata));
  assign f1998_clk = clk;
  assign f1998_rst = rst;
  // Bindings to f1998

  // f2000
  logic [0:0] f2000_wen;
  logic [31:0] f2000_wdata;
  logic [0:0] f2000_clk;
  logic [0:0] f2000_rst;
  logic [31:0] f2000_rdata;
  sr_buffer_32_1 f2000(.wen(f2000_wen), .wdata(f2000_wdata), .clk(f2000_clk), .rst(f2000_rst), .rdata(f2000_rdata));
  assign f2000_clk = clk;
  assign f2000_rst = rst;
  // Bindings to f2000

  // f2002
  logic [0:0] f2002_wen;
  logic [31:0] f2002_wdata;
  logic [0:0] f2002_clk;
  logic [0:0] f2002_rst;
  logic [31:0] f2002_rdata;
  sr_buffer_32_1 f2002(.wen(f2002_wen), .wdata(f2002_wdata), .clk(f2002_clk), .rst(f2002_rst), .rdata(f2002_rdata));
  assign f2002_clk = clk;
  assign f2002_rst = rst;
  // Bindings to f2002

  // f2004
  logic [0:0] f2004_wen;
  logic [31:0] f2004_wdata;
  logic [0:0] f2004_clk;
  logic [0:0] f2004_rst;
  logic [31:0] f2004_rdata;
  sr_buffer_32_1 f2004(.wen(f2004_wen), .wdata(f2004_wdata), .clk(f2004_clk), .rst(f2004_rst), .rdata(f2004_rdata));
  assign f2004_clk = clk;
  assign f2004_rst = rst;
  // Bindings to f2004

  // f2006
  logic [0:0] f2006_wen;
  logic [31:0] f2006_wdata;
  logic [0:0] f2006_clk;
  logic [0:0] f2006_rst;
  logic [31:0] f2006_rdata;
  sr_buffer_32_1 f2006(.wen(f2006_wen), .wdata(f2006_wdata), .clk(f2006_clk), .rst(f2006_rst), .rdata(f2006_rdata));
  assign f2006_clk = clk;
  assign f2006_rst = rst;
  // Bindings to f2006

  // f2008
  logic [0:0] f2008_wen;
  logic [31:0] f2008_wdata;
  logic [0:0] f2008_clk;
  logic [0:0] f2008_rst;
  logic [31:0] f2008_rdata;
  sr_buffer_32_1 f2008(.wen(f2008_wen), .wdata(f2008_wdata), .clk(f2008_clk), .rst(f2008_rst), .rdata(f2008_rdata));
  assign f2008_clk = clk;
  assign f2008_rst = rst;
  // Bindings to f2008

  // f2010
  logic [0:0] f2010_wen;
  logic [31:0] f2010_wdata;
  logic [0:0] f2010_clk;
  logic [0:0] f2010_rst;
  logic [31:0] f2010_rdata;
  sr_buffer_32_1 f2010(.wen(f2010_wen), .wdata(f2010_wdata), .clk(f2010_clk), .rst(f2010_rst), .rdata(f2010_rdata));
  assign f2010_clk = clk;
  assign f2010_rst = rst;
  // Bindings to f2010

  // f2012
  logic [0:0] f2012_wen;
  logic [31:0] f2012_wdata;
  logic [0:0] f2012_clk;
  logic [0:0] f2012_rst;
  logic [31:0] f2012_rdata;
  sr_buffer_32_1 f2012(.wen(f2012_wen), .wdata(f2012_wdata), .clk(f2012_clk), .rst(f2012_rst), .rdata(f2012_rdata));
  assign f2012_clk = clk;
  assign f2012_rst = rst;
  // Bindings to f2012

  // f2014
  logic [0:0] f2014_wen;
  logic [31:0] f2014_wdata;
  logic [0:0] f2014_clk;
  logic [0:0] f2014_rst;
  logic [31:0] f2014_rdata;
  sr_buffer_32_1 f2014(.wen(f2014_wen), .wdata(f2014_wdata), .clk(f2014_clk), .rst(f2014_rst), .rdata(f2014_rdata));
  assign f2014_clk = clk;
  assign f2014_rst = rst;
  // Bindings to f2014

  // f2016
  logic [0:0] f2016_wen;
  logic [31:0] f2016_wdata;
  logic [0:0] f2016_clk;
  logic [0:0] f2016_rst;
  logic [31:0] f2016_rdata;
  sr_buffer_32_1 f2016(.wen(f2016_wen), .wdata(f2016_wdata), .clk(f2016_clk), .rst(f2016_rst), .rdata(f2016_rdata));
  assign f2016_clk = clk;
  assign f2016_rst = rst;
  // Bindings to f2016

  // f2018
  logic [0:0] f2018_wen;
  logic [31:0] f2018_wdata;
  logic [0:0] f2018_clk;
  logic [0:0] f2018_rst;
  logic [31:0] f2018_rdata;
  sr_buffer_32_1 f2018(.wen(f2018_wen), .wdata(f2018_wdata), .clk(f2018_clk), .rst(f2018_rst), .rdata(f2018_rdata));
  assign f2018_clk = clk;
  assign f2018_rst = rst;
  // Bindings to f2018

  // f2020
  logic [0:0] f2020_wen;
  logic [31:0] f2020_wdata;
  logic [0:0] f2020_clk;
  logic [0:0] f2020_rst;
  logic [31:0] f2020_rdata;
  sr_buffer_32_1 f2020(.wen(f2020_wen), .wdata(f2020_wdata), .clk(f2020_clk), .rst(f2020_rst), .rdata(f2020_rdata));
  assign f2020_clk = clk;
  assign f2020_rst = rst;
  // Bindings to f2020

  // f2022
  logic [0:0] f2022_wen;
  logic [31:0] f2022_wdata;
  logic [0:0] f2022_clk;
  logic [0:0] f2022_rst;
  logic [31:0] f2022_rdata;
  sr_buffer_32_1 f2022(.wen(f2022_wen), .wdata(f2022_wdata), .clk(f2022_clk), .rst(f2022_rst), .rdata(f2022_rdata));
  assign f2022_clk = clk;
  assign f2022_rst = rst;
  // Bindings to f2022

  // f2024
  logic [0:0] f2024_wen;
  logic [31:0] f2024_wdata;
  logic [0:0] f2024_clk;
  logic [0:0] f2024_rst;
  logic [31:0] f2024_rdata;
  sr_buffer_32_1 f2024(.wen(f2024_wen), .wdata(f2024_wdata), .clk(f2024_clk), .rst(f2024_rst), .rdata(f2024_rdata));
  assign f2024_clk = clk;
  assign f2024_rst = rst;
  // Bindings to f2024

  // f2026
  logic [0:0] f2026_wen;
  logic [31:0] f2026_wdata;
  logic [0:0] f2026_clk;
  logic [0:0] f2026_rst;
  logic [31:0] f2026_rdata;
  sr_buffer_32_1 f2026(.wen(f2026_wen), .wdata(f2026_wdata), .clk(f2026_clk), .rst(f2026_rst), .rdata(f2026_rdata));
  assign f2026_clk = clk;
  assign f2026_rst = rst;
  // Bindings to f2026

  // f2028
  logic [0:0] f2028_wen;
  logic [31:0] f2028_wdata;
  logic [0:0] f2028_clk;
  logic [0:0] f2028_rst;
  logic [31:0] f2028_rdata;
  sr_buffer_32_1 f2028(.wen(f2028_wen), .wdata(f2028_wdata), .clk(f2028_clk), .rst(f2028_rst), .rdata(f2028_rdata));
  assign f2028_clk = clk;
  assign f2028_rst = rst;
  // Bindings to f2028

  // f2030
  logic [0:0] f2030_wen;
  logic [31:0] f2030_wdata;
  logic [0:0] f2030_clk;
  logic [0:0] f2030_rst;
  logic [31:0] f2030_rdata;
  sr_buffer_32_1 f2030(.wen(f2030_wen), .wdata(f2030_wdata), .clk(f2030_clk), .rst(f2030_rst), .rdata(f2030_rdata));
  assign f2030_clk = clk;
  assign f2030_rst = rst;
  // Bindings to f2030

  // f2032
  logic [0:0] f2032_wen;
  logic [31:0] f2032_wdata;
  logic [0:0] f2032_clk;
  logic [0:0] f2032_rst;
  logic [31:0] f2032_rdata;
  sr_buffer_32_1 f2032(.wen(f2032_wen), .wdata(f2032_wdata), .clk(f2032_clk), .rst(f2032_rst), .rdata(f2032_rdata));
  assign f2032_clk = clk;
  assign f2032_rst = rst;
  // Bindings to f2032

  // f2034
  logic [0:0] f2034_wen;
  logic [31:0] f2034_wdata;
  logic [0:0] f2034_clk;
  logic [0:0] f2034_rst;
  logic [31:0] f2034_rdata;
  sr_buffer_32_1 f2034(.wen(f2034_wen), .wdata(f2034_wdata), .clk(f2034_clk), .rst(f2034_rst), .rdata(f2034_rdata));
  assign f2034_clk = clk;
  assign f2034_rst = rst;
  // Bindings to f2034

  // f2036
  logic [0:0] f2036_wen;
  logic [31:0] f2036_wdata;
  logic [0:0] f2036_clk;
  logic [0:0] f2036_rst;
  logic [31:0] f2036_rdata;
  sr_buffer_32_1 f2036(.wen(f2036_wen), .wdata(f2036_wdata), .clk(f2036_clk), .rst(f2036_rst), .rdata(f2036_rdata));
  assign f2036_clk = clk;
  assign f2036_rst = rst;
  // Bindings to f2036

  // f2038
  logic [0:0] f2038_wen;
  logic [31:0] f2038_wdata;
  logic [0:0] f2038_clk;
  logic [0:0] f2038_rst;
  logic [31:0] f2038_rdata;
  sr_buffer_32_1 f2038(.wen(f2038_wen), .wdata(f2038_wdata), .clk(f2038_clk), .rst(f2038_rst), .rdata(f2038_rdata));
  assign f2038_clk = clk;
  assign f2038_rst = rst;
  // Bindings to f2038

  // f2040
  logic [0:0] f2040_wen;
  logic [31:0] f2040_wdata;
  logic [0:0] f2040_clk;
  logic [0:0] f2040_rst;
  logic [31:0] f2040_rdata;
  sr_buffer_32_1 f2040(.wen(f2040_wen), .wdata(f2040_wdata), .clk(f2040_clk), .rst(f2040_rst), .rdata(f2040_rdata));
  assign f2040_clk = clk;
  assign f2040_rst = rst;
  // Bindings to f2040

  // f2042
  logic [0:0] f2042_wen;
  logic [31:0] f2042_wdata;
  logic [0:0] f2042_clk;
  logic [0:0] f2042_rst;
  logic [31:0] f2042_rdata;
  sr_buffer_32_1 f2042(.wen(f2042_wen), .wdata(f2042_wdata), .clk(f2042_clk), .rst(f2042_rst), .rdata(f2042_rdata));
  assign f2042_clk = clk;
  assign f2042_rst = rst;
  // Bindings to f2042

  // f2044
  logic [0:0] f2044_wen;
  logic [31:0] f2044_wdata;
  logic [0:0] f2044_clk;
  logic [0:0] f2044_rst;
  logic [31:0] f2044_rdata;
  sr_buffer_32_1 f2044(.wen(f2044_wen), .wdata(f2044_wdata), .clk(f2044_clk), .rst(f2044_rst), .rdata(f2044_rdata));
  assign f2044_clk = clk;
  assign f2044_rst = rst;
  // Bindings to f2044

  // f2046
  logic [0:0] f2046_wen;
  logic [31:0] f2046_wdata;
  logic [0:0] f2046_clk;
  logic [0:0] f2046_rst;
  logic [31:0] f2046_rdata;
  sr_buffer_32_1 f2046(.wen(f2046_wen), .wdata(f2046_wdata), .clk(f2046_clk), .rst(f2046_rst), .rdata(f2046_rdata));
  assign f2046_clk = clk;
  assign f2046_rst = rst;
  // Bindings to f2046

  // f2048
  logic [0:0] f2048_wen;
  logic [31:0] f2048_wdata;
  logic [0:0] f2048_clk;
  logic [0:0] f2048_rst;
  logic [31:0] f2048_rdata;
  sr_buffer_32_1 f2048(.wen(f2048_wen), .wdata(f2048_wdata), .clk(f2048_clk), .rst(f2048_rst), .rdata(f2048_rdata));
  assign f2048_clk = clk;
  assign f2048_rst = rst;
  // Bindings to f2048

  // f2050
  logic [0:0] f2050_wen;
  logic [31:0] f2050_wdata;
  logic [0:0] f2050_clk;
  logic [0:0] f2050_rst;
  logic [31:0] f2050_rdata;
  sr_buffer_32_1 f2050(.wen(f2050_wen), .wdata(f2050_wdata), .clk(f2050_clk), .rst(f2050_rst), .rdata(f2050_rdata));
  assign f2050_clk = clk;
  assign f2050_rst = rst;
  // Bindings to f2050

  // f2052
  logic [0:0] f2052_wen;
  logic [31:0] f2052_wdata;
  logic [0:0] f2052_clk;
  logic [0:0] f2052_rst;
  logic [31:0] f2052_rdata;
  sr_buffer_32_1 f2052(.wen(f2052_wen), .wdata(f2052_wdata), .clk(f2052_clk), .rst(f2052_rst), .rdata(f2052_rdata));
  assign f2052_clk = clk;
  assign f2052_rst = rst;
  // Bindings to f2052

  // f2054
  logic [0:0] f2054_wen;
  logic [31:0] f2054_wdata;
  logic [0:0] f2054_clk;
  logic [0:0] f2054_rst;
  logic [31:0] f2054_rdata;
  sr_buffer_32_1 f2054(.wen(f2054_wen), .wdata(f2054_wdata), .clk(f2054_clk), .rst(f2054_rst), .rdata(f2054_rdata));
  assign f2054_clk = clk;
  assign f2054_rst = rst;
  // Bindings to f2054

  // f2056
  logic [0:0] f2056_wen;
  logic [31:0] f2056_wdata;
  logic [0:0] f2056_clk;
  logic [0:0] f2056_rst;
  logic [31:0] f2056_rdata;
  sr_buffer_32_1 f2056(.wen(f2056_wen), .wdata(f2056_wdata), .clk(f2056_clk), .rst(f2056_rst), .rdata(f2056_rdata));
  assign f2056_clk = clk;
  assign f2056_rst = rst;
  // Bindings to f2056

  // f2058
  logic [0:0] f2058_wen;
  logic [31:0] f2058_wdata;
  logic [0:0] f2058_clk;
  logic [0:0] f2058_rst;
  logic [31:0] f2058_rdata;
  sr_buffer_32_1 f2058(.wen(f2058_wen), .wdata(f2058_wdata), .clk(f2058_clk), .rst(f2058_rst), .rdata(f2058_rdata));
  assign f2058_clk = clk;
  assign f2058_rst = rst;
  // Bindings to f2058

  // f2060
  logic [0:0] f2060_wen;
  logic [31:0] f2060_wdata;
  logic [0:0] f2060_clk;
  logic [0:0] f2060_rst;
  logic [31:0] f2060_rdata;
  sr_buffer_32_1 f2060(.wen(f2060_wen), .wdata(f2060_wdata), .clk(f2060_clk), .rst(f2060_rst), .rdata(f2060_rdata));
  assign f2060_clk = clk;
  assign f2060_rst = rst;
  // Bindings to f2060

  // f2062
  logic [0:0] f2062_wen;
  logic [31:0] f2062_wdata;
  logic [0:0] f2062_clk;
  logic [0:0] f2062_rst;
  logic [31:0] f2062_rdata;
  sr_buffer_32_1 f2062(.wen(f2062_wen), .wdata(f2062_wdata), .clk(f2062_clk), .rst(f2062_rst), .rdata(f2062_rdata));
  assign f2062_clk = clk;
  assign f2062_rst = rst;
  // Bindings to f2062

  // f2064
  logic [0:0] f2064_wen;
  logic [31:0] f2064_wdata;
  logic [0:0] f2064_clk;
  logic [0:0] f2064_rst;
  logic [31:0] f2064_rdata;
  sr_buffer_32_1 f2064(.wen(f2064_wen), .wdata(f2064_wdata), .clk(f2064_clk), .rst(f2064_rst), .rdata(f2064_rdata));
  assign f2064_clk = clk;
  assign f2064_rst = rst;
  // Bindings to f2064

  // f2066
  logic [0:0] f2066_wen;
  logic [31:0] f2066_wdata;
  logic [0:0] f2066_clk;
  logic [0:0] f2066_rst;
  logic [31:0] f2066_rdata;
  sr_buffer_32_1 f2066(.wen(f2066_wen), .wdata(f2066_wdata), .clk(f2066_clk), .rst(f2066_rst), .rdata(f2066_rdata));
  assign f2066_clk = clk;
  assign f2066_rst = rst;
  // Bindings to f2066

  // f2068
  logic [0:0] f2068_wen;
  logic [31:0] f2068_wdata;
  logic [0:0] f2068_clk;
  logic [0:0] f2068_rst;
  logic [31:0] f2068_rdata;
  sr_buffer_32_1 f2068(.wen(f2068_wen), .wdata(f2068_wdata), .clk(f2068_clk), .rst(f2068_rst), .rdata(f2068_rdata));
  assign f2068_clk = clk;
  assign f2068_rst = rst;
  // Bindings to f2068

  // f2070
  logic [0:0] f2070_wen;
  logic [31:0] f2070_wdata;
  logic [0:0] f2070_clk;
  logic [0:0] f2070_rst;
  logic [31:0] f2070_rdata;
  sr_buffer_32_1 f2070(.wen(f2070_wen), .wdata(f2070_wdata), .clk(f2070_clk), .rst(f2070_rst), .rdata(f2070_rdata));
  assign f2070_clk = clk;
  assign f2070_rst = rst;
  // Bindings to f2070

  // f2072
  logic [0:0] f2072_wen;
  logic [31:0] f2072_wdata;
  logic [0:0] f2072_clk;
  logic [0:0] f2072_rst;
  logic [31:0] f2072_rdata;
  sr_buffer_32_1 f2072(.wen(f2072_wen), .wdata(f2072_wdata), .clk(f2072_clk), .rst(f2072_rst), .rdata(f2072_rdata));
  assign f2072_clk = clk;
  assign f2072_rst = rst;
  // Bindings to f2072

  // f2074
  logic [0:0] f2074_wen;
  logic [31:0] f2074_wdata;
  logic [0:0] f2074_clk;
  logic [0:0] f2074_rst;
  logic [31:0] f2074_rdata;
  sr_buffer_32_1 f2074(.wen(f2074_wen), .wdata(f2074_wdata), .clk(f2074_clk), .rst(f2074_rst), .rdata(f2074_rdata));
  assign f2074_clk = clk;
  assign f2074_rst = rst;
  // Bindings to f2074

  // f2076
  logic [0:0] f2076_wen;
  logic [31:0] f2076_wdata;
  logic [0:0] f2076_clk;
  logic [0:0] f2076_rst;
  logic [31:0] f2076_rdata;
  sr_buffer_32_1 f2076(.wen(f2076_wen), .wdata(f2076_wdata), .clk(f2076_clk), .rst(f2076_rst), .rdata(f2076_rdata));
  assign f2076_clk = clk;
  assign f2076_rst = rst;
  // Bindings to f2076

  // f2078
  logic [0:0] f2078_wen;
  logic [31:0] f2078_wdata;
  logic [0:0] f2078_clk;
  logic [0:0] f2078_rst;
  logic [31:0] f2078_rdata;
  sr_buffer_32_1 f2078(.wen(f2078_wen), .wdata(f2078_wdata), .clk(f2078_clk), .rst(f2078_rst), .rdata(f2078_rdata));
  assign f2078_clk = clk;
  assign f2078_rst = rst;
  // Bindings to f2078

  // f2080
  logic [0:0] f2080_wen;
  logic [31:0] f2080_wdata;
  logic [0:0] f2080_clk;
  logic [0:0] f2080_rst;
  logic [31:0] f2080_rdata;
  sr_buffer_32_1 f2080(.wen(f2080_wen), .wdata(f2080_wdata), .clk(f2080_clk), .rst(f2080_rst), .rdata(f2080_rdata));
  assign f2080_clk = clk;
  assign f2080_rst = rst;
  // Bindings to f2080

  // f2082
  logic [0:0] f2082_wen;
  logic [31:0] f2082_wdata;
  logic [0:0] f2082_clk;
  logic [0:0] f2082_rst;
  logic [31:0] f2082_rdata;
  sr_buffer_32_1 f2082(.wen(f2082_wen), .wdata(f2082_wdata), .clk(f2082_clk), .rst(f2082_rst), .rdata(f2082_rdata));
  assign f2082_clk = clk;
  assign f2082_rst = rst;
  // Bindings to f2082

  // f2084
  logic [0:0] f2084_wen;
  logic [31:0] f2084_wdata;
  logic [0:0] f2084_clk;
  logic [0:0] f2084_rst;
  logic [31:0] f2084_rdata;
  sr_buffer_32_1 f2084(.wen(f2084_wen), .wdata(f2084_wdata), .clk(f2084_clk), .rst(f2084_rst), .rdata(f2084_rdata));
  assign f2084_clk = clk;
  assign f2084_rst = rst;
  // Bindings to f2084

  // f2086
  logic [0:0] f2086_wen;
  logic [31:0] f2086_wdata;
  logic [0:0] f2086_clk;
  logic [0:0] f2086_rst;
  logic [31:0] f2086_rdata;
  sr_buffer_32_1 f2086(.wen(f2086_wen), .wdata(f2086_wdata), .clk(f2086_clk), .rst(f2086_rst), .rdata(f2086_rdata));
  assign f2086_clk = clk;
  assign f2086_rst = rst;
  // Bindings to f2086

  // f2088
  logic [0:0] f2088_wen;
  logic [31:0] f2088_wdata;
  logic [0:0] f2088_clk;
  logic [0:0] f2088_rst;
  logic [31:0] f2088_rdata;
  sr_buffer_32_1 f2088(.wen(f2088_wen), .wdata(f2088_wdata), .clk(f2088_clk), .rst(f2088_rst), .rdata(f2088_rdata));
  assign f2088_clk = clk;
  assign f2088_rst = rst;
  // Bindings to f2088

  // f2090
  logic [0:0] f2090_wen;
  logic [31:0] f2090_wdata;
  logic [0:0] f2090_clk;
  logic [0:0] f2090_rst;
  logic [31:0] f2090_rdata;
  sr_buffer_32_1 f2090(.wen(f2090_wen), .wdata(f2090_wdata), .clk(f2090_clk), .rst(f2090_rst), .rdata(f2090_rdata));
  assign f2090_clk = clk;
  assign f2090_rst = rst;
  // Bindings to f2090

  // f2092
  logic [0:0] f2092_wen;
  logic [31:0] f2092_wdata;
  logic [0:0] f2092_clk;
  logic [0:0] f2092_rst;
  logic [31:0] f2092_rdata;
  sr_buffer_32_1 f2092(.wen(f2092_wen), .wdata(f2092_wdata), .clk(f2092_clk), .rst(f2092_rst), .rdata(f2092_rdata));
  assign f2092_clk = clk;
  assign f2092_rst = rst;
  // Bindings to f2092

  // f2094
  logic [0:0] f2094_wen;
  logic [31:0] f2094_wdata;
  logic [0:0] f2094_clk;
  logic [0:0] f2094_rst;
  logic [31:0] f2094_rdata;
  sr_buffer_32_1 f2094(.wen(f2094_wen), .wdata(f2094_wdata), .clk(f2094_clk), .rst(f2094_rst), .rdata(f2094_rdata));
  assign f2094_clk = clk;
  assign f2094_rst = rst;
  // Bindings to f2094

  // f2096
  logic [0:0] f2096_wen;
  logic [31:0] f2096_wdata;
  logic [0:0] f2096_clk;
  logic [0:0] f2096_rst;
  logic [31:0] f2096_rdata;
  sr_buffer_32_1 f2096(.wen(f2096_wen), .wdata(f2096_wdata), .clk(f2096_clk), .rst(f2096_rst), .rdata(f2096_rdata));
  assign f2096_clk = clk;
  assign f2096_rst = rst;
  // Bindings to f2096

  // f2098
  logic [0:0] f2098_wen;
  logic [31:0] f2098_wdata;
  logic [0:0] f2098_clk;
  logic [0:0] f2098_rst;
  logic [31:0] f2098_rdata;
  sr_buffer_32_1 f2098(.wen(f2098_wen), .wdata(f2098_wdata), .clk(f2098_clk), .rst(f2098_rst), .rdata(f2098_rdata));
  assign f2098_clk = clk;
  assign f2098_rst = rst;
  // Bindings to f2098

  // f2100
  logic [0:0] f2100_wen;
  logic [31:0] f2100_wdata;
  logic [0:0] f2100_clk;
  logic [0:0] f2100_rst;
  logic [31:0] f2100_rdata;
  sr_buffer_32_1 f2100(.wen(f2100_wen), .wdata(f2100_wdata), .clk(f2100_clk), .rst(f2100_rst), .rdata(f2100_rdata));
  assign f2100_clk = clk;
  assign f2100_rst = rst;
  // Bindings to f2100

  // f2102
  logic [0:0] f2102_wen;
  logic [31:0] f2102_wdata;
  logic [0:0] f2102_clk;
  logic [0:0] f2102_rst;
  logic [31:0] f2102_rdata;
  sr_buffer_32_1 f2102(.wen(f2102_wen), .wdata(f2102_wdata), .clk(f2102_clk), .rst(f2102_rst), .rdata(f2102_rdata));
  assign f2102_clk = clk;
  assign f2102_rst = rst;
  // Bindings to f2102

  // f2104
  logic [0:0] f2104_wen;
  logic [31:0] f2104_wdata;
  logic [0:0] f2104_clk;
  logic [0:0] f2104_rst;
  logic [31:0] f2104_rdata;
  sr_buffer_32_1 f2104(.wen(f2104_wen), .wdata(f2104_wdata), .clk(f2104_clk), .rst(f2104_rst), .rdata(f2104_rdata));
  assign f2104_clk = clk;
  assign f2104_rst = rst;
  // Bindings to f2104

  // f2106
  logic [0:0] f2106_wen;
  logic [31:0] f2106_wdata;
  logic [0:0] f2106_clk;
  logic [0:0] f2106_rst;
  logic [31:0] f2106_rdata;
  sr_buffer_32_1 f2106(.wen(f2106_wen), .wdata(f2106_wdata), .clk(f2106_clk), .rst(f2106_rst), .rdata(f2106_rdata));
  assign f2106_clk = clk;
  assign f2106_rst = rst;
  // Bindings to f2106

  // f2108
  logic [0:0] f2108_wen;
  logic [31:0] f2108_wdata;
  logic [0:0] f2108_clk;
  logic [0:0] f2108_rst;
  logic [31:0] f2108_rdata;
  sr_buffer_32_1 f2108(.wen(f2108_wen), .wdata(f2108_wdata), .clk(f2108_clk), .rst(f2108_rst), .rdata(f2108_rdata));
  assign f2108_clk = clk;
  assign f2108_rst = rst;
  // Bindings to f2108

  // f2110
  logic [0:0] f2110_wen;
  logic [31:0] f2110_wdata;
  logic [0:0] f2110_clk;
  logic [0:0] f2110_rst;
  logic [31:0] f2110_rdata;
  sr_buffer_32_1 f2110(.wen(f2110_wen), .wdata(f2110_wdata), .clk(f2110_clk), .rst(f2110_rst), .rdata(f2110_rdata));
  assign f2110_clk = clk;
  assign f2110_rst = rst;
  // Bindings to f2110

  // f2112
  logic [0:0] f2112_wen;
  logic [31:0] f2112_wdata;
  logic [0:0] f2112_clk;
  logic [0:0] f2112_rst;
  logic [31:0] f2112_rdata;
  sr_buffer_32_1 f2112(.wen(f2112_wen), .wdata(f2112_wdata), .clk(f2112_clk), .rst(f2112_rst), .rdata(f2112_rdata));
  assign f2112_clk = clk;
  assign f2112_rst = rst;
  // Bindings to f2112

  // f2114
  logic [0:0] f2114_wen;
  logic [31:0] f2114_wdata;
  logic [0:0] f2114_clk;
  logic [0:0] f2114_rst;
  logic [31:0] f2114_rdata;
  sr_buffer_32_1 f2114(.wen(f2114_wen), .wdata(f2114_wdata), .clk(f2114_clk), .rst(f2114_rst), .rdata(f2114_rdata));
  assign f2114_clk = clk;
  assign f2114_rst = rst;
  // Bindings to f2114

  // f2116
  logic [0:0] f2116_wen;
  logic [31:0] f2116_wdata;
  logic [0:0] f2116_clk;
  logic [0:0] f2116_rst;
  logic [31:0] f2116_rdata;
  sr_buffer_32_1 f2116(.wen(f2116_wen), .wdata(f2116_wdata), .clk(f2116_clk), .rst(f2116_rst), .rdata(f2116_rdata));
  assign f2116_clk = clk;
  assign f2116_rst = rst;
  // Bindings to f2116

  // f2118
  logic [0:0] f2118_wen;
  logic [31:0] f2118_wdata;
  logic [0:0] f2118_clk;
  logic [0:0] f2118_rst;
  logic [31:0] f2118_rdata;
  sr_buffer_32_1 f2118(.wen(f2118_wen), .wdata(f2118_wdata), .clk(f2118_clk), .rst(f2118_rst), .rdata(f2118_rdata));
  assign f2118_clk = clk;
  assign f2118_rst = rst;
  // Bindings to f2118

  // f2120
  logic [0:0] f2120_wen;
  logic [31:0] f2120_wdata;
  logic [0:0] f2120_clk;
  logic [0:0] f2120_rst;
  logic [31:0] f2120_rdata;
  sr_buffer_32_1 f2120(.wen(f2120_wen), .wdata(f2120_wdata), .clk(f2120_clk), .rst(f2120_rst), .rdata(f2120_rdata));
  assign f2120_clk = clk;
  assign f2120_rst = rst;
  // Bindings to f2120

  // f2122
  logic [0:0] f2122_wen;
  logic [31:0] f2122_wdata;
  logic [0:0] f2122_clk;
  logic [0:0] f2122_rst;
  logic [31:0] f2122_rdata;
  sr_buffer_32_1 f2122(.wen(f2122_wen), .wdata(f2122_wdata), .clk(f2122_clk), .rst(f2122_rst), .rdata(f2122_rdata));
  assign f2122_clk = clk;
  assign f2122_rst = rst;
  // Bindings to f2122

  // f2124
  logic [0:0] f2124_wen;
  logic [31:0] f2124_wdata;
  logic [0:0] f2124_clk;
  logic [0:0] f2124_rst;
  logic [31:0] f2124_rdata;
  sr_buffer_32_1 f2124(.wen(f2124_wen), .wdata(f2124_wdata), .clk(f2124_clk), .rst(f2124_rst), .rdata(f2124_rdata));
  assign f2124_clk = clk;
  assign f2124_rst = rst;
  // Bindings to f2124

  // f2126
  logic [0:0] f2126_wen;
  logic [31:0] f2126_wdata;
  logic [0:0] f2126_clk;
  logic [0:0] f2126_rst;
  logic [31:0] f2126_rdata;
  sr_buffer_32_1 f2126(.wen(f2126_wen), .wdata(f2126_wdata), .clk(f2126_clk), .rst(f2126_rst), .rdata(f2126_rdata));
  assign f2126_clk = clk;
  assign f2126_rst = rst;
  // Bindings to f2126

  // f2128
  logic [0:0] f2128_wen;
  logic [31:0] f2128_wdata;
  logic [0:0] f2128_clk;
  logic [0:0] f2128_rst;
  logic [31:0] f2128_rdata;
  sr_buffer_32_1 f2128(.wen(f2128_wen), .wdata(f2128_wdata), .clk(f2128_clk), .rst(f2128_rst), .rdata(f2128_rdata));
  assign f2128_clk = clk;
  assign f2128_rst = rst;
  // Bindings to f2128

  // f2130
  logic [0:0] f2130_wen;
  logic [31:0] f2130_wdata;
  logic [0:0] f2130_clk;
  logic [0:0] f2130_rst;
  logic [31:0] f2130_rdata;
  sr_buffer_32_1 f2130(.wen(f2130_wen), .wdata(f2130_wdata), .clk(f2130_clk), .rst(f2130_rst), .rdata(f2130_rdata));
  assign f2130_clk = clk;
  assign f2130_rst = rst;
  // Bindings to f2130

  // f2132
  logic [0:0] f2132_wen;
  logic [31:0] f2132_wdata;
  logic [0:0] f2132_clk;
  logic [0:0] f2132_rst;
  logic [31:0] f2132_rdata;
  sr_buffer_32_1 f2132(.wen(f2132_wen), .wdata(f2132_wdata), .clk(f2132_clk), .rst(f2132_rst), .rdata(f2132_rdata));
  assign f2132_clk = clk;
  assign f2132_rst = rst;
  // Bindings to f2132

  // f2134
  logic [0:0] f2134_wen;
  logic [31:0] f2134_wdata;
  logic [0:0] f2134_clk;
  logic [0:0] f2134_rst;
  logic [31:0] f2134_rdata;
  sr_buffer_32_1 f2134(.wen(f2134_wen), .wdata(f2134_wdata), .clk(f2134_clk), .rst(f2134_rst), .rdata(f2134_rdata));
  assign f2134_clk = clk;
  assign f2134_rst = rst;
  // Bindings to f2134

  // f2136
  logic [0:0] f2136_wen;
  logic [31:0] f2136_wdata;
  logic [0:0] f2136_clk;
  logic [0:0] f2136_rst;
  logic [31:0] f2136_rdata;
  sr_buffer_32_1 f2136(.wen(f2136_wen), .wdata(f2136_wdata), .clk(f2136_clk), .rst(f2136_rst), .rdata(f2136_rdata));
  assign f2136_clk = clk;
  assign f2136_rst = rst;
  // Bindings to f2136

  // f2138
  logic [0:0] f2138_wen;
  logic [31:0] f2138_wdata;
  logic [0:0] f2138_clk;
  logic [0:0] f2138_rst;
  logic [31:0] f2138_rdata;
  sr_buffer_32_1 f2138(.wen(f2138_wen), .wdata(f2138_wdata), .clk(f2138_clk), .rst(f2138_rst), .rdata(f2138_rdata));
  assign f2138_clk = clk;
  assign f2138_rst = rst;
  // Bindings to f2138

  // f2140
  logic [0:0] f2140_wen;
  logic [31:0] f2140_wdata;
  logic [0:0] f2140_clk;
  logic [0:0] f2140_rst;
  logic [31:0] f2140_rdata;
  sr_buffer_32_1 f2140(.wen(f2140_wen), .wdata(f2140_wdata), .clk(f2140_clk), .rst(f2140_rst), .rdata(f2140_rdata));
  assign f2140_clk = clk;
  assign f2140_rst = rst;
  // Bindings to f2140

  // f2142
  logic [0:0] f2142_wen;
  logic [31:0] f2142_wdata;
  logic [0:0] f2142_clk;
  logic [0:0] f2142_rst;
  logic [31:0] f2142_rdata;
  sr_buffer_32_1 f2142(.wen(f2142_wen), .wdata(f2142_wdata), .clk(f2142_clk), .rst(f2142_rst), .rdata(f2142_rdata));
  assign f2142_clk = clk;
  assign f2142_rst = rst;
  // Bindings to f2142

  // f2144
  logic [0:0] f2144_wen;
  logic [31:0] f2144_wdata;
  logic [0:0] f2144_clk;
  logic [0:0] f2144_rst;
  logic [31:0] f2144_rdata;
  sr_buffer_32_1 f2144(.wen(f2144_wen), .wdata(f2144_wdata), .clk(f2144_clk), .rst(f2144_rst), .rdata(f2144_rdata));
  assign f2144_clk = clk;
  assign f2144_rst = rst;
  // Bindings to f2144

  // f2146
  logic [0:0] f2146_wen;
  logic [31:0] f2146_wdata;
  logic [0:0] f2146_clk;
  logic [0:0] f2146_rst;
  logic [31:0] f2146_rdata;
  sr_buffer_32_1 f2146(.wen(f2146_wen), .wdata(f2146_wdata), .clk(f2146_clk), .rst(f2146_rst), .rdata(f2146_rdata));
  assign f2146_clk = clk;
  assign f2146_rst = rst;
  // Bindings to f2146

  // f2148
  logic [0:0] f2148_wen;
  logic [31:0] f2148_wdata;
  logic [0:0] f2148_clk;
  logic [0:0] f2148_rst;
  logic [31:0] f2148_rdata;
  sr_buffer_32_1 f2148(.wen(f2148_wen), .wdata(f2148_wdata), .clk(f2148_clk), .rst(f2148_rst), .rdata(f2148_rdata));
  assign f2148_clk = clk;
  assign f2148_rst = rst;
  // Bindings to f2148

  // f2150
  logic [0:0] f2150_wen;
  logic [31:0] f2150_wdata;
  logic [0:0] f2150_clk;
  logic [0:0] f2150_rst;
  logic [31:0] f2150_rdata;
  sr_buffer_32_1 f2150(.wen(f2150_wen), .wdata(f2150_wdata), .clk(f2150_clk), .rst(f2150_rst), .rdata(f2150_rdata));
  assign f2150_clk = clk;
  assign f2150_rst = rst;
  // Bindings to f2150

  // f2152
  logic [0:0] f2152_wen;
  logic [31:0] f2152_wdata;
  logic [0:0] f2152_clk;
  logic [0:0] f2152_rst;
  logic [31:0] f2152_rdata;
  sr_buffer_32_1 f2152(.wen(f2152_wen), .wdata(f2152_wdata), .clk(f2152_clk), .rst(f2152_rst), .rdata(f2152_rdata));
  assign f2152_clk = clk;
  assign f2152_rst = rst;
  // Bindings to f2152

  // f2154
  logic [0:0] f2154_wen;
  logic [31:0] f2154_wdata;
  logic [0:0] f2154_clk;
  logic [0:0] f2154_rst;
  logic [31:0] f2154_rdata;
  sr_buffer_32_1 f2154(.wen(f2154_wen), .wdata(f2154_wdata), .clk(f2154_clk), .rst(f2154_rst), .rdata(f2154_rdata));
  assign f2154_clk = clk;
  assign f2154_rst = rst;
  // Bindings to f2154

  // f2156
  logic [0:0] f2156_wen;
  logic [31:0] f2156_wdata;
  logic [0:0] f2156_clk;
  logic [0:0] f2156_rst;
  logic [31:0] f2156_rdata;
  sr_buffer_32_1 f2156(.wen(f2156_wen), .wdata(f2156_wdata), .clk(f2156_clk), .rst(f2156_rst), .rdata(f2156_rdata));
  assign f2156_clk = clk;
  assign f2156_rst = rst;
  // Bindings to f2156

  // f2158
  logic [0:0] f2158_wen;
  logic [31:0] f2158_wdata;
  logic [0:0] f2158_clk;
  logic [0:0] f2158_rst;
  logic [31:0] f2158_rdata;
  sr_buffer_32_1 f2158(.wen(f2158_wen), .wdata(f2158_wdata), .clk(f2158_clk), .rst(f2158_rst), .rdata(f2158_rdata));
  assign f2158_clk = clk;
  assign f2158_rst = rst;
  // Bindings to f2158

  // f2160
  logic [0:0] f2160_wen;
  logic [31:0] f2160_wdata;
  logic [0:0] f2160_clk;
  logic [0:0] f2160_rst;
  logic [31:0] f2160_rdata;
  sr_buffer_32_1 f2160(.wen(f2160_wen), .wdata(f2160_wdata), .clk(f2160_clk), .rst(f2160_rst), .rdata(f2160_rdata));
  assign f2160_clk = clk;
  assign f2160_rst = rst;
  // Bindings to f2160

  // f2162
  logic [0:0] f2162_wen;
  logic [31:0] f2162_wdata;
  logic [0:0] f2162_clk;
  logic [0:0] f2162_rst;
  logic [31:0] f2162_rdata;
  sr_buffer_32_1 f2162(.wen(f2162_wen), .wdata(f2162_wdata), .clk(f2162_clk), .rst(f2162_rst), .rdata(f2162_rdata));
  assign f2162_clk = clk;
  assign f2162_rst = rst;
  // Bindings to f2162

  // f2164
  logic [0:0] f2164_wen;
  logic [31:0] f2164_wdata;
  logic [0:0] f2164_clk;
  logic [0:0] f2164_rst;
  logic [31:0] f2164_rdata;
  sr_buffer_32_1 f2164(.wen(f2164_wen), .wdata(f2164_wdata), .clk(f2164_clk), .rst(f2164_rst), .rdata(f2164_rdata));
  assign f2164_clk = clk;
  assign f2164_rst = rst;
  // Bindings to f2164

  // f2166
  logic [0:0] f2166_wen;
  logic [31:0] f2166_wdata;
  logic [0:0] f2166_clk;
  logic [0:0] f2166_rst;
  logic [31:0] f2166_rdata;
  sr_buffer_32_1 f2166(.wen(f2166_wen), .wdata(f2166_wdata), .clk(f2166_clk), .rst(f2166_rst), .rdata(f2166_rdata));
  assign f2166_clk = clk;
  assign f2166_rst = rst;
  // Bindings to f2166

  // f2168
  logic [0:0] f2168_wen;
  logic [31:0] f2168_wdata;
  logic [0:0] f2168_clk;
  logic [0:0] f2168_rst;
  logic [31:0] f2168_rdata;
  sr_buffer_32_1 f2168(.wen(f2168_wen), .wdata(f2168_wdata), .clk(f2168_clk), .rst(f2168_rst), .rdata(f2168_rdata));
  assign f2168_clk = clk;
  assign f2168_rst = rst;
  // Bindings to f2168

  // f2170
  logic [0:0] f2170_wen;
  logic [31:0] f2170_wdata;
  logic [0:0] f2170_clk;
  logic [0:0] f2170_rst;
  logic [31:0] f2170_rdata;
  sr_buffer_32_1 f2170(.wen(f2170_wen), .wdata(f2170_wdata), .clk(f2170_clk), .rst(f2170_rst), .rdata(f2170_rdata));
  assign f2170_clk = clk;
  assign f2170_rst = rst;
  // Bindings to f2170

  // f2172
  logic [0:0] f2172_wen;
  logic [31:0] f2172_wdata;
  logic [0:0] f2172_clk;
  logic [0:0] f2172_rst;
  logic [31:0] f2172_rdata;
  sr_buffer_32_1 f2172(.wen(f2172_wen), .wdata(f2172_wdata), .clk(f2172_clk), .rst(f2172_rst), .rdata(f2172_rdata));
  assign f2172_clk = clk;
  assign f2172_rst = rst;
  // Bindings to f2172

  // f2174
  logic [0:0] f2174_wen;
  logic [31:0] f2174_wdata;
  logic [0:0] f2174_clk;
  logic [0:0] f2174_rst;
  logic [31:0] f2174_rdata;
  sr_buffer_32_1 f2174(.wen(f2174_wen), .wdata(f2174_wdata), .clk(f2174_clk), .rst(f2174_rst), .rdata(f2174_rdata));
  assign f2174_clk = clk;
  assign f2174_rst = rst;
  // Bindings to f2174

  // f2176
  logic [0:0] f2176_wen;
  logic [31:0] f2176_wdata;
  logic [0:0] f2176_clk;
  logic [0:0] f2176_rst;
  logic [31:0] f2176_rdata;
  sr_buffer_32_1 f2176(.wen(f2176_wen), .wdata(f2176_wdata), .clk(f2176_clk), .rst(f2176_rst), .rdata(f2176_rdata));
  assign f2176_clk = clk;
  assign f2176_rst = rst;
  // Bindings to f2176

  // f2178
  logic [0:0] f2178_wen;
  logic [31:0] f2178_wdata;
  logic [0:0] f2178_clk;
  logic [0:0] f2178_rst;
  logic [31:0] f2178_rdata;
  sr_buffer_32_1 f2178(.wen(f2178_wen), .wdata(f2178_wdata), .clk(f2178_clk), .rst(f2178_rst), .rdata(f2178_rdata));
  assign f2178_clk = clk;
  assign f2178_rst = rst;
  // Bindings to f2178

  // f2180
  logic [0:0] f2180_wen;
  logic [31:0] f2180_wdata;
  logic [0:0] f2180_clk;
  logic [0:0] f2180_rst;
  logic [31:0] f2180_rdata;
  sr_buffer_32_1 f2180(.wen(f2180_wen), .wdata(f2180_wdata), .clk(f2180_clk), .rst(f2180_rst), .rdata(f2180_rdata));
  assign f2180_clk = clk;
  assign f2180_rst = rst;
  // Bindings to f2180

  // f2182
  logic [0:0] f2182_wen;
  logic [31:0] f2182_wdata;
  logic [0:0] f2182_clk;
  logic [0:0] f2182_rst;
  logic [31:0] f2182_rdata;
  sr_buffer_32_1 f2182(.wen(f2182_wen), .wdata(f2182_wdata), .clk(f2182_clk), .rst(f2182_rst), .rdata(f2182_rdata));
  assign f2182_clk = clk;
  assign f2182_rst = rst;
  // Bindings to f2182

  // f2184
  logic [0:0] f2184_wen;
  logic [31:0] f2184_wdata;
  logic [0:0] f2184_clk;
  logic [0:0] f2184_rst;
  logic [31:0] f2184_rdata;
  sr_buffer_32_1 f2184(.wen(f2184_wen), .wdata(f2184_wdata), .clk(f2184_clk), .rst(f2184_rst), .rdata(f2184_rdata));
  assign f2184_clk = clk;
  assign f2184_rst = rst;
  // Bindings to f2184

  // f2186
  logic [0:0] f2186_wen;
  logic [31:0] f2186_wdata;
  logic [0:0] f2186_clk;
  logic [0:0] f2186_rst;
  logic [31:0] f2186_rdata;
  sr_buffer_32_1 f2186(.wen(f2186_wen), .wdata(f2186_wdata), .clk(f2186_clk), .rst(f2186_rst), .rdata(f2186_rdata));
  assign f2186_clk = clk;
  assign f2186_rst = rst;
  // Bindings to f2186

  // f2188
  logic [0:0] f2188_wen;
  logic [31:0] f2188_wdata;
  logic [0:0] f2188_clk;
  logic [0:0] f2188_rst;
  logic [31:0] f2188_rdata;
  sr_buffer_32_1 f2188(.wen(f2188_wen), .wdata(f2188_wdata), .clk(f2188_clk), .rst(f2188_rst), .rdata(f2188_rdata));
  assign f2188_clk = clk;
  assign f2188_rst = rst;
  // Bindings to f2188

  // f2190
  logic [0:0] f2190_wen;
  logic [31:0] f2190_wdata;
  logic [0:0] f2190_clk;
  logic [0:0] f2190_rst;
  logic [31:0] f2190_rdata;
  sr_buffer_32_1 f2190(.wen(f2190_wen), .wdata(f2190_wdata), .clk(f2190_clk), .rst(f2190_rst), .rdata(f2190_rdata));
  assign f2190_clk = clk;
  assign f2190_rst = rst;
  // Bindings to f2190

  // f2192
  logic [0:0] f2192_wen;
  logic [31:0] f2192_wdata;
  logic [0:0] f2192_clk;
  logic [0:0] f2192_rst;
  logic [31:0] f2192_rdata;
  sr_buffer_32_1 f2192(.wen(f2192_wen), .wdata(f2192_wdata), .clk(f2192_clk), .rst(f2192_rst), .rdata(f2192_rdata));
  assign f2192_clk = clk;
  assign f2192_rst = rst;
  // Bindings to f2192

  // f2194
  logic [0:0] f2194_wen;
  logic [31:0] f2194_wdata;
  logic [0:0] f2194_clk;
  logic [0:0] f2194_rst;
  logic [31:0] f2194_rdata;
  sr_buffer_32_1 f2194(.wen(f2194_wen), .wdata(f2194_wdata), .clk(f2194_clk), .rst(f2194_rst), .rdata(f2194_rdata));
  assign f2194_clk = clk;
  assign f2194_rst = rst;
  // Bindings to f2194

  // f2196
  logic [0:0] f2196_wen;
  logic [31:0] f2196_wdata;
  logic [0:0] f2196_clk;
  logic [0:0] f2196_rst;
  logic [31:0] f2196_rdata;
  sr_buffer_32_1 f2196(.wen(f2196_wen), .wdata(f2196_wdata), .clk(f2196_clk), .rst(f2196_rst), .rdata(f2196_rdata));
  assign f2196_clk = clk;
  assign f2196_rst = rst;
  // Bindings to f2196

  // f2198
  logic [0:0] f2198_wen;
  logic [31:0] f2198_wdata;
  logic [0:0] f2198_clk;
  logic [0:0] f2198_rst;
  logic [31:0] f2198_rdata;
  sr_buffer_32_1 f2198(.wen(f2198_wen), .wdata(f2198_wdata), .clk(f2198_clk), .rst(f2198_rst), .rdata(f2198_rdata));
  assign f2198_clk = clk;
  assign f2198_rst = rst;
  // Bindings to f2198

  // f2200
  logic [0:0] f2200_wen;
  logic [31:0] f2200_wdata;
  logic [0:0] f2200_clk;
  logic [0:0] f2200_rst;
  logic [31:0] f2200_rdata;
  sr_buffer_32_1 f2200(.wen(f2200_wen), .wdata(f2200_wdata), .clk(f2200_clk), .rst(f2200_rst), .rdata(f2200_rdata));
  assign f2200_clk = clk;
  assign f2200_rst = rst;
  // Bindings to f2200

  // f2202
  logic [0:0] f2202_wen;
  logic [31:0] f2202_wdata;
  logic [0:0] f2202_clk;
  logic [0:0] f2202_rst;
  logic [31:0] f2202_rdata;
  sr_buffer_32_1 f2202(.wen(f2202_wen), .wdata(f2202_wdata), .clk(f2202_clk), .rst(f2202_rst), .rdata(f2202_rdata));
  assign f2202_clk = clk;
  assign f2202_rst = rst;
  // Bindings to f2202

  // f2204
  logic [0:0] f2204_wen;
  logic [31:0] f2204_wdata;
  logic [0:0] f2204_clk;
  logic [0:0] f2204_rst;
  logic [31:0] f2204_rdata;
  sr_buffer_32_1 f2204(.wen(f2204_wen), .wdata(f2204_wdata), .clk(f2204_clk), .rst(f2204_rst), .rdata(f2204_rdata));
  assign f2204_clk = clk;
  assign f2204_rst = rst;
  // Bindings to f2204

  // f2206
  logic [0:0] f2206_wen;
  logic [31:0] f2206_wdata;
  logic [0:0] f2206_clk;
  logic [0:0] f2206_rst;
  logic [31:0] f2206_rdata;
  sr_buffer_32_1 f2206(.wen(f2206_wen), .wdata(f2206_wdata), .clk(f2206_clk), .rst(f2206_rst), .rdata(f2206_rdata));
  assign f2206_clk = clk;
  assign f2206_rst = rst;
  // Bindings to f2206

  // f2208
  logic [0:0] f2208_wen;
  logic [31:0] f2208_wdata;
  logic [0:0] f2208_clk;
  logic [0:0] f2208_rst;
  logic [31:0] f2208_rdata;
  sr_buffer_32_1 f2208(.wen(f2208_wen), .wdata(f2208_wdata), .clk(f2208_clk), .rst(f2208_rst), .rdata(f2208_rdata));
  assign f2208_clk = clk;
  assign f2208_rst = rst;
  // Bindings to f2208

  // f2210
  logic [0:0] f2210_wen;
  logic [31:0] f2210_wdata;
  logic [0:0] f2210_clk;
  logic [0:0] f2210_rst;
  logic [31:0] f2210_rdata;
  sr_buffer_32_1 f2210(.wen(f2210_wen), .wdata(f2210_wdata), .clk(f2210_clk), .rst(f2210_rst), .rdata(f2210_rdata));
  assign f2210_clk = clk;
  assign f2210_rst = rst;
  // Bindings to f2210

  // f2212
  logic [0:0] f2212_wen;
  logic [31:0] f2212_wdata;
  logic [0:0] f2212_clk;
  logic [0:0] f2212_rst;
  logic [31:0] f2212_rdata;
  sr_buffer_32_1 f2212(.wen(f2212_wen), .wdata(f2212_wdata), .clk(f2212_clk), .rst(f2212_rst), .rdata(f2212_rdata));
  assign f2212_clk = clk;
  assign f2212_rst = rst;
  // Bindings to f2212

  // f2214
  logic [0:0] f2214_wen;
  logic [31:0] f2214_wdata;
  logic [0:0] f2214_clk;
  logic [0:0] f2214_rst;
  logic [31:0] f2214_rdata;
  sr_buffer_32_1 f2214(.wen(f2214_wen), .wdata(f2214_wdata), .clk(f2214_clk), .rst(f2214_rst), .rdata(f2214_rdata));
  assign f2214_clk = clk;
  assign f2214_rst = rst;
  // Bindings to f2214

  // f2216
  logic [0:0] f2216_wen;
  logic [31:0] f2216_wdata;
  logic [0:0] f2216_clk;
  logic [0:0] f2216_rst;
  logic [31:0] f2216_rdata;
  sr_buffer_32_1 f2216(.wen(f2216_wen), .wdata(f2216_wdata), .clk(f2216_clk), .rst(f2216_rst), .rdata(f2216_rdata));
  assign f2216_clk = clk;
  assign f2216_rst = rst;
  // Bindings to f2216

  // f2218
  logic [0:0] f2218_wen;
  logic [31:0] f2218_wdata;
  logic [0:0] f2218_clk;
  logic [0:0] f2218_rst;
  logic [31:0] f2218_rdata;
  sr_buffer_32_1 f2218(.wen(f2218_wen), .wdata(f2218_wdata), .clk(f2218_clk), .rst(f2218_rst), .rdata(f2218_rdata));
  assign f2218_clk = clk;
  assign f2218_rst = rst;
  // Bindings to f2218

  // f2220
  logic [0:0] f2220_wen;
  logic [31:0] f2220_wdata;
  logic [0:0] f2220_clk;
  logic [0:0] f2220_rst;
  logic [31:0] f2220_rdata;
  sr_buffer_32_1 f2220(.wen(f2220_wen), .wdata(f2220_wdata), .clk(f2220_clk), .rst(f2220_rst), .rdata(f2220_rdata));
  assign f2220_clk = clk;
  assign f2220_rst = rst;
  // Bindings to f2220

  // f2222
  logic [0:0] f2222_wen;
  logic [31:0] f2222_wdata;
  logic [0:0] f2222_clk;
  logic [0:0] f2222_rst;
  logic [31:0] f2222_rdata;
  sr_buffer_32_1 f2222(.wen(f2222_wen), .wdata(f2222_wdata), .clk(f2222_clk), .rst(f2222_rst), .rdata(f2222_rdata));
  assign f2222_clk = clk;
  assign f2222_rst = rst;
  // Bindings to f2222

  // f2224
  logic [0:0] f2224_wen;
  logic [31:0] f2224_wdata;
  logic [0:0] f2224_clk;
  logic [0:0] f2224_rst;
  logic [31:0] f2224_rdata;
  sr_buffer_32_1 f2224(.wen(f2224_wen), .wdata(f2224_wdata), .clk(f2224_clk), .rst(f2224_rst), .rdata(f2224_rdata));
  assign f2224_clk = clk;
  assign f2224_rst = rst;
  // Bindings to f2224

  // f2226
  logic [0:0] f2226_wen;
  logic [31:0] f2226_wdata;
  logic [0:0] f2226_clk;
  logic [0:0] f2226_rst;
  logic [31:0] f2226_rdata;
  sr_buffer_32_1 f2226(.wen(f2226_wen), .wdata(f2226_wdata), .clk(f2226_clk), .rst(f2226_rst), .rdata(f2226_rdata));
  assign f2226_clk = clk;
  assign f2226_rst = rst;
  // Bindings to f2226

  // f2228
  logic [0:0] f2228_wen;
  logic [31:0] f2228_wdata;
  logic [0:0] f2228_clk;
  logic [0:0] f2228_rst;
  logic [31:0] f2228_rdata;
  sr_buffer_32_1 f2228(.wen(f2228_wen), .wdata(f2228_wdata), .clk(f2228_clk), .rst(f2228_rst), .rdata(f2228_rdata));
  assign f2228_clk = clk;
  assign f2228_rst = rst;
  // Bindings to f2228

  // f2230
  logic [0:0] f2230_wen;
  logic [31:0] f2230_wdata;
  logic [0:0] f2230_clk;
  logic [0:0] f2230_rst;
  logic [31:0] f2230_rdata;
  sr_buffer_32_1 f2230(.wen(f2230_wen), .wdata(f2230_wdata), .clk(f2230_clk), .rst(f2230_rst), .rdata(f2230_rdata));
  assign f2230_clk = clk;
  assign f2230_rst = rst;
  // Bindings to f2230

  // f2232
  logic [0:0] f2232_wen;
  logic [31:0] f2232_wdata;
  logic [0:0] f2232_clk;
  logic [0:0] f2232_rst;
  logic [31:0] f2232_rdata;
  sr_buffer_32_1 f2232(.wen(f2232_wen), .wdata(f2232_wdata), .clk(f2232_clk), .rst(f2232_rst), .rdata(f2232_rdata));
  assign f2232_clk = clk;
  assign f2232_rst = rst;
  // Bindings to f2232

  // f2234
  logic [0:0] f2234_wen;
  logic [31:0] f2234_wdata;
  logic [0:0] f2234_clk;
  logic [0:0] f2234_rst;
  logic [31:0] f2234_rdata;
  sr_buffer_32_1 f2234(.wen(f2234_wen), .wdata(f2234_wdata), .clk(f2234_clk), .rst(f2234_rst), .rdata(f2234_rdata));
  assign f2234_clk = clk;
  assign f2234_rst = rst;
  // Bindings to f2234

  // f2236
  logic [0:0] f2236_wen;
  logic [31:0] f2236_wdata;
  logic [0:0] f2236_clk;
  logic [0:0] f2236_rst;
  logic [31:0] f2236_rdata;
  sr_buffer_32_1 f2236(.wen(f2236_wen), .wdata(f2236_wdata), .clk(f2236_clk), .rst(f2236_rst), .rdata(f2236_rdata));
  assign f2236_clk = clk;
  assign f2236_rst = rst;
  // Bindings to f2236

  // f2238
  logic [0:0] f2238_wen;
  logic [31:0] f2238_wdata;
  logic [0:0] f2238_clk;
  logic [0:0] f2238_rst;
  logic [31:0] f2238_rdata;
  sr_buffer_32_1 f2238(.wen(f2238_wen), .wdata(f2238_wdata), .clk(f2238_clk), .rst(f2238_rst), .rdata(f2238_rdata));
  assign f2238_clk = clk;
  assign f2238_rst = rst;
  // Bindings to f2238

  // f2240
  logic [0:0] f2240_wen;
  logic [31:0] f2240_wdata;
  logic [0:0] f2240_clk;
  logic [0:0] f2240_rst;
  logic [31:0] f2240_rdata;
  sr_buffer_32_1 f2240(.wen(f2240_wen), .wdata(f2240_wdata), .clk(f2240_clk), .rst(f2240_rst), .rdata(f2240_rdata));
  assign f2240_clk = clk;
  assign f2240_rst = rst;
  // Bindings to f2240

  // f2242
  logic [0:0] f2242_wen;
  logic [31:0] f2242_wdata;
  logic [0:0] f2242_clk;
  logic [0:0] f2242_rst;
  logic [31:0] f2242_rdata;
  sr_buffer_32_1 f2242(.wen(f2242_wen), .wdata(f2242_wdata), .clk(f2242_clk), .rst(f2242_rst), .rdata(f2242_rdata));
  assign f2242_clk = clk;
  assign f2242_rst = rst;
  // Bindings to f2242

  // f2244
  logic [0:0] f2244_wen;
  logic [31:0] f2244_wdata;
  logic [0:0] f2244_clk;
  logic [0:0] f2244_rst;
  logic [31:0] f2244_rdata;
  sr_buffer_32_1 f2244(.wen(f2244_wen), .wdata(f2244_wdata), .clk(f2244_clk), .rst(f2244_rst), .rdata(f2244_rdata));
  assign f2244_clk = clk;
  assign f2244_rst = rst;
  // Bindings to f2244

  // f2246
  logic [0:0] f2246_wen;
  logic [31:0] f2246_wdata;
  logic [0:0] f2246_clk;
  logic [0:0] f2246_rst;
  logic [31:0] f2246_rdata;
  sr_buffer_32_1 f2246(.wen(f2246_wen), .wdata(f2246_wdata), .clk(f2246_clk), .rst(f2246_rst), .rdata(f2246_rdata));
  assign f2246_clk = clk;
  assign f2246_rst = rst;
  // Bindings to f2246

  // f2248
  logic [0:0] f2248_wen;
  logic [31:0] f2248_wdata;
  logic [0:0] f2248_clk;
  logic [0:0] f2248_rst;
  logic [31:0] f2248_rdata;
  sr_buffer_32_1 f2248(.wen(f2248_wen), .wdata(f2248_wdata), .clk(f2248_clk), .rst(f2248_rst), .rdata(f2248_rdata));
  assign f2248_clk = clk;
  assign f2248_rst = rst;
  // Bindings to f2248

  // f2250
  logic [0:0] f2250_wen;
  logic [31:0] f2250_wdata;
  logic [0:0] f2250_clk;
  logic [0:0] f2250_rst;
  logic [31:0] f2250_rdata;
  sr_buffer_32_1 f2250(.wen(f2250_wen), .wdata(f2250_wdata), .clk(f2250_clk), .rst(f2250_rst), .rdata(f2250_rdata));
  assign f2250_clk = clk;
  assign f2250_rst = rst;
  // Bindings to f2250

  // f2252
  logic [0:0] f2252_wen;
  logic [31:0] f2252_wdata;
  logic [0:0] f2252_clk;
  logic [0:0] f2252_rst;
  logic [31:0] f2252_rdata;
  sr_buffer_32_1 f2252(.wen(f2252_wen), .wdata(f2252_wdata), .clk(f2252_clk), .rst(f2252_rst), .rdata(f2252_rdata));
  assign f2252_clk = clk;
  assign f2252_rst = rst;
  // Bindings to f2252

  // f2254
  logic [0:0] f2254_wen;
  logic [31:0] f2254_wdata;
  logic [0:0] f2254_clk;
  logic [0:0] f2254_rst;
  logic [31:0] f2254_rdata;
  sr_buffer_32_1 f2254(.wen(f2254_wen), .wdata(f2254_wdata), .clk(f2254_clk), .rst(f2254_rst), .rdata(f2254_rdata));
  assign f2254_clk = clk;
  assign f2254_rst = rst;
  // Bindings to f2254

  // f2256
  logic [0:0] f2256_wen;
  logic [31:0] f2256_wdata;
  logic [0:0] f2256_clk;
  logic [0:0] f2256_rst;
  logic [31:0] f2256_rdata;
  sr_buffer_32_1 f2256(.wen(f2256_wen), .wdata(f2256_wdata), .clk(f2256_clk), .rst(f2256_rst), .rdata(f2256_rdata));
  assign f2256_clk = clk;
  assign f2256_rst = rst;
  // Bindings to f2256

  // f2258
  logic [0:0] f2258_wen;
  logic [31:0] f2258_wdata;
  logic [0:0] f2258_clk;
  logic [0:0] f2258_rst;
  logic [31:0] f2258_rdata;
  sr_buffer_32_1 f2258(.wen(f2258_wen), .wdata(f2258_wdata), .clk(f2258_clk), .rst(f2258_rst), .rdata(f2258_rdata));
  assign f2258_clk = clk;
  assign f2258_rst = rst;
  // Bindings to f2258

  // f2260
  logic [0:0] f2260_wen;
  logic [31:0] f2260_wdata;
  logic [0:0] f2260_clk;
  logic [0:0] f2260_rst;
  logic [31:0] f2260_rdata;
  sr_buffer_32_1 f2260(.wen(f2260_wen), .wdata(f2260_wdata), .clk(f2260_clk), .rst(f2260_rst), .rdata(f2260_rdata));
  assign f2260_clk = clk;
  assign f2260_rst = rst;
  // Bindings to f2260

  // f2262
  logic [0:0] f2262_wen;
  logic [31:0] f2262_wdata;
  logic [0:0] f2262_clk;
  logic [0:0] f2262_rst;
  logic [31:0] f2262_rdata;
  sr_buffer_32_1 f2262(.wen(f2262_wen), .wdata(f2262_wdata), .clk(f2262_clk), .rst(f2262_rst), .rdata(f2262_rdata));
  assign f2262_clk = clk;
  assign f2262_rst = rst;
  // Bindings to f2262

  // f2264
  logic [0:0] f2264_wen;
  logic [31:0] f2264_wdata;
  logic [0:0] f2264_clk;
  logic [0:0] f2264_rst;
  logic [31:0] f2264_rdata;
  sr_buffer_32_1 f2264(.wen(f2264_wen), .wdata(f2264_wdata), .clk(f2264_clk), .rst(f2264_rst), .rdata(f2264_rdata));
  assign f2264_clk = clk;
  assign f2264_rst = rst;
  // Bindings to f2264

  // f2266
  logic [0:0] f2266_wen;
  logic [31:0] f2266_wdata;
  logic [0:0] f2266_clk;
  logic [0:0] f2266_rst;
  logic [31:0] f2266_rdata;
  sr_buffer_32_1 f2266(.wen(f2266_wen), .wdata(f2266_wdata), .clk(f2266_clk), .rst(f2266_rst), .rdata(f2266_rdata));
  assign f2266_clk = clk;
  assign f2266_rst = rst;
  // Bindings to f2266

  // f2268
  logic [0:0] f2268_wen;
  logic [31:0] f2268_wdata;
  logic [0:0] f2268_clk;
  logic [0:0] f2268_rst;
  logic [31:0] f2268_rdata;
  sr_buffer_32_1 f2268(.wen(f2268_wen), .wdata(f2268_wdata), .clk(f2268_clk), .rst(f2268_rst), .rdata(f2268_rdata));
  assign f2268_clk = clk;
  assign f2268_rst = rst;
  // Bindings to f2268

  // f2270
  logic [0:0] f2270_wen;
  logic [31:0] f2270_wdata;
  logic [0:0] f2270_clk;
  logic [0:0] f2270_rst;
  logic [31:0] f2270_rdata;
  sr_buffer_32_1 f2270(.wen(f2270_wen), .wdata(f2270_wdata), .clk(f2270_clk), .rst(f2270_rst), .rdata(f2270_rdata));
  assign f2270_clk = clk;
  assign f2270_rst = rst;
  // Bindings to f2270

  // f2272
  logic [0:0] f2272_wen;
  logic [31:0] f2272_wdata;
  logic [0:0] f2272_clk;
  logic [0:0] f2272_rst;
  logic [31:0] f2272_rdata;
  sr_buffer_32_1 f2272(.wen(f2272_wen), .wdata(f2272_wdata), .clk(f2272_clk), .rst(f2272_rst), .rdata(f2272_rdata));
  assign f2272_clk = clk;
  assign f2272_rst = rst;
  // Bindings to f2272

  // f2274
  logic [0:0] f2274_wen;
  logic [31:0] f2274_wdata;
  logic [0:0] f2274_clk;
  logic [0:0] f2274_rst;
  logic [31:0] f2274_rdata;
  sr_buffer_32_1 f2274(.wen(f2274_wen), .wdata(f2274_wdata), .clk(f2274_clk), .rst(f2274_rst), .rdata(f2274_rdata));
  assign f2274_clk = clk;
  assign f2274_rst = rst;
  // Bindings to f2274

  // f2276
  logic [0:0] f2276_wen;
  logic [31:0] f2276_wdata;
  logic [0:0] f2276_clk;
  logic [0:0] f2276_rst;
  logic [31:0] f2276_rdata;
  sr_buffer_32_1 f2276(.wen(f2276_wen), .wdata(f2276_wdata), .clk(f2276_clk), .rst(f2276_rst), .rdata(f2276_rdata));
  assign f2276_clk = clk;
  assign f2276_rst = rst;
  // Bindings to f2276

  // f2278
  logic [0:0] f2278_wen;
  logic [31:0] f2278_wdata;
  logic [0:0] f2278_clk;
  logic [0:0] f2278_rst;
  logic [31:0] f2278_rdata;
  sr_buffer_32_1 f2278(.wen(f2278_wen), .wdata(f2278_wdata), .clk(f2278_clk), .rst(f2278_rst), .rdata(f2278_rdata));
  assign f2278_clk = clk;
  assign f2278_rst = rst;
  // Bindings to f2278

  // f2280
  logic [0:0] f2280_wen;
  logic [31:0] f2280_wdata;
  logic [0:0] f2280_clk;
  logic [0:0] f2280_rst;
  logic [31:0] f2280_rdata;
  sr_buffer_32_1 f2280(.wen(f2280_wen), .wdata(f2280_wdata), .clk(f2280_clk), .rst(f2280_rst), .rdata(f2280_rdata));
  assign f2280_clk = clk;
  assign f2280_rst = rst;
  // Bindings to f2280

  // f2282
  logic [0:0] f2282_wen;
  logic [31:0] f2282_wdata;
  logic [0:0] f2282_clk;
  logic [0:0] f2282_rst;
  logic [31:0] f2282_rdata;
  sr_buffer_32_1 f2282(.wen(f2282_wen), .wdata(f2282_wdata), .clk(f2282_clk), .rst(f2282_rst), .rdata(f2282_rdata));
  assign f2282_clk = clk;
  assign f2282_rst = rst;
  // Bindings to f2282

  // f2284
  logic [0:0] f2284_wen;
  logic [31:0] f2284_wdata;
  logic [0:0] f2284_clk;
  logic [0:0] f2284_rst;
  logic [31:0] f2284_rdata;
  sr_buffer_32_1 f2284(.wen(f2284_wen), .wdata(f2284_wdata), .clk(f2284_clk), .rst(f2284_rst), .rdata(f2284_rdata));
  assign f2284_clk = clk;
  assign f2284_rst = rst;
  // Bindings to f2284

  // f2286
  logic [0:0] f2286_wen;
  logic [31:0] f2286_wdata;
  logic [0:0] f2286_clk;
  logic [0:0] f2286_rst;
  logic [31:0] f2286_rdata;
  sr_buffer_32_1 f2286(.wen(f2286_wen), .wdata(f2286_wdata), .clk(f2286_clk), .rst(f2286_rst), .rdata(f2286_rdata));
  assign f2286_clk = clk;
  assign f2286_rst = rst;
  // Bindings to f2286

  // f2288
  logic [0:0] f2288_wen;
  logic [31:0] f2288_wdata;
  logic [0:0] f2288_clk;
  logic [0:0] f2288_rst;
  logic [31:0] f2288_rdata;
  sr_buffer_32_1 f2288(.wen(f2288_wen), .wdata(f2288_wdata), .clk(f2288_clk), .rst(f2288_rst), .rdata(f2288_rdata));
  assign f2288_clk = clk;
  assign f2288_rst = rst;
  // Bindings to f2288

  // f2290
  logic [0:0] f2290_wen;
  logic [31:0] f2290_wdata;
  logic [0:0] f2290_clk;
  logic [0:0] f2290_rst;
  logic [31:0] f2290_rdata;
  sr_buffer_32_1 f2290(.wen(f2290_wen), .wdata(f2290_wdata), .clk(f2290_clk), .rst(f2290_rst), .rdata(f2290_rdata));
  assign f2290_clk = clk;
  assign f2290_rst = rst;
  // Bindings to f2290

  // f2292
  logic [0:0] f2292_wen;
  logic [31:0] f2292_wdata;
  logic [0:0] f2292_clk;
  logic [0:0] f2292_rst;
  logic [31:0] f2292_rdata;
  sr_buffer_32_1 f2292(.wen(f2292_wen), .wdata(f2292_wdata), .clk(f2292_clk), .rst(f2292_rst), .rdata(f2292_rdata));
  assign f2292_clk = clk;
  assign f2292_rst = rst;
  // Bindings to f2292

  // f2294
  logic [0:0] f2294_wen;
  logic [31:0] f2294_wdata;
  logic [0:0] f2294_clk;
  logic [0:0] f2294_rst;
  logic [31:0] f2294_rdata;
  sr_buffer_32_1 f2294(.wen(f2294_wen), .wdata(f2294_wdata), .clk(f2294_clk), .rst(f2294_rst), .rdata(f2294_rdata));
  assign f2294_clk = clk;
  assign f2294_rst = rst;
  // Bindings to f2294

  // f2296
  logic [0:0] f2296_wen;
  logic [31:0] f2296_wdata;
  logic [0:0] f2296_clk;
  logic [0:0] f2296_rst;
  logic [31:0] f2296_rdata;
  sr_buffer_32_1 f2296(.wen(f2296_wen), .wdata(f2296_wdata), .clk(f2296_clk), .rst(f2296_rst), .rdata(f2296_rdata));
  assign f2296_clk = clk;
  assign f2296_rst = rst;
  // Bindings to f2296

  // f2298
  logic [0:0] f2298_wen;
  logic [31:0] f2298_wdata;
  logic [0:0] f2298_clk;
  logic [0:0] f2298_rst;
  logic [31:0] f2298_rdata;
  sr_buffer_32_1 f2298(.wen(f2298_wen), .wdata(f2298_wdata), .clk(f2298_clk), .rst(f2298_rst), .rdata(f2298_rdata));
  assign f2298_clk = clk;
  assign f2298_rst = rst;
  // Bindings to f2298

  // f2300
  logic [0:0] f2300_wen;
  logic [31:0] f2300_wdata;
  logic [0:0] f2300_clk;
  logic [0:0] f2300_rst;
  logic [31:0] f2300_rdata;
  sr_buffer_32_1 f2300(.wen(f2300_wen), .wdata(f2300_wdata), .clk(f2300_clk), .rst(f2300_rst), .rdata(f2300_rdata));
  assign f2300_clk = clk;
  assign f2300_rst = rst;
  // Bindings to f2300

  // f2302
  logic [0:0] f2302_wen;
  logic [31:0] f2302_wdata;
  logic [0:0] f2302_clk;
  logic [0:0] f2302_rst;
  logic [31:0] f2302_rdata;
  sr_buffer_32_1 f2302(.wen(f2302_wen), .wdata(f2302_wdata), .clk(f2302_clk), .rst(f2302_rst), .rdata(f2302_rdata));
  assign f2302_clk = clk;
  assign f2302_rst = rst;
  // Bindings to f2302

  // f2304
  logic [0:0] f2304_wen;
  logic [31:0] f2304_wdata;
  logic [0:0] f2304_clk;
  logic [0:0] f2304_rst;
  logic [31:0] f2304_rdata;
  sr_buffer_32_1 f2304(.wen(f2304_wen), .wdata(f2304_wdata), .clk(f2304_clk), .rst(f2304_rst), .rdata(f2304_rdata));
  assign f2304_clk = clk;
  assign f2304_rst = rst;
  // Bindings to f2304

  // f2306
  logic [0:0] f2306_wen;
  logic [31:0] f2306_wdata;
  logic [0:0] f2306_clk;
  logic [0:0] f2306_rst;
  logic [31:0] f2306_rdata;
  sr_buffer_32_1 f2306(.wen(f2306_wen), .wdata(f2306_wdata), .clk(f2306_clk), .rst(f2306_rst), .rdata(f2306_rdata));
  assign f2306_clk = clk;
  assign f2306_rst = rst;
  // Bindings to f2306

  // f2308
  logic [0:0] f2308_wen;
  logic [31:0] f2308_wdata;
  logic [0:0] f2308_clk;
  logic [0:0] f2308_rst;
  logic [31:0] f2308_rdata;
  sr_buffer_32_1 f2308(.wen(f2308_wen), .wdata(f2308_wdata), .clk(f2308_clk), .rst(f2308_rst), .rdata(f2308_rdata));
  assign f2308_clk = clk;
  assign f2308_rst = rst;
  // Bindings to f2308

  // f2310
  logic [0:0] f2310_wen;
  logic [31:0] f2310_wdata;
  logic [0:0] f2310_clk;
  logic [0:0] f2310_rst;
  logic [31:0] f2310_rdata;
  sr_buffer_32_1 f2310(.wen(f2310_wen), .wdata(f2310_wdata), .clk(f2310_clk), .rst(f2310_rst), .rdata(f2310_rdata));
  assign f2310_clk = clk;
  assign f2310_rst = rst;
  // Bindings to f2310

  // f2312
  logic [0:0] f2312_wen;
  logic [31:0] f2312_wdata;
  logic [0:0] f2312_clk;
  logic [0:0] f2312_rst;
  logic [31:0] f2312_rdata;
  sr_buffer_32_1 f2312(.wen(f2312_wen), .wdata(f2312_wdata), .clk(f2312_clk), .rst(f2312_rst), .rdata(f2312_rdata));
  assign f2312_clk = clk;
  assign f2312_rst = rst;
  // Bindings to f2312

  // f2314
  logic [0:0] f2314_wen;
  logic [31:0] f2314_wdata;
  logic [0:0] f2314_clk;
  logic [0:0] f2314_rst;
  logic [31:0] f2314_rdata;
  sr_buffer_32_1 f2314(.wen(f2314_wen), .wdata(f2314_wdata), .clk(f2314_clk), .rst(f2314_rst), .rdata(f2314_rdata));
  assign f2314_clk = clk;
  assign f2314_rst = rst;
  // Bindings to f2314

  // f2316
  logic [0:0] f2316_wen;
  logic [31:0] f2316_wdata;
  logic [0:0] f2316_clk;
  logic [0:0] f2316_rst;
  logic [31:0] f2316_rdata;
  sr_buffer_32_1 f2316(.wen(f2316_wen), .wdata(f2316_wdata), .clk(f2316_clk), .rst(f2316_rst), .rdata(f2316_rdata));
  assign f2316_clk = clk;
  assign f2316_rst = rst;
  // Bindings to f2316

  // f2318
  logic [0:0] f2318_wen;
  logic [31:0] f2318_wdata;
  logic [0:0] f2318_clk;
  logic [0:0] f2318_rst;
  logic [31:0] f2318_rdata;
  sr_buffer_32_1 f2318(.wen(f2318_wen), .wdata(f2318_wdata), .clk(f2318_clk), .rst(f2318_rst), .rdata(f2318_rdata));
  assign f2318_clk = clk;
  assign f2318_rst = rst;
  // Bindings to f2318

  // f2320
  logic [0:0] f2320_wen;
  logic [31:0] f2320_wdata;
  logic [0:0] f2320_clk;
  logic [0:0] f2320_rst;
  logic [31:0] f2320_rdata;
  sr_buffer_32_1 f2320(.wen(f2320_wen), .wdata(f2320_wdata), .clk(f2320_clk), .rst(f2320_rst), .rdata(f2320_rdata));
  assign f2320_clk = clk;
  assign f2320_rst = rst;
  // Bindings to f2320

  // f2322
  logic [0:0] f2322_wen;
  logic [31:0] f2322_wdata;
  logic [0:0] f2322_clk;
  logic [0:0] f2322_rst;
  logic [31:0] f2322_rdata;
  sr_buffer_32_1 f2322(.wen(f2322_wen), .wdata(f2322_wdata), .clk(f2322_clk), .rst(f2322_rst), .rdata(f2322_rdata));
  assign f2322_clk = clk;
  assign f2322_rst = rst;
  // Bindings to f2322

  // f2324
  logic [0:0] f2324_wen;
  logic [31:0] f2324_wdata;
  logic [0:0] f2324_clk;
  logic [0:0] f2324_rst;
  logic [31:0] f2324_rdata;
  sr_buffer_32_1 f2324(.wen(f2324_wen), .wdata(f2324_wdata), .clk(f2324_clk), .rst(f2324_rst), .rdata(f2324_rdata));
  assign f2324_clk = clk;
  assign f2324_rst = rst;
  // Bindings to f2324

  // f2326
  logic [0:0] f2326_wen;
  logic [31:0] f2326_wdata;
  logic [0:0] f2326_clk;
  logic [0:0] f2326_rst;
  logic [31:0] f2326_rdata;
  sr_buffer_32_1 f2326(.wen(f2326_wen), .wdata(f2326_wdata), .clk(f2326_clk), .rst(f2326_rst), .rdata(f2326_rdata));
  assign f2326_clk = clk;
  assign f2326_rst = rst;
  // Bindings to f2326

  // f2328
  logic [0:0] f2328_wen;
  logic [31:0] f2328_wdata;
  logic [0:0] f2328_clk;
  logic [0:0] f2328_rst;
  logic [31:0] f2328_rdata;
  sr_buffer_32_1 f2328(.wen(f2328_wen), .wdata(f2328_wdata), .clk(f2328_clk), .rst(f2328_rst), .rdata(f2328_rdata));
  assign f2328_clk = clk;
  assign f2328_rst = rst;
  // Bindings to f2328

  // f2330
  logic [0:0] f2330_wen;
  logic [31:0] f2330_wdata;
  logic [0:0] f2330_clk;
  logic [0:0] f2330_rst;
  logic [31:0] f2330_rdata;
  sr_buffer_32_1 f2330(.wen(f2330_wen), .wdata(f2330_wdata), .clk(f2330_clk), .rst(f2330_rst), .rdata(f2330_rdata));
  assign f2330_clk = clk;
  assign f2330_rst = rst;
  // Bindings to f2330

  // f2332
  logic [0:0] f2332_wen;
  logic [31:0] f2332_wdata;
  logic [0:0] f2332_clk;
  logic [0:0] f2332_rst;
  logic [31:0] f2332_rdata;
  sr_buffer_32_1 f2332(.wen(f2332_wen), .wdata(f2332_wdata), .clk(f2332_clk), .rst(f2332_rst), .rdata(f2332_rdata));
  assign f2332_clk = clk;
  assign f2332_rst = rst;
  // Bindings to f2332

  // f2334
  logic [0:0] f2334_wen;
  logic [31:0] f2334_wdata;
  logic [0:0] f2334_clk;
  logic [0:0] f2334_rst;
  logic [31:0] f2334_rdata;
  sr_buffer_32_1 f2334(.wen(f2334_wen), .wdata(f2334_wdata), .clk(f2334_clk), .rst(f2334_rst), .rdata(f2334_rdata));
  assign f2334_clk = clk;
  assign f2334_rst = rst;
  // Bindings to f2334

  // f2336
  logic [0:0] f2336_wen;
  logic [31:0] f2336_wdata;
  logic [0:0] f2336_clk;
  logic [0:0] f2336_rst;
  logic [31:0] f2336_rdata;
  sr_buffer_32_1 f2336(.wen(f2336_wen), .wdata(f2336_wdata), .clk(f2336_clk), .rst(f2336_rst), .rdata(f2336_rdata));
  assign f2336_clk = clk;
  assign f2336_rst = rst;
  // Bindings to f2336

  // f2338
  logic [0:0] f2338_wen;
  logic [31:0] f2338_wdata;
  logic [0:0] f2338_clk;
  logic [0:0] f2338_rst;
  logic [31:0] f2338_rdata;
  sr_buffer_32_1 f2338(.wen(f2338_wen), .wdata(f2338_wdata), .clk(f2338_clk), .rst(f2338_rst), .rdata(f2338_rdata));
  assign f2338_clk = clk;
  assign f2338_rst = rst;
  // Bindings to f2338

  // f2340
  logic [0:0] f2340_wen;
  logic [31:0] f2340_wdata;
  logic [0:0] f2340_clk;
  logic [0:0] f2340_rst;
  logic [31:0] f2340_rdata;
  sr_buffer_32_1 f2340(.wen(f2340_wen), .wdata(f2340_wdata), .clk(f2340_clk), .rst(f2340_rst), .rdata(f2340_rdata));
  assign f2340_clk = clk;
  assign f2340_rst = rst;
  // Bindings to f2340

  // f2342
  logic [0:0] f2342_wen;
  logic [31:0] f2342_wdata;
  logic [0:0] f2342_clk;
  logic [0:0] f2342_rst;
  logic [31:0] f2342_rdata;
  sr_buffer_32_1 f2342(.wen(f2342_wen), .wdata(f2342_wdata), .clk(f2342_clk), .rst(f2342_rst), .rdata(f2342_rdata));
  assign f2342_clk = clk;
  assign f2342_rst = rst;
  // Bindings to f2342

  // f2344
  logic [0:0] f2344_wen;
  logic [31:0] f2344_wdata;
  logic [0:0] f2344_clk;
  logic [0:0] f2344_rst;
  logic [31:0] f2344_rdata;
  sr_buffer_32_1 f2344(.wen(f2344_wen), .wdata(f2344_wdata), .clk(f2344_clk), .rst(f2344_rst), .rdata(f2344_rdata));
  assign f2344_clk = clk;
  assign f2344_rst = rst;
  // Bindings to f2344

  // f2346
  logic [0:0] f2346_wen;
  logic [31:0] f2346_wdata;
  logic [0:0] f2346_clk;
  logic [0:0] f2346_rst;
  logic [31:0] f2346_rdata;
  sr_buffer_32_1 f2346(.wen(f2346_wen), .wdata(f2346_wdata), .clk(f2346_clk), .rst(f2346_rst), .rdata(f2346_rdata));
  assign f2346_clk = clk;
  assign f2346_rst = rst;
  // Bindings to f2346

  // f2348
  logic [0:0] f2348_wen;
  logic [31:0] f2348_wdata;
  logic [0:0] f2348_clk;
  logic [0:0] f2348_rst;
  logic [31:0] f2348_rdata;
  sr_buffer_32_1 f2348(.wen(f2348_wen), .wdata(f2348_wdata), .clk(f2348_clk), .rst(f2348_rst), .rdata(f2348_rdata));
  assign f2348_clk = clk;
  assign f2348_rst = rst;
  // Bindings to f2348

  // f2350
  logic [0:0] f2350_wen;
  logic [31:0] f2350_wdata;
  logic [0:0] f2350_clk;
  logic [0:0] f2350_rst;
  logic [31:0] f2350_rdata;
  sr_buffer_32_1 f2350(.wen(f2350_wen), .wdata(f2350_wdata), .clk(f2350_clk), .rst(f2350_rst), .rdata(f2350_rdata));
  assign f2350_clk = clk;
  assign f2350_rst = rst;
  // Bindings to f2350

  // f2352
  logic [0:0] f2352_wen;
  logic [31:0] f2352_wdata;
  logic [0:0] f2352_clk;
  logic [0:0] f2352_rst;
  logic [31:0] f2352_rdata;
  sr_buffer_32_1 f2352(.wen(f2352_wen), .wdata(f2352_wdata), .clk(f2352_clk), .rst(f2352_rst), .rdata(f2352_rdata));
  assign f2352_clk = clk;
  assign f2352_rst = rst;
  // Bindings to f2352

  // f2354
  logic [0:0] f2354_wen;
  logic [31:0] f2354_wdata;
  logic [0:0] f2354_clk;
  logic [0:0] f2354_rst;
  logic [31:0] f2354_rdata;
  sr_buffer_32_1 f2354(.wen(f2354_wen), .wdata(f2354_wdata), .clk(f2354_clk), .rst(f2354_rst), .rdata(f2354_rdata));
  assign f2354_clk = clk;
  assign f2354_rst = rst;
  // Bindings to f2354

  // f2356
  logic [0:0] f2356_wen;
  logic [31:0] f2356_wdata;
  logic [0:0] f2356_clk;
  logic [0:0] f2356_rst;
  logic [31:0] f2356_rdata;
  sr_buffer_32_1 f2356(.wen(f2356_wen), .wdata(f2356_wdata), .clk(f2356_clk), .rst(f2356_rst), .rdata(f2356_rdata));
  assign f2356_clk = clk;
  assign f2356_rst = rst;
  // Bindings to f2356

  // f2358
  logic [0:0] f2358_wen;
  logic [31:0] f2358_wdata;
  logic [0:0] f2358_clk;
  logic [0:0] f2358_rst;
  logic [31:0] f2358_rdata;
  sr_buffer_32_1 f2358(.wen(f2358_wen), .wdata(f2358_wdata), .clk(f2358_clk), .rst(f2358_rst), .rdata(f2358_rdata));
  assign f2358_clk = clk;
  assign f2358_rst = rst;
  // Bindings to f2358

  // f2360
  logic [0:0] f2360_wen;
  logic [31:0] f2360_wdata;
  logic [0:0] f2360_clk;
  logic [0:0] f2360_rst;
  logic [31:0] f2360_rdata;
  sr_buffer_32_1 f2360(.wen(f2360_wen), .wdata(f2360_wdata), .clk(f2360_clk), .rst(f2360_rst), .rdata(f2360_rdata));
  assign f2360_clk = clk;
  assign f2360_rst = rst;
  // Bindings to f2360

  // f2362
  logic [0:0] f2362_wen;
  logic [31:0] f2362_wdata;
  logic [0:0] f2362_clk;
  logic [0:0] f2362_rst;
  logic [31:0] f2362_rdata;
  sr_buffer_32_1 f2362(.wen(f2362_wen), .wdata(f2362_wdata), .clk(f2362_clk), .rst(f2362_rst), .rdata(f2362_rdata));
  assign f2362_clk = clk;
  assign f2362_rst = rst;
  // Bindings to f2362

  // f2364
  logic [0:0] f2364_wen;
  logic [31:0] f2364_wdata;
  logic [0:0] f2364_clk;
  logic [0:0] f2364_rst;
  logic [31:0] f2364_rdata;
  sr_buffer_32_1 f2364(.wen(f2364_wen), .wdata(f2364_wdata), .clk(f2364_clk), .rst(f2364_rst), .rdata(f2364_rdata));
  assign f2364_clk = clk;
  assign f2364_rst = rst;
  // Bindings to f2364

  // f2366
  logic [0:0] f2366_wen;
  logic [31:0] f2366_wdata;
  logic [0:0] f2366_clk;
  logic [0:0] f2366_rst;
  logic [31:0] f2366_rdata;
  sr_buffer_32_1 f2366(.wen(f2366_wen), .wdata(f2366_wdata), .clk(f2366_clk), .rst(f2366_rst), .rdata(f2366_rdata));
  assign f2366_clk = clk;
  assign f2366_rst = rst;
  // Bindings to f2366

  // f2368
  logic [0:0] f2368_wen;
  logic [31:0] f2368_wdata;
  logic [0:0] f2368_clk;
  logic [0:0] f2368_rst;
  logic [31:0] f2368_rdata;
  sr_buffer_32_1 f2368(.wen(f2368_wen), .wdata(f2368_wdata), .clk(f2368_clk), .rst(f2368_rst), .rdata(f2368_rdata));
  assign f2368_clk = clk;
  assign f2368_rst = rst;
  // Bindings to f2368

  // f2370
  logic [0:0] f2370_wen;
  logic [31:0] f2370_wdata;
  logic [0:0] f2370_clk;
  logic [0:0] f2370_rst;
  logic [31:0] f2370_rdata;
  sr_buffer_32_1 f2370(.wen(f2370_wen), .wdata(f2370_wdata), .clk(f2370_clk), .rst(f2370_rst), .rdata(f2370_rdata));
  assign f2370_clk = clk;
  assign f2370_rst = rst;
  // Bindings to f2370

  // f2372
  logic [0:0] f2372_wen;
  logic [31:0] f2372_wdata;
  logic [0:0] f2372_clk;
  logic [0:0] f2372_rst;
  logic [31:0] f2372_rdata;
  sr_buffer_32_1 f2372(.wen(f2372_wen), .wdata(f2372_wdata), .clk(f2372_clk), .rst(f2372_rst), .rdata(f2372_rdata));
  assign f2372_clk = clk;
  assign f2372_rst = rst;
  // Bindings to f2372

  // f2374
  logic [0:0] f2374_wen;
  logic [31:0] f2374_wdata;
  logic [0:0] f2374_clk;
  logic [0:0] f2374_rst;
  logic [31:0] f2374_rdata;
  sr_buffer_32_1 f2374(.wen(f2374_wen), .wdata(f2374_wdata), .clk(f2374_clk), .rst(f2374_rst), .rdata(f2374_rdata));
  assign f2374_clk = clk;
  assign f2374_rst = rst;
  // Bindings to f2374

  // f2376
  logic [0:0] f2376_wen;
  logic [31:0] f2376_wdata;
  logic [0:0] f2376_clk;
  logic [0:0] f2376_rst;
  logic [31:0] f2376_rdata;
  sr_buffer_32_1 f2376(.wen(f2376_wen), .wdata(f2376_wdata), .clk(f2376_clk), .rst(f2376_rst), .rdata(f2376_rdata));
  assign f2376_clk = clk;
  assign f2376_rst = rst;
  // Bindings to f2376

  // f2378
  logic [0:0] f2378_wen;
  logic [31:0] f2378_wdata;
  logic [0:0] f2378_clk;
  logic [0:0] f2378_rst;
  logic [31:0] f2378_rdata;
  sr_buffer_32_1 f2378(.wen(f2378_wen), .wdata(f2378_wdata), .clk(f2378_clk), .rst(f2378_rst), .rdata(f2378_rdata));
  assign f2378_clk = clk;
  assign f2378_rst = rst;
  // Bindings to f2378

  // f2380
  logic [0:0] f2380_wen;
  logic [31:0] f2380_wdata;
  logic [0:0] f2380_clk;
  logic [0:0] f2380_rst;
  logic [31:0] f2380_rdata;
  sr_buffer_32_1 f2380(.wen(f2380_wen), .wdata(f2380_wdata), .clk(f2380_clk), .rst(f2380_rst), .rdata(f2380_rdata));
  assign f2380_clk = clk;
  assign f2380_rst = rst;
  // Bindings to f2380

  // f2382
  logic [0:0] f2382_wen;
  logic [31:0] f2382_wdata;
  logic [0:0] f2382_clk;
  logic [0:0] f2382_rst;
  logic [31:0] f2382_rdata;
  sr_buffer_32_1 f2382(.wen(f2382_wen), .wdata(f2382_wdata), .clk(f2382_clk), .rst(f2382_rst), .rdata(f2382_rdata));
  assign f2382_clk = clk;
  assign f2382_rst = rst;
  // Bindings to f2382

  // f2384
  logic [0:0] f2384_wen;
  logic [31:0] f2384_wdata;
  logic [0:0] f2384_clk;
  logic [0:0] f2384_rst;
  logic [31:0] f2384_rdata;
  sr_buffer_32_1 f2384(.wen(f2384_wen), .wdata(f2384_wdata), .clk(f2384_clk), .rst(f2384_rst), .rdata(f2384_rdata));
  assign f2384_clk = clk;
  assign f2384_rst = rst;
  // Bindings to f2384

  // f2386
  logic [0:0] f2386_wen;
  logic [31:0] f2386_wdata;
  logic [0:0] f2386_clk;
  logic [0:0] f2386_rst;
  logic [31:0] f2386_rdata;
  sr_buffer_32_1 f2386(.wen(f2386_wen), .wdata(f2386_wdata), .clk(f2386_clk), .rst(f2386_rst), .rdata(f2386_rdata));
  assign f2386_clk = clk;
  assign f2386_rst = rst;
  // Bindings to f2386

  // f2388
  logic [0:0] f2388_wen;
  logic [31:0] f2388_wdata;
  logic [0:0] f2388_clk;
  logic [0:0] f2388_rst;
  logic [31:0] f2388_rdata;
  sr_buffer_32_1 f2388(.wen(f2388_wen), .wdata(f2388_wdata), .clk(f2388_clk), .rst(f2388_rst), .rdata(f2388_rdata));
  assign f2388_clk = clk;
  assign f2388_rst = rst;
  // Bindings to f2388

  // f2390
  logic [0:0] f2390_wen;
  logic [31:0] f2390_wdata;
  logic [0:0] f2390_clk;
  logic [0:0] f2390_rst;
  logic [31:0] f2390_rdata;
  sr_buffer_32_1 f2390(.wen(f2390_wen), .wdata(f2390_wdata), .clk(f2390_clk), .rst(f2390_rst), .rdata(f2390_rdata));
  assign f2390_clk = clk;
  assign f2390_rst = rst;
  // Bindings to f2390

  // f2392
  logic [0:0] f2392_wen;
  logic [31:0] f2392_wdata;
  logic [0:0] f2392_clk;
  logic [0:0] f2392_rst;
  logic [31:0] f2392_rdata;
  sr_buffer_32_1 f2392(.wen(f2392_wen), .wdata(f2392_wdata), .clk(f2392_clk), .rst(f2392_rst), .rdata(f2392_rdata));
  assign f2392_clk = clk;
  assign f2392_rst = rst;
  // Bindings to f2392

  // f2394
  logic [0:0] f2394_wen;
  logic [31:0] f2394_wdata;
  logic [0:0] f2394_clk;
  logic [0:0] f2394_rst;
  logic [31:0] f2394_rdata;
  sr_buffer_32_1 f2394(.wen(f2394_wen), .wdata(f2394_wdata), .clk(f2394_clk), .rst(f2394_rst), .rdata(f2394_rdata));
  assign f2394_clk = clk;
  assign f2394_rst = rst;
  // Bindings to f2394

  // f2396
  logic [0:0] f2396_wen;
  logic [31:0] f2396_wdata;
  logic [0:0] f2396_clk;
  logic [0:0] f2396_rst;
  logic [31:0] f2396_rdata;
  sr_buffer_32_1 f2396(.wen(f2396_wen), .wdata(f2396_wdata), .clk(f2396_clk), .rst(f2396_rst), .rdata(f2396_rdata));
  assign f2396_clk = clk;
  assign f2396_rst = rst;
  // Bindings to f2396

  // f2398
  logic [0:0] f2398_wen;
  logic [31:0] f2398_wdata;
  logic [0:0] f2398_clk;
  logic [0:0] f2398_rst;
  logic [31:0] f2398_rdata;
  sr_buffer_32_1 f2398(.wen(f2398_wen), .wdata(f2398_wdata), .clk(f2398_clk), .rst(f2398_rst), .rdata(f2398_rdata));
  assign f2398_clk = clk;
  assign f2398_rst = rst;
  // Bindings to f2398

  // f2400
  logic [0:0] f2400_wen;
  logic [31:0] f2400_wdata;
  logic [0:0] f2400_clk;
  logic [0:0] f2400_rst;
  logic [31:0] f2400_rdata;
  sr_buffer_32_1 f2400(.wen(f2400_wen), .wdata(f2400_wdata), .clk(f2400_clk), .rst(f2400_rst), .rdata(f2400_rdata));
  assign f2400_clk = clk;
  assign f2400_rst = rst;
  // Bindings to f2400

  // f2402
  logic [0:0] f2402_wen;
  logic [31:0] f2402_wdata;
  logic [0:0] f2402_clk;
  logic [0:0] f2402_rst;
  logic [31:0] f2402_rdata;
  sr_buffer_32_1 f2402(.wen(f2402_wen), .wdata(f2402_wdata), .clk(f2402_clk), .rst(f2402_rst), .rdata(f2402_rdata));
  assign f2402_clk = clk;
  assign f2402_rst = rst;
  // Bindings to f2402

  // f2404
  logic [0:0] f2404_wen;
  logic [31:0] f2404_wdata;
  logic [0:0] f2404_clk;
  logic [0:0] f2404_rst;
  logic [31:0] f2404_rdata;
  sr_buffer_32_1 f2404(.wen(f2404_wen), .wdata(f2404_wdata), .clk(f2404_clk), .rst(f2404_rst), .rdata(f2404_rdata));
  assign f2404_clk = clk;
  assign f2404_rst = rst;
  // Bindings to f2404

  // f2406
  logic [0:0] f2406_wen;
  logic [31:0] f2406_wdata;
  logic [0:0] f2406_clk;
  logic [0:0] f2406_rst;
  logic [31:0] f2406_rdata;
  sr_buffer_32_1 f2406(.wen(f2406_wen), .wdata(f2406_wdata), .clk(f2406_clk), .rst(f2406_rst), .rdata(f2406_rdata));
  assign f2406_clk = clk;
  assign f2406_rst = rst;
  // Bindings to f2406

  // f2408
  logic [0:0] f2408_wen;
  logic [31:0] f2408_wdata;
  logic [0:0] f2408_clk;
  logic [0:0] f2408_rst;
  logic [31:0] f2408_rdata;
  sr_buffer_32_1 f2408(.wen(f2408_wen), .wdata(f2408_wdata), .clk(f2408_clk), .rst(f2408_rst), .rdata(f2408_rdata));
  assign f2408_clk = clk;
  assign f2408_rst = rst;
  // Bindings to f2408

  // f2410
  logic [0:0] f2410_wen;
  logic [31:0] f2410_wdata;
  logic [0:0] f2410_clk;
  logic [0:0] f2410_rst;
  logic [31:0] f2410_rdata;
  sr_buffer_32_1 f2410(.wen(f2410_wen), .wdata(f2410_wdata), .clk(f2410_clk), .rst(f2410_rst), .rdata(f2410_rdata));
  assign f2410_clk = clk;
  assign f2410_rst = rst;
  // Bindings to f2410

  // f2412
  logic [0:0] f2412_wen;
  logic [31:0] f2412_wdata;
  logic [0:0] f2412_clk;
  logic [0:0] f2412_rst;
  logic [31:0] f2412_rdata;
  sr_buffer_32_1 f2412(.wen(f2412_wen), .wdata(f2412_wdata), .clk(f2412_clk), .rst(f2412_rst), .rdata(f2412_rdata));
  assign f2412_clk = clk;
  assign f2412_rst = rst;
  // Bindings to f2412

  // f2414
  logic [0:0] f2414_wen;
  logic [31:0] f2414_wdata;
  logic [0:0] f2414_clk;
  logic [0:0] f2414_rst;
  logic [31:0] f2414_rdata;
  sr_buffer_32_1 f2414(.wen(f2414_wen), .wdata(f2414_wdata), .clk(f2414_clk), .rst(f2414_rst), .rdata(f2414_rdata));
  assign f2414_clk = clk;
  assign f2414_rst = rst;
  // Bindings to f2414

  // f2416
  logic [0:0] f2416_wen;
  logic [31:0] f2416_wdata;
  logic [0:0] f2416_clk;
  logic [0:0] f2416_rst;
  logic [31:0] f2416_rdata;
  sr_buffer_32_1 f2416(.wen(f2416_wen), .wdata(f2416_wdata), .clk(f2416_clk), .rst(f2416_rst), .rdata(f2416_rdata));
  assign f2416_clk = clk;
  assign f2416_rst = rst;
  // Bindings to f2416

  // f2418
  logic [0:0] f2418_wen;
  logic [31:0] f2418_wdata;
  logic [0:0] f2418_clk;
  logic [0:0] f2418_rst;
  logic [31:0] f2418_rdata;
  sr_buffer_32_1 f2418(.wen(f2418_wen), .wdata(f2418_wdata), .clk(f2418_clk), .rst(f2418_rst), .rdata(f2418_rdata));
  assign f2418_clk = clk;
  assign f2418_rst = rst;
  // Bindings to f2418

  // f2420
  logic [0:0] f2420_wen;
  logic [31:0] f2420_wdata;
  logic [0:0] f2420_clk;
  logic [0:0] f2420_rst;
  logic [31:0] f2420_rdata;
  sr_buffer_32_1 f2420(.wen(f2420_wen), .wdata(f2420_wdata), .clk(f2420_clk), .rst(f2420_rst), .rdata(f2420_rdata));
  assign f2420_clk = clk;
  assign f2420_rst = rst;
  // Bindings to f2420

  // f2422
  logic [0:0] f2422_wen;
  logic [31:0] f2422_wdata;
  logic [0:0] f2422_clk;
  logic [0:0] f2422_rst;
  logic [31:0] f2422_rdata;
  sr_buffer_32_1 f2422(.wen(f2422_wen), .wdata(f2422_wdata), .clk(f2422_clk), .rst(f2422_rst), .rdata(f2422_rdata));
  assign f2422_clk = clk;
  assign f2422_rst = rst;
  // Bindings to f2422

  // f2424
  logic [0:0] f2424_wen;
  logic [31:0] f2424_wdata;
  logic [0:0] f2424_clk;
  logic [0:0] f2424_rst;
  logic [31:0] f2424_rdata;
  sr_buffer_32_1 f2424(.wen(f2424_wen), .wdata(f2424_wdata), .clk(f2424_clk), .rst(f2424_rst), .rdata(f2424_rdata));
  assign f2424_clk = clk;
  assign f2424_rst = rst;
  // Bindings to f2424

  // f2426
  logic [0:0] f2426_wen;
  logic [31:0] f2426_wdata;
  logic [0:0] f2426_clk;
  logic [0:0] f2426_rst;
  logic [31:0] f2426_rdata;
  sr_buffer_32_1 f2426(.wen(f2426_wen), .wdata(f2426_wdata), .clk(f2426_clk), .rst(f2426_rst), .rdata(f2426_rdata));
  assign f2426_clk = clk;
  assign f2426_rst = rst;
  // Bindings to f2426

  // f2428
  logic [0:0] f2428_wen;
  logic [31:0] f2428_wdata;
  logic [0:0] f2428_clk;
  logic [0:0] f2428_rst;
  logic [31:0] f2428_rdata;
  sr_buffer_32_1 f2428(.wen(f2428_wen), .wdata(f2428_wdata), .clk(f2428_clk), .rst(f2428_rst), .rdata(f2428_rdata));
  assign f2428_clk = clk;
  assign f2428_rst = rst;
  // Bindings to f2428

  // f2430
  logic [0:0] f2430_wen;
  logic [31:0] f2430_wdata;
  logic [0:0] f2430_clk;
  logic [0:0] f2430_rst;
  logic [31:0] f2430_rdata;
  sr_buffer_32_1 f2430(.wen(f2430_wen), .wdata(f2430_wdata), .clk(f2430_clk), .rst(f2430_rst), .rdata(f2430_rdata));
  assign f2430_clk = clk;
  assign f2430_rst = rst;
  // Bindings to f2430

  // f2432
  logic [0:0] f2432_wen;
  logic [31:0] f2432_wdata;
  logic [0:0] f2432_clk;
  logic [0:0] f2432_rst;
  logic [31:0] f2432_rdata;
  sr_buffer_32_1 f2432(.wen(f2432_wen), .wdata(f2432_wdata), .clk(f2432_clk), .rst(f2432_rst), .rdata(f2432_rdata));
  assign f2432_clk = clk;
  assign f2432_rst = rst;
  // Bindings to f2432

  // f2434
  logic [0:0] f2434_wen;
  logic [31:0] f2434_wdata;
  logic [0:0] f2434_clk;
  logic [0:0] f2434_rst;
  logic [31:0] f2434_rdata;
  sr_buffer_32_1 f2434(.wen(f2434_wen), .wdata(f2434_wdata), .clk(f2434_clk), .rst(f2434_rst), .rdata(f2434_rdata));
  assign f2434_clk = clk;
  assign f2434_rst = rst;
  // Bindings to f2434

  // f2436
  logic [0:0] f2436_wen;
  logic [31:0] f2436_wdata;
  logic [0:0] f2436_clk;
  logic [0:0] f2436_rst;
  logic [31:0] f2436_rdata;
  sr_buffer_32_1 f2436(.wen(f2436_wen), .wdata(f2436_wdata), .clk(f2436_clk), .rst(f2436_rst), .rdata(f2436_rdata));
  assign f2436_clk = clk;
  assign f2436_rst = rst;
  // Bindings to f2436

  // f2438
  logic [0:0] f2438_wen;
  logic [31:0] f2438_wdata;
  logic [0:0] f2438_clk;
  logic [0:0] f2438_rst;
  logic [31:0] f2438_rdata;
  sr_buffer_32_1 f2438(.wen(f2438_wen), .wdata(f2438_wdata), .clk(f2438_clk), .rst(f2438_rst), .rdata(f2438_rdata));
  assign f2438_clk = clk;
  assign f2438_rst = rst;
  // Bindings to f2438

  // f2440
  logic [0:0] f2440_wen;
  logic [31:0] f2440_wdata;
  logic [0:0] f2440_clk;
  logic [0:0] f2440_rst;
  logic [31:0] f2440_rdata;
  sr_buffer_32_1 f2440(.wen(f2440_wen), .wdata(f2440_wdata), .clk(f2440_clk), .rst(f2440_rst), .rdata(f2440_rdata));
  assign f2440_clk = clk;
  assign f2440_rst = rst;
  // Bindings to f2440

  // f2442
  logic [0:0] f2442_wen;
  logic [31:0] f2442_wdata;
  logic [0:0] f2442_clk;
  logic [0:0] f2442_rst;
  logic [31:0] f2442_rdata;
  sr_buffer_32_1 f2442(.wen(f2442_wen), .wdata(f2442_wdata), .clk(f2442_clk), .rst(f2442_rst), .rdata(f2442_rdata));
  assign f2442_clk = clk;
  assign f2442_rst = rst;
  // Bindings to f2442

  // f2444
  logic [0:0] f2444_wen;
  logic [31:0] f2444_wdata;
  logic [0:0] f2444_clk;
  logic [0:0] f2444_rst;
  logic [31:0] f2444_rdata;
  sr_buffer_32_1 f2444(.wen(f2444_wen), .wdata(f2444_wdata), .clk(f2444_clk), .rst(f2444_rst), .rdata(f2444_rdata));
  assign f2444_clk = clk;
  assign f2444_rst = rst;
  // Bindings to f2444

  // f2446
  logic [0:0] f2446_wen;
  logic [31:0] f2446_wdata;
  logic [0:0] f2446_clk;
  logic [0:0] f2446_rst;
  logic [31:0] f2446_rdata;
  sr_buffer_32_1 f2446(.wen(f2446_wen), .wdata(f2446_wdata), .clk(f2446_clk), .rst(f2446_rst), .rdata(f2446_rdata));
  assign f2446_clk = clk;
  assign f2446_rst = rst;
  // Bindings to f2446

  // f2448
  logic [0:0] f2448_wen;
  logic [31:0] f2448_wdata;
  logic [0:0] f2448_clk;
  logic [0:0] f2448_rst;
  logic [31:0] f2448_rdata;
  sr_buffer_32_1 f2448(.wen(f2448_wen), .wdata(f2448_wdata), .clk(f2448_clk), .rst(f2448_rst), .rdata(f2448_rdata));
  assign f2448_clk = clk;
  assign f2448_rst = rst;
  // Bindings to f2448

  // f2450
  logic [0:0] f2450_wen;
  logic [31:0] f2450_wdata;
  logic [0:0] f2450_clk;
  logic [0:0] f2450_rst;
  logic [31:0] f2450_rdata;
  sr_buffer_32_1 f2450(.wen(f2450_wen), .wdata(f2450_wdata), .clk(f2450_clk), .rst(f2450_rst), .rdata(f2450_rdata));
  assign f2450_clk = clk;
  assign f2450_rst = rst;
  // Bindings to f2450

  // f2452
  logic [0:0] f2452_wen;
  logic [31:0] f2452_wdata;
  logic [0:0] f2452_clk;
  logic [0:0] f2452_rst;
  logic [31:0] f2452_rdata;
  sr_buffer_32_1 f2452(.wen(f2452_wen), .wdata(f2452_wdata), .clk(f2452_clk), .rst(f2452_rst), .rdata(f2452_rdata));
  assign f2452_clk = clk;
  assign f2452_rst = rst;
  // Bindings to f2452

  // f2454
  logic [0:0] f2454_wen;
  logic [31:0] f2454_wdata;
  logic [0:0] f2454_clk;
  logic [0:0] f2454_rst;
  logic [31:0] f2454_rdata;
  sr_buffer_32_1 f2454(.wen(f2454_wen), .wdata(f2454_wdata), .clk(f2454_clk), .rst(f2454_rst), .rdata(f2454_rdata));
  assign f2454_clk = clk;
  assign f2454_rst = rst;
  // Bindings to f2454

  // f2456
  logic [0:0] f2456_wen;
  logic [31:0] f2456_wdata;
  logic [0:0] f2456_clk;
  logic [0:0] f2456_rst;
  logic [31:0] f2456_rdata;
  sr_buffer_32_1 f2456(.wen(f2456_wen), .wdata(f2456_wdata), .clk(f2456_clk), .rst(f2456_rst), .rdata(f2456_rdata));
  assign f2456_clk = clk;
  assign f2456_rst = rst;
  // Bindings to f2456

  // f2458
  logic [0:0] f2458_wen;
  logic [31:0] f2458_wdata;
  logic [0:0] f2458_clk;
  logic [0:0] f2458_rst;
  logic [31:0] f2458_rdata;
  sr_buffer_32_1 f2458(.wen(f2458_wen), .wdata(f2458_wdata), .clk(f2458_clk), .rst(f2458_rst), .rdata(f2458_rdata));
  assign f2458_clk = clk;
  assign f2458_rst = rst;
  // Bindings to f2458

  // f2460
  logic [0:0] f2460_wen;
  logic [31:0] f2460_wdata;
  logic [0:0] f2460_clk;
  logic [0:0] f2460_rst;
  logic [31:0] f2460_rdata;
  sr_buffer_32_1 f2460(.wen(f2460_wen), .wdata(f2460_wdata), .clk(f2460_clk), .rst(f2460_rst), .rdata(f2460_rdata));
  assign f2460_clk = clk;
  assign f2460_rst = rst;
  // Bindings to f2460

  // f2462
  logic [0:0] f2462_wen;
  logic [31:0] f2462_wdata;
  logic [0:0] f2462_clk;
  logic [0:0] f2462_rst;
  logic [31:0] f2462_rdata;
  sr_buffer_32_1 f2462(.wen(f2462_wen), .wdata(f2462_wdata), .clk(f2462_clk), .rst(f2462_rst), .rdata(f2462_rdata));
  assign f2462_clk = clk;
  assign f2462_rst = rst;
  // Bindings to f2462

  // f2464
  logic [0:0] f2464_wen;
  logic [31:0] f2464_wdata;
  logic [0:0] f2464_clk;
  logic [0:0] f2464_rst;
  logic [31:0] f2464_rdata;
  sr_buffer_32_1 f2464(.wen(f2464_wen), .wdata(f2464_wdata), .clk(f2464_clk), .rst(f2464_rst), .rdata(f2464_rdata));
  assign f2464_clk = clk;
  assign f2464_rst = rst;
  // Bindings to f2464

  // f2466
  logic [0:0] f2466_wen;
  logic [31:0] f2466_wdata;
  logic [0:0] f2466_clk;
  logic [0:0] f2466_rst;
  logic [31:0] f2466_rdata;
  sr_buffer_32_1 f2466(.wen(f2466_wen), .wdata(f2466_wdata), .clk(f2466_clk), .rst(f2466_rst), .rdata(f2466_rdata));
  assign f2466_clk = clk;
  assign f2466_rst = rst;
  // Bindings to f2466

  // f2468
  logic [0:0] f2468_wen;
  logic [31:0] f2468_wdata;
  logic [0:0] f2468_clk;
  logic [0:0] f2468_rst;
  logic [31:0] f2468_rdata;
  sr_buffer_32_1 f2468(.wen(f2468_wen), .wdata(f2468_wdata), .clk(f2468_clk), .rst(f2468_rst), .rdata(f2468_rdata));
  assign f2468_clk = clk;
  assign f2468_rst = rst;
  // Bindings to f2468

  // f2470
  logic [0:0] f2470_wen;
  logic [31:0] f2470_wdata;
  logic [0:0] f2470_clk;
  logic [0:0] f2470_rst;
  logic [31:0] f2470_rdata;
  sr_buffer_32_1 f2470(.wen(f2470_wen), .wdata(f2470_wdata), .clk(f2470_clk), .rst(f2470_rst), .rdata(f2470_rdata));
  assign f2470_clk = clk;
  assign f2470_rst = rst;
  // Bindings to f2470

  // f2472
  logic [0:0] f2472_wen;
  logic [31:0] f2472_wdata;
  logic [0:0] f2472_clk;
  logic [0:0] f2472_rst;
  logic [31:0] f2472_rdata;
  sr_buffer_32_1 f2472(.wen(f2472_wen), .wdata(f2472_wdata), .clk(f2472_clk), .rst(f2472_rst), .rdata(f2472_rdata));
  assign f2472_clk = clk;
  assign f2472_rst = rst;
  // Bindings to f2472

  // f2474
  logic [0:0] f2474_wen;
  logic [31:0] f2474_wdata;
  logic [0:0] f2474_clk;
  logic [0:0] f2474_rst;
  logic [31:0] f2474_rdata;
  sr_buffer_32_1 f2474(.wen(f2474_wen), .wdata(f2474_wdata), .clk(f2474_clk), .rst(f2474_rst), .rdata(f2474_rdata));
  assign f2474_clk = clk;
  assign f2474_rst = rst;
  // Bindings to f2474

  // f2476
  logic [0:0] f2476_wen;
  logic [31:0] f2476_wdata;
  logic [0:0] f2476_clk;
  logic [0:0] f2476_rst;
  logic [31:0] f2476_rdata;
  sr_buffer_32_1 f2476(.wen(f2476_wen), .wdata(f2476_wdata), .clk(f2476_clk), .rst(f2476_rst), .rdata(f2476_rdata));
  assign f2476_clk = clk;
  assign f2476_rst = rst;
  // Bindings to f2476

  // f2478
  logic [0:0] f2478_wen;
  logic [31:0] f2478_wdata;
  logic [0:0] f2478_clk;
  logic [0:0] f2478_rst;
  logic [31:0] f2478_rdata;
  sr_buffer_32_1 f2478(.wen(f2478_wen), .wdata(f2478_wdata), .clk(f2478_clk), .rst(f2478_rst), .rdata(f2478_rdata));
  assign f2478_clk = clk;
  assign f2478_rst = rst;
  // Bindings to f2478

  // f2480
  logic [0:0] f2480_wen;
  logic [31:0] f2480_wdata;
  logic [0:0] f2480_clk;
  logic [0:0] f2480_rst;
  logic [31:0] f2480_rdata;
  sr_buffer_32_1 f2480(.wen(f2480_wen), .wdata(f2480_wdata), .clk(f2480_clk), .rst(f2480_rst), .rdata(f2480_rdata));
  assign f2480_clk = clk;
  assign f2480_rst = rst;
  // Bindings to f2480

  // f2482
  logic [0:0] f2482_wen;
  logic [31:0] f2482_wdata;
  logic [0:0] f2482_clk;
  logic [0:0] f2482_rst;
  logic [31:0] f2482_rdata;
  sr_buffer_32_1 f2482(.wen(f2482_wen), .wdata(f2482_wdata), .clk(f2482_clk), .rst(f2482_rst), .rdata(f2482_rdata));
  assign f2482_clk = clk;
  assign f2482_rst = rst;
  // Bindings to f2482

  // f2484
  logic [0:0] f2484_wen;
  logic [31:0] f2484_wdata;
  logic [0:0] f2484_clk;
  logic [0:0] f2484_rst;
  logic [31:0] f2484_rdata;
  sr_buffer_32_1 f2484(.wen(f2484_wen), .wdata(f2484_wdata), .clk(f2484_clk), .rst(f2484_rst), .rdata(f2484_rdata));
  assign f2484_clk = clk;
  assign f2484_rst = rst;
  // Bindings to f2484

  // f2486
  logic [0:0] f2486_wen;
  logic [31:0] f2486_wdata;
  logic [0:0] f2486_clk;
  logic [0:0] f2486_rst;
  logic [31:0] f2486_rdata;
  sr_buffer_32_1 f2486(.wen(f2486_wen), .wdata(f2486_wdata), .clk(f2486_clk), .rst(f2486_rst), .rdata(f2486_rdata));
  assign f2486_clk = clk;
  assign f2486_rst = rst;
  // Bindings to f2486

  // f2488
  logic [0:0] f2488_wen;
  logic [31:0] f2488_wdata;
  logic [0:0] f2488_clk;
  logic [0:0] f2488_rst;
  logic [31:0] f2488_rdata;
  sr_buffer_32_1 f2488(.wen(f2488_wen), .wdata(f2488_wdata), .clk(f2488_clk), .rst(f2488_rst), .rdata(f2488_rdata));
  assign f2488_clk = clk;
  assign f2488_rst = rst;
  // Bindings to f2488

  // f2490
  logic [0:0] f2490_wen;
  logic [31:0] f2490_wdata;
  logic [0:0] f2490_clk;
  logic [0:0] f2490_rst;
  logic [31:0] f2490_rdata;
  sr_buffer_32_1 f2490(.wen(f2490_wen), .wdata(f2490_wdata), .clk(f2490_clk), .rst(f2490_rst), .rdata(f2490_rdata));
  assign f2490_clk = clk;
  assign f2490_rst = rst;
  // Bindings to f2490

  // f2492
  logic [0:0] f2492_wen;
  logic [31:0] f2492_wdata;
  logic [0:0] f2492_clk;
  logic [0:0] f2492_rst;
  logic [31:0] f2492_rdata;
  sr_buffer_32_1 f2492(.wen(f2492_wen), .wdata(f2492_wdata), .clk(f2492_clk), .rst(f2492_rst), .rdata(f2492_rdata));
  assign f2492_clk = clk;
  assign f2492_rst = rst;
  // Bindings to f2492

  // f2494
  logic [0:0] f2494_wen;
  logic [31:0] f2494_wdata;
  logic [0:0] f2494_clk;
  logic [0:0] f2494_rst;
  logic [31:0] f2494_rdata;
  sr_buffer_32_1 f2494(.wen(f2494_wen), .wdata(f2494_wdata), .clk(f2494_clk), .rst(f2494_rst), .rdata(f2494_rdata));
  assign f2494_clk = clk;
  assign f2494_rst = rst;
  // Bindings to f2494

  // f2496
  logic [0:0] f2496_wen;
  logic [31:0] f2496_wdata;
  logic [0:0] f2496_clk;
  logic [0:0] f2496_rst;
  logic [31:0] f2496_rdata;
  sr_buffer_32_1 f2496(.wen(f2496_wen), .wdata(f2496_wdata), .clk(f2496_clk), .rst(f2496_rst), .rdata(f2496_rdata));
  assign f2496_clk = clk;
  assign f2496_rst = rst;
  // Bindings to f2496

  // f2498
  logic [0:0] f2498_wen;
  logic [31:0] f2498_wdata;
  logic [0:0] f2498_clk;
  logic [0:0] f2498_rst;
  logic [31:0] f2498_rdata;
  sr_buffer_32_1 f2498(.wen(f2498_wen), .wdata(f2498_wdata), .clk(f2498_clk), .rst(f2498_rst), .rdata(f2498_rdata));
  assign f2498_clk = clk;
  assign f2498_rst = rst;
  // Bindings to f2498

  // f2500
  logic [0:0] f2500_wen;
  logic [31:0] f2500_wdata;
  logic [0:0] f2500_clk;
  logic [0:0] f2500_rst;
  logic [31:0] f2500_rdata;
  sr_buffer_32_1 f2500(.wen(f2500_wen), .wdata(f2500_wdata), .clk(f2500_clk), .rst(f2500_rst), .rdata(f2500_rdata));
  assign f2500_clk = clk;
  assign f2500_rst = rst;
  // Bindings to f2500

  // f2502
  logic [0:0] f2502_wen;
  logic [31:0] f2502_wdata;
  logic [0:0] f2502_clk;
  logic [0:0] f2502_rst;
  logic [31:0] f2502_rdata;
  sr_buffer_32_1 f2502(.wen(f2502_wen), .wdata(f2502_wdata), .clk(f2502_clk), .rst(f2502_rst), .rdata(f2502_rdata));
  assign f2502_clk = clk;
  assign f2502_rst = rst;
  // Bindings to f2502

  // f2504
  logic [0:0] f2504_wen;
  logic [31:0] f2504_wdata;
  logic [0:0] f2504_clk;
  logic [0:0] f2504_rst;
  logic [31:0] f2504_rdata;
  sr_buffer_32_1 f2504(.wen(f2504_wen), .wdata(f2504_wdata), .clk(f2504_clk), .rst(f2504_rst), .rdata(f2504_rdata));
  assign f2504_clk = clk;
  assign f2504_rst = rst;
  // Bindings to f2504

  // f2506
  logic [0:0] f2506_wen;
  logic [31:0] f2506_wdata;
  logic [0:0] f2506_clk;
  logic [0:0] f2506_rst;
  logic [31:0] f2506_rdata;
  sr_buffer_32_1 f2506(.wen(f2506_wen), .wdata(f2506_wdata), .clk(f2506_clk), .rst(f2506_rst), .rdata(f2506_rdata));
  assign f2506_clk = clk;
  assign f2506_rst = rst;
  // Bindings to f2506

  // f2508
  logic [0:0] f2508_wen;
  logic [31:0] f2508_wdata;
  logic [0:0] f2508_clk;
  logic [0:0] f2508_rst;
  logic [31:0] f2508_rdata;
  sr_buffer_32_1 f2508(.wen(f2508_wen), .wdata(f2508_wdata), .clk(f2508_clk), .rst(f2508_rst), .rdata(f2508_rdata));
  assign f2508_clk = clk;
  assign f2508_rst = rst;
  // Bindings to f2508

  // f2510
  logic [0:0] f2510_wen;
  logic [31:0] f2510_wdata;
  logic [0:0] f2510_clk;
  logic [0:0] f2510_rst;
  logic [31:0] f2510_rdata;
  sr_buffer_32_1 f2510(.wen(f2510_wen), .wdata(f2510_wdata), .clk(f2510_clk), .rst(f2510_rst), .rdata(f2510_rdata));
  assign f2510_clk = clk;
  assign f2510_rst = rst;
  // Bindings to f2510

  // f2512
  logic [0:0] f2512_wen;
  logic [31:0] f2512_wdata;
  logic [0:0] f2512_clk;
  logic [0:0] f2512_rst;
  logic [31:0] f2512_rdata;
  sr_buffer_32_1 f2512(.wen(f2512_wen), .wdata(f2512_wdata), .clk(f2512_clk), .rst(f2512_rst), .rdata(f2512_rdata));
  assign f2512_clk = clk;
  assign f2512_rst = rst;
  // Bindings to f2512

  // f2514
  logic [0:0] f2514_wen;
  logic [31:0] f2514_wdata;
  logic [0:0] f2514_clk;
  logic [0:0] f2514_rst;
  logic [31:0] f2514_rdata;
  sr_buffer_32_1 f2514(.wen(f2514_wen), .wdata(f2514_wdata), .clk(f2514_clk), .rst(f2514_rst), .rdata(f2514_rdata));
  assign f2514_clk = clk;
  assign f2514_rst = rst;
  // Bindings to f2514

  // f2516
  logic [0:0] f2516_wen;
  logic [31:0] f2516_wdata;
  logic [0:0] f2516_clk;
  logic [0:0] f2516_rst;
  logic [31:0] f2516_rdata;
  sr_buffer_32_1 f2516(.wen(f2516_wen), .wdata(f2516_wdata), .clk(f2516_clk), .rst(f2516_rst), .rdata(f2516_rdata));
  assign f2516_clk = clk;
  assign f2516_rst = rst;
  // Bindings to f2516

  // f2518
  logic [0:0] f2518_wen;
  logic [31:0] f2518_wdata;
  logic [0:0] f2518_clk;
  logic [0:0] f2518_rst;
  logic [31:0] f2518_rdata;
  sr_buffer_32_1 f2518(.wen(f2518_wen), .wdata(f2518_wdata), .clk(f2518_clk), .rst(f2518_rst), .rdata(f2518_rdata));
  assign f2518_clk = clk;
  assign f2518_rst = rst;
  // Bindings to f2518

  // f2520
  logic [0:0] f2520_wen;
  logic [31:0] f2520_wdata;
  logic [0:0] f2520_clk;
  logic [0:0] f2520_rst;
  logic [31:0] f2520_rdata;
  sr_buffer_32_1 f2520(.wen(f2520_wen), .wdata(f2520_wdata), .clk(f2520_clk), .rst(f2520_rst), .rdata(f2520_rdata));
  assign f2520_clk = clk;
  assign f2520_rst = rst;
  // Bindings to f2520

  // f2522
  logic [0:0] f2522_wen;
  logic [31:0] f2522_wdata;
  logic [0:0] f2522_clk;
  logic [0:0] f2522_rst;
  logic [31:0] f2522_rdata;
  sr_buffer_32_1 f2522(.wen(f2522_wen), .wdata(f2522_wdata), .clk(f2522_clk), .rst(f2522_rst), .rdata(f2522_rdata));
  assign f2522_clk = clk;
  assign f2522_rst = rst;
  // Bindings to f2522

  // f2524
  logic [0:0] f2524_wen;
  logic [31:0] f2524_wdata;
  logic [0:0] f2524_clk;
  logic [0:0] f2524_rst;
  logic [31:0] f2524_rdata;
  sr_buffer_32_1 f2524(.wen(f2524_wen), .wdata(f2524_wdata), .clk(f2524_clk), .rst(f2524_rst), .rdata(f2524_rdata));
  assign f2524_clk = clk;
  assign f2524_rst = rst;
  // Bindings to f2524

  // f2526
  logic [0:0] f2526_wen;
  logic [31:0] f2526_wdata;
  logic [0:0] f2526_clk;
  logic [0:0] f2526_rst;
  logic [31:0] f2526_rdata;
  sr_buffer_32_1 f2526(.wen(f2526_wen), .wdata(f2526_wdata), .clk(f2526_clk), .rst(f2526_rst), .rdata(f2526_rdata));
  assign f2526_clk = clk;
  assign f2526_rst = rst;
  // Bindings to f2526

  // f2528
  logic [0:0] f2528_wen;
  logic [31:0] f2528_wdata;
  logic [0:0] f2528_clk;
  logic [0:0] f2528_rst;
  logic [31:0] f2528_rdata;
  sr_buffer_32_1 f2528(.wen(f2528_wen), .wdata(f2528_wdata), .clk(f2528_clk), .rst(f2528_rst), .rdata(f2528_rdata));
  assign f2528_clk = clk;
  assign f2528_rst = rst;
  // Bindings to f2528

  // f2530
  logic [0:0] f2530_wen;
  logic [31:0] f2530_wdata;
  logic [0:0] f2530_clk;
  logic [0:0] f2530_rst;
  logic [31:0] f2530_rdata;
  sr_buffer_32_1 f2530(.wen(f2530_wen), .wdata(f2530_wdata), .clk(f2530_clk), .rst(f2530_rst), .rdata(f2530_rdata));
  assign f2530_clk = clk;
  assign f2530_rst = rst;
  // Bindings to f2530

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f1450
  logic [0:0] f1450_wen;
  logic [31:0] f1450_wdata;
  logic [0:0] f1450_clk;
  logic [0:0] f1450_rst;
  logic [31:0] f1450_rdata;
  sr_buffer_32_1 f1450(.wen(f1450_wen), .wdata(f1450_wdata), .clk(f1450_clk), .rst(f1450_rst), .rdata(f1450_rdata));
  assign f1450_clk = clk;
  assign f1450_rst = rst;
  // Bindings to f1450

  // f1452
  logic [0:0] f1452_wen;
  logic [31:0] f1452_wdata;
  logic [0:0] f1452_clk;
  logic [0:0] f1452_rst;
  logic [31:0] f1452_rdata;
  sr_buffer_32_1 f1452(.wen(f1452_wen), .wdata(f1452_wdata), .clk(f1452_clk), .rst(f1452_rst), .rdata(f1452_rdata));
  assign f1452_clk = clk;
  assign f1452_rst = rst;
  // Bindings to f1452

  // f1448
  logic [0:0] f1448_wen;
  logic [31:0] f1448_wdata;
  logic [0:0] f1448_clk;
  logic [0:0] f1448_rst;
  logic [31:0] f1448_rdata;
  sr_buffer_32_1 f1448(.wen(f1448_wen), .wdata(f1448_wdata), .clk(f1448_clk), .rst(f1448_rst), .rdata(f1448_rdata));
  assign f1448_clk = clk;
  assign f1448_rst = rst;
  // Bindings to f1448

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_16431 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f314
  logic [0:0] f314_wen;
  logic [31:0] f314_wdata;
  logic [0:0] f314_clk;
  logic [0:0] f314_rst;
  logic [31:0] f314_rdata;
  sr_buffer_32_1 f314(.wen(f314_wen), .wdata(f314_wdata), .clk(f314_clk), .rst(f314_rst), .rdata(f314_rdata));
  assign f314_clk = clk;
  assign f314_rst = rst;
  // Bindings to f314

  // f316
  logic [0:0] f316_wen;
  logic [31:0] f316_wdata;
  logic [0:0] f316_clk;
  logic [0:0] f316_rst;
  logic [31:0] f316_rdata;
  sr_buffer_32_1 f316(.wen(f316_wen), .wdata(f316_wdata), .clk(f316_clk), .rst(f316_rst), .rdata(f316_rdata));
  assign f316_clk = clk;
  assign f316_rst = rst;
  // Bindings to f316

  // f318
  logic [0:0] f318_wen;
  logic [31:0] f318_wdata;
  logic [0:0] f318_clk;
  logic [0:0] f318_rst;
  logic [31:0] f318_rdata;
  sr_buffer_32_1 f318(.wen(f318_wen), .wdata(f318_wdata), .clk(f318_clk), .rst(f318_rst), .rdata(f318_rdata));
  assign f318_clk = clk;
  assign f318_rst = rst;
  // Bindings to f318

  // f320
  logic [0:0] f320_wen;
  logic [31:0] f320_wdata;
  logic [0:0] f320_clk;
  logic [0:0] f320_rst;
  logic [31:0] f320_rdata;
  sr_buffer_32_1 f320(.wen(f320_wen), .wdata(f320_wdata), .clk(f320_clk), .rst(f320_rst), .rdata(f320_rdata));
  assign f320_clk = clk;
  assign f320_rst = rst;
  // Bindings to f320

  // f322
  logic [0:0] f322_wen;
  logic [31:0] f322_wdata;
  logic [0:0] f322_clk;
  logic [0:0] f322_rst;
  logic [31:0] f322_rdata;
  sr_buffer_32_1 f322(.wen(f322_wen), .wdata(f322_wdata), .clk(f322_clk), .rst(f322_rst), .rdata(f322_rdata));
  assign f322_clk = clk;
  assign f322_rst = rst;
  // Bindings to f322

  // f324
  logic [0:0] f324_wen;
  logic [31:0] f324_wdata;
  logic [0:0] f324_clk;
  logic [0:0] f324_rst;
  logic [31:0] f324_rdata;
  sr_buffer_32_1 f324(.wen(f324_wen), .wdata(f324_wdata), .clk(f324_clk), .rst(f324_rst), .rdata(f324_rdata));
  assign f324_clk = clk;
  assign f324_rst = rst;
  // Bindings to f324

  // f326
  logic [0:0] f326_wen;
  logic [31:0] f326_wdata;
  logic [0:0] f326_clk;
  logic [0:0] f326_rst;
  logic [31:0] f326_rdata;
  sr_buffer_32_1 f326(.wen(f326_wen), .wdata(f326_wdata), .clk(f326_clk), .rst(f326_rst), .rdata(f326_rdata));
  assign f326_clk = clk;
  assign f326_rst = rst;
  // Bindings to f326

  // f328
  logic [0:0] f328_wen;
  logic [31:0] f328_wdata;
  logic [0:0] f328_clk;
  logic [0:0] f328_rst;
  logic [31:0] f328_rdata;
  sr_buffer_32_1 f328(.wen(f328_wen), .wdata(f328_wdata), .clk(f328_clk), .rst(f328_rst), .rdata(f328_rdata));
  assign f328_clk = clk;
  assign f328_rst = rst;
  // Bindings to f328

  // f330
  logic [0:0] f330_wen;
  logic [31:0] f330_wdata;
  logic [0:0] f330_clk;
  logic [0:0] f330_rst;
  logic [31:0] f330_rdata;
  sr_buffer_32_1 f330(.wen(f330_wen), .wdata(f330_wdata), .clk(f330_clk), .rst(f330_rst), .rdata(f330_rdata));
  assign f330_clk = clk;
  assign f330_rst = rst;
  // Bindings to f330

  // f332
  logic [0:0] f332_wen;
  logic [31:0] f332_wdata;
  logic [0:0] f332_clk;
  logic [0:0] f332_rst;
  logic [31:0] f332_rdata;
  sr_buffer_32_1 f332(.wen(f332_wen), .wdata(f332_wdata), .clk(f332_clk), .rst(f332_rst), .rdata(f332_rdata));
  assign f332_clk = clk;
  assign f332_rst = rst;
  // Bindings to f332

  // f334
  logic [0:0] f334_wen;
  logic [31:0] f334_wdata;
  logic [0:0] f334_clk;
  logic [0:0] f334_rst;
  logic [31:0] f334_rdata;
  sr_buffer_32_1 f334(.wen(f334_wen), .wdata(f334_wdata), .clk(f334_clk), .rst(f334_rst), .rdata(f334_rdata));
  assign f334_clk = clk;
  assign f334_rst = rst;
  // Bindings to f334

  // f336
  logic [0:0] f336_wen;
  logic [31:0] f336_wdata;
  logic [0:0] f336_clk;
  logic [0:0] f336_rst;
  logic [31:0] f336_rdata;
  sr_buffer_32_1 f336(.wen(f336_wen), .wdata(f336_wdata), .clk(f336_clk), .rst(f336_rst), .rdata(f336_rdata));
  assign f336_clk = clk;
  assign f336_rst = rst;
  // Bindings to f336

  // f338
  logic [0:0] f338_wen;
  logic [31:0] f338_wdata;
  logic [0:0] f338_clk;
  logic [0:0] f338_rst;
  logic [31:0] f338_rdata;
  sr_buffer_32_1 f338(.wen(f338_wen), .wdata(f338_wdata), .clk(f338_clk), .rst(f338_rst), .rdata(f338_rdata));
  assign f338_clk = clk;
  assign f338_rst = rst;
  // Bindings to f338

  // f340
  logic [0:0] f340_wen;
  logic [31:0] f340_wdata;
  logic [0:0] f340_clk;
  logic [0:0] f340_rst;
  logic [31:0] f340_rdata;
  sr_buffer_32_1 f340(.wen(f340_wen), .wdata(f340_wdata), .clk(f340_clk), .rst(f340_rst), .rdata(f340_rdata));
  assign f340_clk = clk;
  assign f340_rst = rst;
  // Bindings to f340

  // f342
  logic [0:0] f342_wen;
  logic [31:0] f342_wdata;
  logic [0:0] f342_clk;
  logic [0:0] f342_rst;
  logic [31:0] f342_rdata;
  sr_buffer_32_1 f342(.wen(f342_wen), .wdata(f342_wdata), .clk(f342_clk), .rst(f342_rst), .rdata(f342_rdata));
  assign f342_clk = clk;
  assign f342_rst = rst;
  // Bindings to f342

  // f344
  logic [0:0] f344_wen;
  logic [31:0] f344_wdata;
  logic [0:0] f344_clk;
  logic [0:0] f344_rst;
  logic [31:0] f344_rdata;
  sr_buffer_32_1 f344(.wen(f344_wen), .wdata(f344_wdata), .clk(f344_clk), .rst(f344_rst), .rdata(f344_rdata));
  assign f344_clk = clk;
  assign f344_rst = rst;
  // Bindings to f344

  // f346
  logic [0:0] f346_wen;
  logic [31:0] f346_wdata;
  logic [0:0] f346_clk;
  logic [0:0] f346_rst;
  logic [31:0] f346_rdata;
  sr_buffer_32_1 f346(.wen(f346_wen), .wdata(f346_wdata), .clk(f346_clk), .rst(f346_rst), .rdata(f346_rdata));
  assign f346_clk = clk;
  assign f346_rst = rst;
  // Bindings to f346

  // f348
  logic [0:0] f348_wen;
  logic [31:0] f348_wdata;
  logic [0:0] f348_clk;
  logic [0:0] f348_rst;
  logic [31:0] f348_rdata;
  sr_buffer_32_1 f348(.wen(f348_wen), .wdata(f348_wdata), .clk(f348_clk), .rst(f348_rst), .rdata(f348_rdata));
  assign f348_clk = clk;
  assign f348_rst = rst;
  // Bindings to f348

  // f350
  logic [0:0] f350_wen;
  logic [31:0] f350_wdata;
  logic [0:0] f350_clk;
  logic [0:0] f350_rst;
  logic [31:0] f350_rdata;
  sr_buffer_32_1 f350(.wen(f350_wen), .wdata(f350_wdata), .clk(f350_clk), .rst(f350_rst), .rdata(f350_rdata));
  assign f350_clk = clk;
  assign f350_rst = rst;
  // Bindings to f350

  // f352
  logic [0:0] f352_wen;
  logic [31:0] f352_wdata;
  logic [0:0] f352_clk;
  logic [0:0] f352_rst;
  logic [31:0] f352_rdata;
  sr_buffer_32_1 f352(.wen(f352_wen), .wdata(f352_wdata), .clk(f352_clk), .rst(f352_rst), .rdata(f352_rdata));
  assign f352_clk = clk;
  assign f352_rst = rst;
  // Bindings to f352

  // f354
  logic [0:0] f354_wen;
  logic [31:0] f354_wdata;
  logic [0:0] f354_clk;
  logic [0:0] f354_rst;
  logic [31:0] f354_rdata;
  sr_buffer_32_1 f354(.wen(f354_wen), .wdata(f354_wdata), .clk(f354_clk), .rst(f354_rst), .rdata(f354_rdata));
  assign f354_clk = clk;
  assign f354_rst = rst;
  // Bindings to f354

  // f356
  logic [0:0] f356_wen;
  logic [31:0] f356_wdata;
  logic [0:0] f356_clk;
  logic [0:0] f356_rst;
  logic [31:0] f356_rdata;
  sr_buffer_32_1 f356(.wen(f356_wen), .wdata(f356_wdata), .clk(f356_clk), .rst(f356_rst), .rdata(f356_rdata));
  assign f356_clk = clk;
  assign f356_rst = rst;
  // Bindings to f356

  // f358
  logic [0:0] f358_wen;
  logic [31:0] f358_wdata;
  logic [0:0] f358_clk;
  logic [0:0] f358_rst;
  logic [31:0] f358_rdata;
  sr_buffer_32_1 f358(.wen(f358_wen), .wdata(f358_wdata), .clk(f358_clk), .rst(f358_rst), .rdata(f358_rdata));
  assign f358_clk = clk;
  assign f358_rst = rst;
  // Bindings to f358

  // f360
  logic [0:0] f360_wen;
  logic [31:0] f360_wdata;
  logic [0:0] f360_clk;
  logic [0:0] f360_rst;
  logic [31:0] f360_rdata;
  sr_buffer_32_1 f360(.wen(f360_wen), .wdata(f360_wdata), .clk(f360_clk), .rst(f360_rst), .rdata(f360_rdata));
  assign f360_clk = clk;
  assign f360_rst = rst;
  // Bindings to f360

  // f362
  logic [0:0] f362_wen;
  logic [31:0] f362_wdata;
  logic [0:0] f362_clk;
  logic [0:0] f362_rst;
  logic [31:0] f362_rdata;
  sr_buffer_32_1 f362(.wen(f362_wen), .wdata(f362_wdata), .clk(f362_clk), .rst(f362_rst), .rdata(f362_rdata));
  assign f362_clk = clk;
  assign f362_rst = rst;
  // Bindings to f362

  // f364
  logic [0:0] f364_wen;
  logic [31:0] f364_wdata;
  logic [0:0] f364_clk;
  logic [0:0] f364_rst;
  logic [31:0] f364_rdata;
  sr_buffer_32_1 f364(.wen(f364_wen), .wdata(f364_wdata), .clk(f364_clk), .rst(f364_rst), .rdata(f364_rdata));
  assign f364_clk = clk;
  assign f364_rst = rst;
  // Bindings to f364

  // f366
  logic [0:0] f366_wen;
  logic [31:0] f366_wdata;
  logic [0:0] f366_clk;
  logic [0:0] f366_rst;
  logic [31:0] f366_rdata;
  sr_buffer_32_1 f366(.wen(f366_wen), .wdata(f366_wdata), .clk(f366_clk), .rst(f366_rst), .rdata(f366_rdata));
  assign f366_clk = clk;
  assign f366_rst = rst;
  // Bindings to f366

  // f368
  logic [0:0] f368_wen;
  logic [31:0] f368_wdata;
  logic [0:0] f368_clk;
  logic [0:0] f368_rst;
  logic [31:0] f368_rdata;
  sr_buffer_32_1 f368(.wen(f368_wen), .wdata(f368_wdata), .clk(f368_clk), .rst(f368_rst), .rdata(f368_rdata));
  assign f368_clk = clk;
  assign f368_rst = rst;
  // Bindings to f368

  // f370
  logic [0:0] f370_wen;
  logic [31:0] f370_wdata;
  logic [0:0] f370_clk;
  logic [0:0] f370_rst;
  logic [31:0] f370_rdata;
  sr_buffer_32_1 f370(.wen(f370_wen), .wdata(f370_wdata), .clk(f370_clk), .rst(f370_rst), .rdata(f370_rdata));
  assign f370_clk = clk;
  assign f370_rst = rst;
  // Bindings to f370

  // f372
  logic [0:0] f372_wen;
  logic [31:0] f372_wdata;
  logic [0:0] f372_clk;
  logic [0:0] f372_rst;
  logic [31:0] f372_rdata;
  sr_buffer_32_1 f372(.wen(f372_wen), .wdata(f372_wdata), .clk(f372_clk), .rst(f372_rst), .rdata(f372_rdata));
  assign f372_clk = clk;
  assign f372_rst = rst;
  // Bindings to f372

  // f374
  logic [0:0] f374_wen;
  logic [31:0] f374_wdata;
  logic [0:0] f374_clk;
  logic [0:0] f374_rst;
  logic [31:0] f374_rdata;
  sr_buffer_32_1 f374(.wen(f374_wen), .wdata(f374_wdata), .clk(f374_clk), .rst(f374_rst), .rdata(f374_rdata));
  assign f374_clk = clk;
  assign f374_rst = rst;
  // Bindings to f374

  // f376
  logic [0:0] f376_wen;
  logic [31:0] f376_wdata;
  logic [0:0] f376_clk;
  logic [0:0] f376_rst;
  logic [31:0] f376_rdata;
  sr_buffer_32_1 f376(.wen(f376_wen), .wdata(f376_wdata), .clk(f376_clk), .rst(f376_rst), .rdata(f376_rdata));
  assign f376_clk = clk;
  assign f376_rst = rst;
  // Bindings to f376

  // f378
  logic [0:0] f378_wen;
  logic [31:0] f378_wdata;
  logic [0:0] f378_clk;
  logic [0:0] f378_rst;
  logic [31:0] f378_rdata;
  sr_buffer_32_1 f378(.wen(f378_wen), .wdata(f378_wdata), .clk(f378_clk), .rst(f378_rst), .rdata(f378_rdata));
  assign f378_clk = clk;
  assign f378_rst = rst;
  // Bindings to f378

  // f380
  logic [0:0] f380_wen;
  logic [31:0] f380_wdata;
  logic [0:0] f380_clk;
  logic [0:0] f380_rst;
  logic [31:0] f380_rdata;
  sr_buffer_32_1 f380(.wen(f380_wen), .wdata(f380_wdata), .clk(f380_clk), .rst(f380_rst), .rdata(f380_rdata));
  assign f380_clk = clk;
  assign f380_rst = rst;
  // Bindings to f380

  // f382
  logic [0:0] f382_wen;
  logic [31:0] f382_wdata;
  logic [0:0] f382_clk;
  logic [0:0] f382_rst;
  logic [31:0] f382_rdata;
  sr_buffer_32_1 f382(.wen(f382_wen), .wdata(f382_wdata), .clk(f382_clk), .rst(f382_rst), .rdata(f382_rdata));
  assign f382_clk = clk;
  assign f382_rst = rst;
  // Bindings to f382

  // f384
  logic [0:0] f384_wen;
  logic [31:0] f384_wdata;
  logic [0:0] f384_clk;
  logic [0:0] f384_rst;
  logic [31:0] f384_rdata;
  sr_buffer_32_1 f384(.wen(f384_wen), .wdata(f384_wdata), .clk(f384_clk), .rst(f384_rst), .rdata(f384_rdata));
  assign f384_clk = clk;
  assign f384_rst = rst;
  // Bindings to f384

  // f386
  logic [0:0] f386_wen;
  logic [31:0] f386_wdata;
  logic [0:0] f386_clk;
  logic [0:0] f386_rst;
  logic [31:0] f386_rdata;
  sr_buffer_32_1 f386(.wen(f386_wen), .wdata(f386_wdata), .clk(f386_clk), .rst(f386_rst), .rdata(f386_rdata));
  assign f386_clk = clk;
  assign f386_rst = rst;
  // Bindings to f386

  // f388
  logic [0:0] f388_wen;
  logic [31:0] f388_wdata;
  logic [0:0] f388_clk;
  logic [0:0] f388_rst;
  logic [31:0] f388_rdata;
  sr_buffer_32_1 f388(.wen(f388_wen), .wdata(f388_wdata), .clk(f388_clk), .rst(f388_rst), .rdata(f388_rdata));
  assign f388_clk = clk;
  assign f388_rst = rst;
  // Bindings to f388

  // f390
  logic [0:0] f390_wen;
  logic [31:0] f390_wdata;
  logic [0:0] f390_clk;
  logic [0:0] f390_rst;
  logic [31:0] f390_rdata;
  sr_buffer_32_1 f390(.wen(f390_wen), .wdata(f390_wdata), .clk(f390_clk), .rst(f390_rst), .rdata(f390_rdata));
  assign f390_clk = clk;
  assign f390_rst = rst;
  // Bindings to f390

  // f392
  logic [0:0] f392_wen;
  logic [31:0] f392_wdata;
  logic [0:0] f392_clk;
  logic [0:0] f392_rst;
  logic [31:0] f392_rdata;
  sr_buffer_32_1 f392(.wen(f392_wen), .wdata(f392_wdata), .clk(f392_clk), .rst(f392_rst), .rdata(f392_rdata));
  assign f392_clk = clk;
  assign f392_rst = rst;
  // Bindings to f392

  // f394
  logic [0:0] f394_wen;
  logic [31:0] f394_wdata;
  logic [0:0] f394_clk;
  logic [0:0] f394_rst;
  logic [31:0] f394_rdata;
  sr_buffer_32_1 f394(.wen(f394_wen), .wdata(f394_wdata), .clk(f394_clk), .rst(f394_rst), .rdata(f394_rdata));
  assign f394_clk = clk;
  assign f394_rst = rst;
  // Bindings to f394

  // f396
  logic [0:0] f396_wen;
  logic [31:0] f396_wdata;
  logic [0:0] f396_clk;
  logic [0:0] f396_rst;
  logic [31:0] f396_rdata;
  sr_buffer_32_1 f396(.wen(f396_wen), .wdata(f396_wdata), .clk(f396_clk), .rst(f396_rst), .rdata(f396_rdata));
  assign f396_clk = clk;
  assign f396_rst = rst;
  // Bindings to f396

  // f398
  logic [0:0] f398_wen;
  logic [31:0] f398_wdata;
  logic [0:0] f398_clk;
  logic [0:0] f398_rst;
  logic [31:0] f398_rdata;
  sr_buffer_32_1 f398(.wen(f398_wen), .wdata(f398_wdata), .clk(f398_clk), .rst(f398_rst), .rdata(f398_rdata));
  assign f398_clk = clk;
  assign f398_rst = rst;
  // Bindings to f398

  // f400
  logic [0:0] f400_wen;
  logic [31:0] f400_wdata;
  logic [0:0] f400_clk;
  logic [0:0] f400_rst;
  logic [31:0] f400_rdata;
  sr_buffer_32_1 f400(.wen(f400_wen), .wdata(f400_wdata), .clk(f400_clk), .rst(f400_rst), .rdata(f400_rdata));
  assign f400_clk = clk;
  assign f400_rst = rst;
  // Bindings to f400

  // f402
  logic [0:0] f402_wen;
  logic [31:0] f402_wdata;
  logic [0:0] f402_clk;
  logic [0:0] f402_rst;
  logic [31:0] f402_rdata;
  sr_buffer_32_1 f402(.wen(f402_wen), .wdata(f402_wdata), .clk(f402_clk), .rst(f402_rst), .rdata(f402_rdata));
  assign f402_clk = clk;
  assign f402_rst = rst;
  // Bindings to f402

  // f404
  logic [0:0] f404_wen;
  logic [31:0] f404_wdata;
  logic [0:0] f404_clk;
  logic [0:0] f404_rst;
  logic [31:0] f404_rdata;
  sr_buffer_32_1 f404(.wen(f404_wen), .wdata(f404_wdata), .clk(f404_clk), .rst(f404_rst), .rdata(f404_rdata));
  assign f404_clk = clk;
  assign f404_rst = rst;
  // Bindings to f404

  // f406
  logic [0:0] f406_wen;
  logic [31:0] f406_wdata;
  logic [0:0] f406_clk;
  logic [0:0] f406_rst;
  logic [31:0] f406_rdata;
  sr_buffer_32_1 f406(.wen(f406_wen), .wdata(f406_wdata), .clk(f406_clk), .rst(f406_rst), .rdata(f406_rdata));
  assign f406_clk = clk;
  assign f406_rst = rst;
  // Bindings to f406

  // f408
  logic [0:0] f408_wen;
  logic [31:0] f408_wdata;
  logic [0:0] f408_clk;
  logic [0:0] f408_rst;
  logic [31:0] f408_rdata;
  sr_buffer_32_1 f408(.wen(f408_wen), .wdata(f408_wdata), .clk(f408_clk), .rst(f408_rst), .rdata(f408_rdata));
  assign f408_clk = clk;
  assign f408_rst = rst;
  // Bindings to f408

  // f410
  logic [0:0] f410_wen;
  logic [31:0] f410_wdata;
  logic [0:0] f410_clk;
  logic [0:0] f410_rst;
  logic [31:0] f410_rdata;
  sr_buffer_32_1 f410(.wen(f410_wen), .wdata(f410_wdata), .clk(f410_clk), .rst(f410_rst), .rdata(f410_rdata));
  assign f410_clk = clk;
  assign f410_rst = rst;
  // Bindings to f410

  // f412
  logic [0:0] f412_wen;
  logic [31:0] f412_wdata;
  logic [0:0] f412_clk;
  logic [0:0] f412_rst;
  logic [31:0] f412_rdata;
  sr_buffer_32_1 f412(.wen(f412_wen), .wdata(f412_wdata), .clk(f412_clk), .rst(f412_rst), .rdata(f412_rdata));
  assign f412_clk = clk;
  assign f412_rst = rst;
  // Bindings to f412

  // f414
  logic [0:0] f414_wen;
  logic [31:0] f414_wdata;
  logic [0:0] f414_clk;
  logic [0:0] f414_rst;
  logic [31:0] f414_rdata;
  sr_buffer_32_1 f414(.wen(f414_wen), .wdata(f414_wdata), .clk(f414_clk), .rst(f414_rst), .rdata(f414_rdata));
  assign f414_clk = clk;
  assign f414_rst = rst;
  // Bindings to f414

  // f416
  logic [0:0] f416_wen;
  logic [31:0] f416_wdata;
  logic [0:0] f416_clk;
  logic [0:0] f416_rst;
  logic [31:0] f416_rdata;
  sr_buffer_32_1 f416(.wen(f416_wen), .wdata(f416_wdata), .clk(f416_clk), .rst(f416_rst), .rdata(f416_rdata));
  assign f416_clk = clk;
  assign f416_rst = rst;
  // Bindings to f416

  // f418
  logic [0:0] f418_wen;
  logic [31:0] f418_wdata;
  logic [0:0] f418_clk;
  logic [0:0] f418_rst;
  logic [31:0] f418_rdata;
  sr_buffer_32_1 f418(.wen(f418_wen), .wdata(f418_wdata), .clk(f418_clk), .rst(f418_rst), .rdata(f418_rdata));
  assign f418_clk = clk;
  assign f418_rst = rst;
  // Bindings to f418

  // f420
  logic [0:0] f420_wen;
  logic [31:0] f420_wdata;
  logic [0:0] f420_clk;
  logic [0:0] f420_rst;
  logic [31:0] f420_rdata;
  sr_buffer_32_1 f420(.wen(f420_wen), .wdata(f420_wdata), .clk(f420_clk), .rst(f420_rst), .rdata(f420_rdata));
  assign f420_clk = clk;
  assign f420_rst = rst;
  // Bindings to f420

  // f422
  logic [0:0] f422_wen;
  logic [31:0] f422_wdata;
  logic [0:0] f422_clk;
  logic [0:0] f422_rst;
  logic [31:0] f422_rdata;
  sr_buffer_32_1 f422(.wen(f422_wen), .wdata(f422_wdata), .clk(f422_clk), .rst(f422_rst), .rdata(f422_rdata));
  assign f422_clk = clk;
  assign f422_rst = rst;
  // Bindings to f422

  // f424
  logic [0:0] f424_wen;
  logic [31:0] f424_wdata;
  logic [0:0] f424_clk;
  logic [0:0] f424_rst;
  logic [31:0] f424_rdata;
  sr_buffer_32_1 f424(.wen(f424_wen), .wdata(f424_wdata), .clk(f424_clk), .rst(f424_rst), .rdata(f424_rdata));
  assign f424_clk = clk;
  assign f424_rst = rst;
  // Bindings to f424

  // f426
  logic [0:0] f426_wen;
  logic [31:0] f426_wdata;
  logic [0:0] f426_clk;
  logic [0:0] f426_rst;
  logic [31:0] f426_rdata;
  sr_buffer_32_1 f426(.wen(f426_wen), .wdata(f426_wdata), .clk(f426_clk), .rst(f426_rst), .rdata(f426_rdata));
  assign f426_clk = clk;
  assign f426_rst = rst;
  // Bindings to f426

  // f428
  logic [0:0] f428_wen;
  logic [31:0] f428_wdata;
  logic [0:0] f428_clk;
  logic [0:0] f428_rst;
  logic [31:0] f428_rdata;
  sr_buffer_32_1 f428(.wen(f428_wen), .wdata(f428_wdata), .clk(f428_clk), .rst(f428_rst), .rdata(f428_rdata));
  assign f428_clk = clk;
  assign f428_rst = rst;
  // Bindings to f428

  // f430
  logic [0:0] f430_wen;
  logic [31:0] f430_wdata;
  logic [0:0] f430_clk;
  logic [0:0] f430_rst;
  logic [31:0] f430_rdata;
  sr_buffer_32_1 f430(.wen(f430_wen), .wdata(f430_wdata), .clk(f430_clk), .rst(f430_rst), .rdata(f430_rdata));
  assign f430_clk = clk;
  assign f430_rst = rst;
  // Bindings to f430

  // f432
  logic [0:0] f432_wen;
  logic [31:0] f432_wdata;
  logic [0:0] f432_clk;
  logic [0:0] f432_rst;
  logic [31:0] f432_rdata;
  sr_buffer_32_1 f432(.wen(f432_wen), .wdata(f432_wdata), .clk(f432_clk), .rst(f432_rst), .rdata(f432_rdata));
  assign f432_clk = clk;
  assign f432_rst = rst;
  // Bindings to f432

  // f434
  logic [0:0] f434_wen;
  logic [31:0] f434_wdata;
  logic [0:0] f434_clk;
  logic [0:0] f434_rst;
  logic [31:0] f434_rdata;
  sr_buffer_32_1 f434(.wen(f434_wen), .wdata(f434_wdata), .clk(f434_clk), .rst(f434_rst), .rdata(f434_rdata));
  assign f434_clk = clk;
  assign f434_rst = rst;
  // Bindings to f434

  // f436
  logic [0:0] f436_wen;
  logic [31:0] f436_wdata;
  logic [0:0] f436_clk;
  logic [0:0] f436_rst;
  logic [31:0] f436_rdata;
  sr_buffer_32_1 f436(.wen(f436_wen), .wdata(f436_wdata), .clk(f436_clk), .rst(f436_rst), .rdata(f436_rdata));
  assign f436_clk = clk;
  assign f436_rst = rst;
  // Bindings to f436

  // f438
  logic [0:0] f438_wen;
  logic [31:0] f438_wdata;
  logic [0:0] f438_clk;
  logic [0:0] f438_rst;
  logic [31:0] f438_rdata;
  sr_buffer_32_1 f438(.wen(f438_wen), .wdata(f438_wdata), .clk(f438_clk), .rst(f438_rst), .rdata(f438_rdata));
  assign f438_clk = clk;
  assign f438_rst = rst;
  // Bindings to f438

  // f440
  logic [0:0] f440_wen;
  logic [31:0] f440_wdata;
  logic [0:0] f440_clk;
  logic [0:0] f440_rst;
  logic [31:0] f440_rdata;
  sr_buffer_32_1 f440(.wen(f440_wen), .wdata(f440_wdata), .clk(f440_clk), .rst(f440_rst), .rdata(f440_rdata));
  assign f440_clk = clk;
  assign f440_rst = rst;
  // Bindings to f440

  // f442
  logic [0:0] f442_wen;
  logic [31:0] f442_wdata;
  logic [0:0] f442_clk;
  logic [0:0] f442_rst;
  logic [31:0] f442_rdata;
  sr_buffer_32_1 f442(.wen(f442_wen), .wdata(f442_wdata), .clk(f442_clk), .rst(f442_rst), .rdata(f442_rdata));
  assign f442_clk = clk;
  assign f442_rst = rst;
  // Bindings to f442

  // f444
  logic [0:0] f444_wen;
  logic [31:0] f444_wdata;
  logic [0:0] f444_clk;
  logic [0:0] f444_rst;
  logic [31:0] f444_rdata;
  sr_buffer_32_1 f444(.wen(f444_wen), .wdata(f444_wdata), .clk(f444_clk), .rst(f444_rst), .rdata(f444_rdata));
  assign f444_clk = clk;
  assign f444_rst = rst;
  // Bindings to f444

  // f446
  logic [0:0] f446_wen;
  logic [31:0] f446_wdata;
  logic [0:0] f446_clk;
  logic [0:0] f446_rst;
  logic [31:0] f446_rdata;
  sr_buffer_32_1 f446(.wen(f446_wen), .wdata(f446_wdata), .clk(f446_clk), .rst(f446_rst), .rdata(f446_rdata));
  assign f446_clk = clk;
  assign f446_rst = rst;
  // Bindings to f446

  // f448
  logic [0:0] f448_wen;
  logic [31:0] f448_wdata;
  logic [0:0] f448_clk;
  logic [0:0] f448_rst;
  logic [31:0] f448_rdata;
  sr_buffer_32_1 f448(.wen(f448_wen), .wdata(f448_wdata), .clk(f448_clk), .rst(f448_rst), .rdata(f448_rdata));
  assign f448_clk = clk;
  assign f448_rst = rst;
  // Bindings to f448

  // f450
  logic [0:0] f450_wen;
  logic [31:0] f450_wdata;
  logic [0:0] f450_clk;
  logic [0:0] f450_rst;
  logic [31:0] f450_rdata;
  sr_buffer_32_1 f450(.wen(f450_wen), .wdata(f450_wdata), .clk(f450_clk), .rst(f450_rst), .rdata(f450_rdata));
  assign f450_clk = clk;
  assign f450_rst = rst;
  // Bindings to f450

  // f452
  logic [0:0] f452_wen;
  logic [31:0] f452_wdata;
  logic [0:0] f452_clk;
  logic [0:0] f452_rst;
  logic [31:0] f452_rdata;
  sr_buffer_32_1 f452(.wen(f452_wen), .wdata(f452_wdata), .clk(f452_clk), .rst(f452_rst), .rdata(f452_rdata));
  assign f452_clk = clk;
  assign f452_rst = rst;
  // Bindings to f452

  // f454
  logic [0:0] f454_wen;
  logic [31:0] f454_wdata;
  logic [0:0] f454_clk;
  logic [0:0] f454_rst;
  logic [31:0] f454_rdata;
  sr_buffer_32_1 f454(.wen(f454_wen), .wdata(f454_wdata), .clk(f454_clk), .rst(f454_rst), .rdata(f454_rdata));
  assign f454_clk = clk;
  assign f454_rst = rst;
  // Bindings to f454

  // f456
  logic [0:0] f456_wen;
  logic [31:0] f456_wdata;
  logic [0:0] f456_clk;
  logic [0:0] f456_rst;
  logic [31:0] f456_rdata;
  sr_buffer_32_1 f456(.wen(f456_wen), .wdata(f456_wdata), .clk(f456_clk), .rst(f456_rst), .rdata(f456_rdata));
  assign f456_clk = clk;
  assign f456_rst = rst;
  // Bindings to f456

  // f458
  logic [0:0] f458_wen;
  logic [31:0] f458_wdata;
  logic [0:0] f458_clk;
  logic [0:0] f458_rst;
  logic [31:0] f458_rdata;
  sr_buffer_32_1 f458(.wen(f458_wen), .wdata(f458_wdata), .clk(f458_clk), .rst(f458_rst), .rdata(f458_rdata));
  assign f458_clk = clk;
  assign f458_rst = rst;
  // Bindings to f458

  // f460
  logic [0:0] f460_wen;
  logic [31:0] f460_wdata;
  logic [0:0] f460_clk;
  logic [0:0] f460_rst;
  logic [31:0] f460_rdata;
  sr_buffer_32_1 f460(.wen(f460_wen), .wdata(f460_wdata), .clk(f460_clk), .rst(f460_rst), .rdata(f460_rdata));
  assign f460_clk = clk;
  assign f460_rst = rst;
  // Bindings to f460

  // f462
  logic [0:0] f462_wen;
  logic [31:0] f462_wdata;
  logic [0:0] f462_clk;
  logic [0:0] f462_rst;
  logic [31:0] f462_rdata;
  sr_buffer_32_1 f462(.wen(f462_wen), .wdata(f462_wdata), .clk(f462_clk), .rst(f462_rst), .rdata(f462_rdata));
  assign f462_clk = clk;
  assign f462_rst = rst;
  // Bindings to f462

  // f464
  logic [0:0] f464_wen;
  logic [31:0] f464_wdata;
  logic [0:0] f464_clk;
  logic [0:0] f464_rst;
  logic [31:0] f464_rdata;
  sr_buffer_32_1 f464(.wen(f464_wen), .wdata(f464_wdata), .clk(f464_clk), .rst(f464_rst), .rdata(f464_rdata));
  assign f464_clk = clk;
  assign f464_rst = rst;
  // Bindings to f464

  // f466
  logic [0:0] f466_wen;
  logic [31:0] f466_wdata;
  logic [0:0] f466_clk;
  logic [0:0] f466_rst;
  logic [31:0] f466_rdata;
  sr_buffer_32_1 f466(.wen(f466_wen), .wdata(f466_wdata), .clk(f466_clk), .rst(f466_rst), .rdata(f466_rdata));
  assign f466_clk = clk;
  assign f466_rst = rst;
  // Bindings to f466

  // f468
  logic [0:0] f468_wen;
  logic [31:0] f468_wdata;
  logic [0:0] f468_clk;
  logic [0:0] f468_rst;
  logic [31:0] f468_rdata;
  sr_buffer_32_1 f468(.wen(f468_wen), .wdata(f468_wdata), .clk(f468_clk), .rst(f468_rst), .rdata(f468_rdata));
  assign f468_clk = clk;
  assign f468_rst = rst;
  // Bindings to f468

  // f470
  logic [0:0] f470_wen;
  logic [31:0] f470_wdata;
  logic [0:0] f470_clk;
  logic [0:0] f470_rst;
  logic [31:0] f470_rdata;
  sr_buffer_32_1 f470(.wen(f470_wen), .wdata(f470_wdata), .clk(f470_clk), .rst(f470_rst), .rdata(f470_rdata));
  assign f470_clk = clk;
  assign f470_rst = rst;
  // Bindings to f470

  // f472
  logic [0:0] f472_wen;
  logic [31:0] f472_wdata;
  logic [0:0] f472_clk;
  logic [0:0] f472_rst;
  logic [31:0] f472_rdata;
  sr_buffer_32_1 f472(.wen(f472_wen), .wdata(f472_wdata), .clk(f472_clk), .rst(f472_rst), .rdata(f472_rdata));
  assign f472_clk = clk;
  assign f472_rst = rst;
  // Bindings to f472

  // f474
  logic [0:0] f474_wen;
  logic [31:0] f474_wdata;
  logic [0:0] f474_clk;
  logic [0:0] f474_rst;
  logic [31:0] f474_rdata;
  sr_buffer_32_1 f474(.wen(f474_wen), .wdata(f474_wdata), .clk(f474_clk), .rst(f474_rst), .rdata(f474_rdata));
  assign f474_clk = clk;
  assign f474_rst = rst;
  // Bindings to f474

  // f476
  logic [0:0] f476_wen;
  logic [31:0] f476_wdata;
  logic [0:0] f476_clk;
  logic [0:0] f476_rst;
  logic [31:0] f476_rdata;
  sr_buffer_32_1 f476(.wen(f476_wen), .wdata(f476_wdata), .clk(f476_clk), .rst(f476_rst), .rdata(f476_rdata));
  assign f476_clk = clk;
  assign f476_rst = rst;
  // Bindings to f476

  // f478
  logic [0:0] f478_wen;
  logic [31:0] f478_wdata;
  logic [0:0] f478_clk;
  logic [0:0] f478_rst;
  logic [31:0] f478_rdata;
  sr_buffer_32_1 f478(.wen(f478_wen), .wdata(f478_wdata), .clk(f478_clk), .rst(f478_rst), .rdata(f478_rdata));
  assign f478_clk = clk;
  assign f478_rst = rst;
  // Bindings to f478

  // f480
  logic [0:0] f480_wen;
  logic [31:0] f480_wdata;
  logic [0:0] f480_clk;
  logic [0:0] f480_rst;
  logic [31:0] f480_rdata;
  sr_buffer_32_1 f480(.wen(f480_wen), .wdata(f480_wdata), .clk(f480_clk), .rst(f480_rst), .rdata(f480_rdata));
  assign f480_clk = clk;
  assign f480_rst = rst;
  // Bindings to f480

  // f482
  logic [0:0] f482_wen;
  logic [31:0] f482_wdata;
  logic [0:0] f482_clk;
  logic [0:0] f482_rst;
  logic [31:0] f482_rdata;
  sr_buffer_32_1 f482(.wen(f482_wen), .wdata(f482_wdata), .clk(f482_clk), .rst(f482_rst), .rdata(f482_rdata));
  assign f482_clk = clk;
  assign f482_rst = rst;
  // Bindings to f482

  // f484
  logic [0:0] f484_wen;
  logic [31:0] f484_wdata;
  logic [0:0] f484_clk;
  logic [0:0] f484_rst;
  logic [31:0] f484_rdata;
  sr_buffer_32_1 f484(.wen(f484_wen), .wdata(f484_wdata), .clk(f484_clk), .rst(f484_rst), .rdata(f484_rdata));
  assign f484_clk = clk;
  assign f484_rst = rst;
  // Bindings to f484

  // f486
  logic [0:0] f486_wen;
  logic [31:0] f486_wdata;
  logic [0:0] f486_clk;
  logic [0:0] f486_rst;
  logic [31:0] f486_rdata;
  sr_buffer_32_1 f486(.wen(f486_wen), .wdata(f486_wdata), .clk(f486_clk), .rst(f486_rst), .rdata(f486_rdata));
  assign f486_clk = clk;
  assign f486_rst = rst;
  // Bindings to f486

  // f488
  logic [0:0] f488_wen;
  logic [31:0] f488_wdata;
  logic [0:0] f488_clk;
  logic [0:0] f488_rst;
  logic [31:0] f488_rdata;
  sr_buffer_32_1 f488(.wen(f488_wen), .wdata(f488_wdata), .clk(f488_clk), .rst(f488_rst), .rdata(f488_rdata));
  assign f488_clk = clk;
  assign f488_rst = rst;
  // Bindings to f488

  // f490
  logic [0:0] f490_wen;
  logic [31:0] f490_wdata;
  logic [0:0] f490_clk;
  logic [0:0] f490_rst;
  logic [31:0] f490_rdata;
  sr_buffer_32_1 f490(.wen(f490_wen), .wdata(f490_wdata), .clk(f490_clk), .rst(f490_rst), .rdata(f490_rdata));
  assign f490_clk = clk;
  assign f490_rst = rst;
  // Bindings to f490

  // f492
  logic [0:0] f492_wen;
  logic [31:0] f492_wdata;
  logic [0:0] f492_clk;
  logic [0:0] f492_rst;
  logic [31:0] f492_rdata;
  sr_buffer_32_1 f492(.wen(f492_wen), .wdata(f492_wdata), .clk(f492_clk), .rst(f492_rst), .rdata(f492_rdata));
  assign f492_clk = clk;
  assign f492_rst = rst;
  // Bindings to f492

  // f494
  logic [0:0] f494_wen;
  logic [31:0] f494_wdata;
  logic [0:0] f494_clk;
  logic [0:0] f494_rst;
  logic [31:0] f494_rdata;
  sr_buffer_32_1 f494(.wen(f494_wen), .wdata(f494_wdata), .clk(f494_clk), .rst(f494_rst), .rdata(f494_rdata));
  assign f494_clk = clk;
  assign f494_rst = rst;
  // Bindings to f494

  // f496
  logic [0:0] f496_wen;
  logic [31:0] f496_wdata;
  logic [0:0] f496_clk;
  logic [0:0] f496_rst;
  logic [31:0] f496_rdata;
  sr_buffer_32_1 f496(.wen(f496_wen), .wdata(f496_wdata), .clk(f496_clk), .rst(f496_rst), .rdata(f496_rdata));
  assign f496_clk = clk;
  assign f496_rst = rst;
  // Bindings to f496

  // f498
  logic [0:0] f498_wen;
  logic [31:0] f498_wdata;
  logic [0:0] f498_clk;
  logic [0:0] f498_rst;
  logic [31:0] f498_rdata;
  sr_buffer_32_1 f498(.wen(f498_wen), .wdata(f498_wdata), .clk(f498_clk), .rst(f498_rst), .rdata(f498_rdata));
  assign f498_clk = clk;
  assign f498_rst = rst;
  // Bindings to f498

  // f500
  logic [0:0] f500_wen;
  logic [31:0] f500_wdata;
  logic [0:0] f500_clk;
  logic [0:0] f500_rst;
  logic [31:0] f500_rdata;
  sr_buffer_32_1 f500(.wen(f500_wen), .wdata(f500_wdata), .clk(f500_clk), .rst(f500_rst), .rdata(f500_rdata));
  assign f500_clk = clk;
  assign f500_rst = rst;
  // Bindings to f500

  // f502
  logic [0:0] f502_wen;
  logic [31:0] f502_wdata;
  logic [0:0] f502_clk;
  logic [0:0] f502_rst;
  logic [31:0] f502_rdata;
  sr_buffer_32_1 f502(.wen(f502_wen), .wdata(f502_wdata), .clk(f502_clk), .rst(f502_rst), .rdata(f502_rdata));
  assign f502_clk = clk;
  assign f502_rst = rst;
  // Bindings to f502

  // f504
  logic [0:0] f504_wen;
  logic [31:0] f504_wdata;
  logic [0:0] f504_clk;
  logic [0:0] f504_rst;
  logic [31:0] f504_rdata;
  sr_buffer_32_1 f504(.wen(f504_wen), .wdata(f504_wdata), .clk(f504_clk), .rst(f504_rst), .rdata(f504_rdata));
  assign f504_clk = clk;
  assign f504_rst = rst;
  // Bindings to f504

  // f506
  logic [0:0] f506_wen;
  logic [31:0] f506_wdata;
  logic [0:0] f506_clk;
  logic [0:0] f506_rst;
  logic [31:0] f506_rdata;
  sr_buffer_32_1 f506(.wen(f506_wen), .wdata(f506_wdata), .clk(f506_clk), .rst(f506_rst), .rdata(f506_rdata));
  assign f506_clk = clk;
  assign f506_rst = rst;
  // Bindings to f506

  // f508
  logic [0:0] f508_wen;
  logic [31:0] f508_wdata;
  logic [0:0] f508_clk;
  logic [0:0] f508_rst;
  logic [31:0] f508_rdata;
  sr_buffer_32_1 f508(.wen(f508_wen), .wdata(f508_wdata), .clk(f508_clk), .rst(f508_rst), .rdata(f508_rdata));
  assign f508_clk = clk;
  assign f508_rst = rst;
  // Bindings to f508

  // f510
  logic [0:0] f510_wen;
  logic [31:0] f510_wdata;
  logic [0:0] f510_clk;
  logic [0:0] f510_rst;
  logic [31:0] f510_rdata;
  sr_buffer_32_1 f510(.wen(f510_wen), .wdata(f510_wdata), .clk(f510_clk), .rst(f510_rst), .rdata(f510_rdata));
  assign f510_clk = clk;
  assign f510_rst = rst;
  // Bindings to f510

  // f512
  logic [0:0] f512_wen;
  logic [31:0] f512_wdata;
  logic [0:0] f512_clk;
  logic [0:0] f512_rst;
  logic [31:0] f512_rdata;
  sr_buffer_32_1 f512(.wen(f512_wen), .wdata(f512_wdata), .clk(f512_clk), .rst(f512_rst), .rdata(f512_rdata));
  assign f512_clk = clk;
  assign f512_rst = rst;
  // Bindings to f512

  // f514
  logic [0:0] f514_wen;
  logic [31:0] f514_wdata;
  logic [0:0] f514_clk;
  logic [0:0] f514_rst;
  logic [31:0] f514_rdata;
  sr_buffer_32_1 f514(.wen(f514_wen), .wdata(f514_wdata), .clk(f514_clk), .rst(f514_rst), .rdata(f514_rdata));
  assign f514_clk = clk;
  assign f514_rst = rst;
  // Bindings to f514

  // f516
  logic [0:0] f516_wen;
  logic [31:0] f516_wdata;
  logic [0:0] f516_clk;
  logic [0:0] f516_rst;
  logic [31:0] f516_rdata;
  sr_buffer_32_1 f516(.wen(f516_wen), .wdata(f516_wdata), .clk(f516_clk), .rst(f516_rst), .rdata(f516_rdata));
  assign f516_clk = clk;
  assign f516_rst = rst;
  // Bindings to f516

  // f518
  logic [0:0] f518_wen;
  logic [31:0] f518_wdata;
  logic [0:0] f518_clk;
  logic [0:0] f518_rst;
  logic [31:0] f518_rdata;
  sr_buffer_32_1 f518(.wen(f518_wen), .wdata(f518_wdata), .clk(f518_clk), .rst(f518_rst), .rdata(f518_rdata));
  assign f518_clk = clk;
  assign f518_rst = rst;
  // Bindings to f518

  // f520
  logic [0:0] f520_wen;
  logic [31:0] f520_wdata;
  logic [0:0] f520_clk;
  logic [0:0] f520_rst;
  logic [31:0] f520_rdata;
  sr_buffer_32_1 f520(.wen(f520_wen), .wdata(f520_wdata), .clk(f520_clk), .rst(f520_rst), .rdata(f520_rdata));
  assign f520_clk = clk;
  assign f520_rst = rst;
  // Bindings to f520

  // f522
  logic [0:0] f522_wen;
  logic [31:0] f522_wdata;
  logic [0:0] f522_clk;
  logic [0:0] f522_rst;
  logic [31:0] f522_rdata;
  sr_buffer_32_1 f522(.wen(f522_wen), .wdata(f522_wdata), .clk(f522_clk), .rst(f522_rst), .rdata(f522_rdata));
  assign f522_clk = clk;
  assign f522_rst = rst;
  // Bindings to f522

  // f524
  logic [0:0] f524_wen;
  logic [31:0] f524_wdata;
  logic [0:0] f524_clk;
  logic [0:0] f524_rst;
  logic [31:0] f524_rdata;
  sr_buffer_32_1 f524(.wen(f524_wen), .wdata(f524_wdata), .clk(f524_clk), .rst(f524_rst), .rdata(f524_rdata));
  assign f524_clk = clk;
  assign f524_rst = rst;
  // Bindings to f524

  // f526
  logic [0:0] f526_wen;
  logic [31:0] f526_wdata;
  logic [0:0] f526_clk;
  logic [0:0] f526_rst;
  logic [31:0] f526_rdata;
  sr_buffer_32_1 f526(.wen(f526_wen), .wdata(f526_wdata), .clk(f526_clk), .rst(f526_rst), .rdata(f526_rdata));
  assign f526_clk = clk;
  assign f526_rst = rst;
  // Bindings to f526

  // f528
  logic [0:0] f528_wen;
  logic [31:0] f528_wdata;
  logic [0:0] f528_clk;
  logic [0:0] f528_rst;
  logic [31:0] f528_rdata;
  sr_buffer_32_1 f528(.wen(f528_wen), .wdata(f528_wdata), .clk(f528_clk), .rst(f528_rst), .rdata(f528_rdata));
  assign f528_clk = clk;
  assign f528_rst = rst;
  // Bindings to f528

  // f530
  logic [0:0] f530_wen;
  logic [31:0] f530_wdata;
  logic [0:0] f530_clk;
  logic [0:0] f530_rst;
  logic [31:0] f530_rdata;
  sr_buffer_32_1 f530(.wen(f530_wen), .wdata(f530_wdata), .clk(f530_clk), .rst(f530_rst), .rdata(f530_rdata));
  assign f530_clk = clk;
  assign f530_rst = rst;
  // Bindings to f530

  // f532
  logic [0:0] f532_wen;
  logic [31:0] f532_wdata;
  logic [0:0] f532_clk;
  logic [0:0] f532_rst;
  logic [31:0] f532_rdata;
  sr_buffer_32_1 f532(.wen(f532_wen), .wdata(f532_wdata), .clk(f532_clk), .rst(f532_rst), .rdata(f532_rdata));
  assign f532_clk = clk;
  assign f532_rst = rst;
  // Bindings to f532

  // f534
  logic [0:0] f534_wen;
  logic [31:0] f534_wdata;
  logic [0:0] f534_clk;
  logic [0:0] f534_rst;
  logic [31:0] f534_rdata;
  sr_buffer_32_1 f534(.wen(f534_wen), .wdata(f534_wdata), .clk(f534_clk), .rst(f534_rst), .rdata(f534_rdata));
  assign f534_clk = clk;
  assign f534_rst = rst;
  // Bindings to f534

  // f536
  logic [0:0] f536_wen;
  logic [31:0] f536_wdata;
  logic [0:0] f536_clk;
  logic [0:0] f536_rst;
  logic [31:0] f536_rdata;
  sr_buffer_32_1 f536(.wen(f536_wen), .wdata(f536_wdata), .clk(f536_clk), .rst(f536_rst), .rdata(f536_rdata));
  assign f536_clk = clk;
  assign f536_rst = rst;
  // Bindings to f536

  // f538
  logic [0:0] f538_wen;
  logic [31:0] f538_wdata;
  logic [0:0] f538_clk;
  logic [0:0] f538_rst;
  logic [31:0] f538_rdata;
  sr_buffer_32_1 f538(.wen(f538_wen), .wdata(f538_wdata), .clk(f538_clk), .rst(f538_rst), .rdata(f538_rdata));
  assign f538_clk = clk;
  assign f538_rst = rst;
  // Bindings to f538

  // f540
  logic [0:0] f540_wen;
  logic [31:0] f540_wdata;
  logic [0:0] f540_clk;
  logic [0:0] f540_rst;
  logic [31:0] f540_rdata;
  sr_buffer_32_1 f540(.wen(f540_wen), .wdata(f540_wdata), .clk(f540_clk), .rst(f540_rst), .rdata(f540_rdata));
  assign f540_clk = clk;
  assign f540_rst = rst;
  // Bindings to f540

  // f542
  logic [0:0] f542_wen;
  logic [31:0] f542_wdata;
  logic [0:0] f542_clk;
  logic [0:0] f542_rst;
  logic [31:0] f542_rdata;
  sr_buffer_32_1 f542(.wen(f542_wen), .wdata(f542_wdata), .clk(f542_clk), .rst(f542_rst), .rdata(f542_rdata));
  assign f542_clk = clk;
  assign f542_rst = rst;
  // Bindings to f542

  // f544
  logic [0:0] f544_wen;
  logic [31:0] f544_wdata;
  logic [0:0] f544_clk;
  logic [0:0] f544_rst;
  logic [31:0] f544_rdata;
  sr_buffer_32_1 f544(.wen(f544_wen), .wdata(f544_wdata), .clk(f544_clk), .rst(f544_rst), .rdata(f544_rdata));
  assign f544_clk = clk;
  assign f544_rst = rst;
  // Bindings to f544

  // f546
  logic [0:0] f546_wen;
  logic [31:0] f546_wdata;
  logic [0:0] f546_clk;
  logic [0:0] f546_rst;
  logic [31:0] f546_rdata;
  sr_buffer_32_1 f546(.wen(f546_wen), .wdata(f546_wdata), .clk(f546_clk), .rst(f546_rst), .rdata(f546_rdata));
  assign f546_clk = clk;
  assign f546_rst = rst;
  // Bindings to f546

  // f548
  logic [0:0] f548_wen;
  logic [31:0] f548_wdata;
  logic [0:0] f548_clk;
  logic [0:0] f548_rst;
  logic [31:0] f548_rdata;
  sr_buffer_32_1 f548(.wen(f548_wen), .wdata(f548_wdata), .clk(f548_clk), .rst(f548_rst), .rdata(f548_rdata));
  assign f548_clk = clk;
  assign f548_rst = rst;
  // Bindings to f548

  // f550
  logic [0:0] f550_wen;
  logic [31:0] f550_wdata;
  logic [0:0] f550_clk;
  logic [0:0] f550_rst;
  logic [31:0] f550_rdata;
  sr_buffer_32_1 f550(.wen(f550_wen), .wdata(f550_wdata), .clk(f550_clk), .rst(f550_rst), .rdata(f550_rdata));
  assign f550_clk = clk;
  assign f550_rst = rst;
  // Bindings to f550

  // f552
  logic [0:0] f552_wen;
  logic [31:0] f552_wdata;
  logic [0:0] f552_clk;
  logic [0:0] f552_rst;
  logic [31:0] f552_rdata;
  sr_buffer_32_1 f552(.wen(f552_wen), .wdata(f552_wdata), .clk(f552_clk), .rst(f552_rst), .rdata(f552_rdata));
  assign f552_clk = clk;
  assign f552_rst = rst;
  // Bindings to f552

  // f554
  logic [0:0] f554_wen;
  logic [31:0] f554_wdata;
  logic [0:0] f554_clk;
  logic [0:0] f554_rst;
  logic [31:0] f554_rdata;
  sr_buffer_32_1 f554(.wen(f554_wen), .wdata(f554_wdata), .clk(f554_clk), .rst(f554_rst), .rdata(f554_rdata));
  assign f554_clk = clk;
  assign f554_rst = rst;
  // Bindings to f554

  // f556
  logic [0:0] f556_wen;
  logic [31:0] f556_wdata;
  logic [0:0] f556_clk;
  logic [0:0] f556_rst;
  logic [31:0] f556_rdata;
  sr_buffer_32_1 f556(.wen(f556_wen), .wdata(f556_wdata), .clk(f556_clk), .rst(f556_rst), .rdata(f556_rdata));
  assign f556_clk = clk;
  assign f556_rst = rst;
  // Bindings to f556

  // f558
  logic [0:0] f558_wen;
  logic [31:0] f558_wdata;
  logic [0:0] f558_clk;
  logic [0:0] f558_rst;
  logic [31:0] f558_rdata;
  sr_buffer_32_1 f558(.wen(f558_wen), .wdata(f558_wdata), .clk(f558_clk), .rst(f558_rst), .rdata(f558_rdata));
  assign f558_clk = clk;
  assign f558_rst = rst;
  // Bindings to f558

  // f560
  logic [0:0] f560_wen;
  logic [31:0] f560_wdata;
  logic [0:0] f560_clk;
  logic [0:0] f560_rst;
  logic [31:0] f560_rdata;
  sr_buffer_32_1 f560(.wen(f560_wen), .wdata(f560_wdata), .clk(f560_clk), .rst(f560_rst), .rdata(f560_rdata));
  assign f560_clk = clk;
  assign f560_rst = rst;
  // Bindings to f560

  // f562
  logic [0:0] f562_wen;
  logic [31:0] f562_wdata;
  logic [0:0] f562_clk;
  logic [0:0] f562_rst;
  logic [31:0] f562_rdata;
  sr_buffer_32_1 f562(.wen(f562_wen), .wdata(f562_wdata), .clk(f562_clk), .rst(f562_rst), .rdata(f562_rdata));
  assign f562_clk = clk;
  assign f562_rst = rst;
  // Bindings to f562

  // f564
  logic [0:0] f564_wen;
  logic [31:0] f564_wdata;
  logic [0:0] f564_clk;
  logic [0:0] f564_rst;
  logic [31:0] f564_rdata;
  sr_buffer_32_1 f564(.wen(f564_wen), .wdata(f564_wdata), .clk(f564_clk), .rst(f564_rst), .rdata(f564_rdata));
  assign f564_clk = clk;
  assign f564_rst = rst;
  // Bindings to f564

  // f566
  logic [0:0] f566_wen;
  logic [31:0] f566_wdata;
  logic [0:0] f566_clk;
  logic [0:0] f566_rst;
  logic [31:0] f566_rdata;
  sr_buffer_32_1 f566(.wen(f566_wen), .wdata(f566_wdata), .clk(f566_clk), .rst(f566_rst), .rdata(f566_rdata));
  assign f566_clk = clk;
  assign f566_rst = rst;
  // Bindings to f566

  // f568
  logic [0:0] f568_wen;
  logic [31:0] f568_wdata;
  logic [0:0] f568_clk;
  logic [0:0] f568_rst;
  logic [31:0] f568_rdata;
  sr_buffer_32_1 f568(.wen(f568_wen), .wdata(f568_wdata), .clk(f568_clk), .rst(f568_rst), .rdata(f568_rdata));
  assign f568_clk = clk;
  assign f568_rst = rst;
  // Bindings to f568

  // f570
  logic [0:0] f570_wen;
  logic [31:0] f570_wdata;
  logic [0:0] f570_clk;
  logic [0:0] f570_rst;
  logic [31:0] f570_rdata;
  sr_buffer_32_1 f570(.wen(f570_wen), .wdata(f570_wdata), .clk(f570_clk), .rst(f570_rst), .rdata(f570_rdata));
  assign f570_clk = clk;
  assign f570_rst = rst;
  // Bindings to f570

  // f572
  logic [0:0] f572_wen;
  logic [31:0] f572_wdata;
  logic [0:0] f572_clk;
  logic [0:0] f572_rst;
  logic [31:0] f572_rdata;
  sr_buffer_32_1 f572(.wen(f572_wen), .wdata(f572_wdata), .clk(f572_clk), .rst(f572_rst), .rdata(f572_rdata));
  assign f572_clk = clk;
  assign f572_rst = rst;
  // Bindings to f572

  // f574
  logic [0:0] f574_wen;
  logic [31:0] f574_wdata;
  logic [0:0] f574_clk;
  logic [0:0] f574_rst;
  logic [31:0] f574_rdata;
  sr_buffer_32_1 f574(.wen(f574_wen), .wdata(f574_wdata), .clk(f574_clk), .rst(f574_rst), .rdata(f574_rdata));
  assign f574_clk = clk;
  assign f574_rst = rst;
  // Bindings to f574

  // f576
  logic [0:0] f576_wen;
  logic [31:0] f576_wdata;
  logic [0:0] f576_clk;
  logic [0:0] f576_rst;
  logic [31:0] f576_rdata;
  sr_buffer_32_1 f576(.wen(f576_wen), .wdata(f576_wdata), .clk(f576_clk), .rst(f576_rst), .rdata(f576_rdata));
  assign f576_clk = clk;
  assign f576_rst = rst;
  // Bindings to f576

  // f578
  logic [0:0] f578_wen;
  logic [31:0] f578_wdata;
  logic [0:0] f578_clk;
  logic [0:0] f578_rst;
  logic [31:0] f578_rdata;
  sr_buffer_32_1 f578(.wen(f578_wen), .wdata(f578_wdata), .clk(f578_clk), .rst(f578_rst), .rdata(f578_rdata));
  assign f578_clk = clk;
  assign f578_rst = rst;
  // Bindings to f578

  // f580
  logic [0:0] f580_wen;
  logic [31:0] f580_wdata;
  logic [0:0] f580_clk;
  logic [0:0] f580_rst;
  logic [31:0] f580_rdata;
  sr_buffer_32_1 f580(.wen(f580_wen), .wdata(f580_wdata), .clk(f580_clk), .rst(f580_rst), .rdata(f580_rdata));
  assign f580_clk = clk;
  assign f580_rst = rst;
  // Bindings to f580

  // f582
  logic [0:0] f582_wen;
  logic [31:0] f582_wdata;
  logic [0:0] f582_clk;
  logic [0:0] f582_rst;
  logic [31:0] f582_rdata;
  sr_buffer_32_1 f582(.wen(f582_wen), .wdata(f582_wdata), .clk(f582_clk), .rst(f582_rst), .rdata(f582_rdata));
  assign f582_clk = clk;
  assign f582_rst = rst;
  // Bindings to f582

  // f584
  logic [0:0] f584_wen;
  logic [31:0] f584_wdata;
  logic [0:0] f584_clk;
  logic [0:0] f584_rst;
  logic [31:0] f584_rdata;
  sr_buffer_32_1 f584(.wen(f584_wen), .wdata(f584_wdata), .clk(f584_clk), .rst(f584_rst), .rdata(f584_rdata));
  assign f584_clk = clk;
  assign f584_rst = rst;
  // Bindings to f584

  // f586
  logic [0:0] f586_wen;
  logic [31:0] f586_wdata;
  logic [0:0] f586_clk;
  logic [0:0] f586_rst;
  logic [31:0] f586_rdata;
  sr_buffer_32_1 f586(.wen(f586_wen), .wdata(f586_wdata), .clk(f586_clk), .rst(f586_rst), .rdata(f586_rdata));
  assign f586_clk = clk;
  assign f586_rst = rst;
  // Bindings to f586

  // f588
  logic [0:0] f588_wen;
  logic [31:0] f588_wdata;
  logic [0:0] f588_clk;
  logic [0:0] f588_rst;
  logic [31:0] f588_rdata;
  sr_buffer_32_1 f588(.wen(f588_wen), .wdata(f588_wdata), .clk(f588_clk), .rst(f588_rst), .rdata(f588_rdata));
  assign f588_clk = clk;
  assign f588_rst = rst;
  // Bindings to f588

  // f590
  logic [0:0] f590_wen;
  logic [31:0] f590_wdata;
  logic [0:0] f590_clk;
  logic [0:0] f590_rst;
  logic [31:0] f590_rdata;
  sr_buffer_32_1 f590(.wen(f590_wen), .wdata(f590_wdata), .clk(f590_clk), .rst(f590_rst), .rdata(f590_rdata));
  assign f590_clk = clk;
  assign f590_rst = rst;
  // Bindings to f590

  // f592
  logic [0:0] f592_wen;
  logic [31:0] f592_wdata;
  logic [0:0] f592_clk;
  logic [0:0] f592_rst;
  logic [31:0] f592_rdata;
  sr_buffer_32_1 f592(.wen(f592_wen), .wdata(f592_wdata), .clk(f592_clk), .rst(f592_rst), .rdata(f592_rdata));
  assign f592_clk = clk;
  assign f592_rst = rst;
  // Bindings to f592

  // f594
  logic [0:0] f594_wen;
  logic [31:0] f594_wdata;
  logic [0:0] f594_clk;
  logic [0:0] f594_rst;
  logic [31:0] f594_rdata;
  sr_buffer_32_1 f594(.wen(f594_wen), .wdata(f594_wdata), .clk(f594_clk), .rst(f594_rst), .rdata(f594_rdata));
  assign f594_clk = clk;
  assign f594_rst = rst;
  // Bindings to f594

  // f596
  logic [0:0] f596_wen;
  logic [31:0] f596_wdata;
  logic [0:0] f596_clk;
  logic [0:0] f596_rst;
  logic [31:0] f596_rdata;
  sr_buffer_32_1 f596(.wen(f596_wen), .wdata(f596_wdata), .clk(f596_clk), .rst(f596_rst), .rdata(f596_rdata));
  assign f596_clk = clk;
  assign f596_rst = rst;
  // Bindings to f596

  // f598
  logic [0:0] f598_wen;
  logic [31:0] f598_wdata;
  logic [0:0] f598_clk;
  logic [0:0] f598_rst;
  logic [31:0] f598_rdata;
  sr_buffer_32_1 f598(.wen(f598_wen), .wdata(f598_wdata), .clk(f598_clk), .rst(f598_rst), .rdata(f598_rdata));
  assign f598_clk = clk;
  assign f598_rst = rst;
  // Bindings to f598

  // f600
  logic [0:0] f600_wen;
  logic [31:0] f600_wdata;
  logic [0:0] f600_clk;
  logic [0:0] f600_rst;
  logic [31:0] f600_rdata;
  sr_buffer_32_1 f600(.wen(f600_wen), .wdata(f600_wdata), .clk(f600_clk), .rst(f600_rst), .rdata(f600_rdata));
  assign f600_clk = clk;
  assign f600_rst = rst;
  // Bindings to f600

  // f602
  logic [0:0] f602_wen;
  logic [31:0] f602_wdata;
  logic [0:0] f602_clk;
  logic [0:0] f602_rst;
  logic [31:0] f602_rdata;
  sr_buffer_32_1 f602(.wen(f602_wen), .wdata(f602_wdata), .clk(f602_clk), .rst(f602_rst), .rdata(f602_rdata));
  assign f602_clk = clk;
  assign f602_rst = rst;
  // Bindings to f602

  // f604
  logic [0:0] f604_wen;
  logic [31:0] f604_wdata;
  logic [0:0] f604_clk;
  logic [0:0] f604_rst;
  logic [31:0] f604_rdata;
  sr_buffer_32_1 f604(.wen(f604_wen), .wdata(f604_wdata), .clk(f604_clk), .rst(f604_rst), .rdata(f604_rdata));
  assign f604_clk = clk;
  assign f604_rst = rst;
  // Bindings to f604

  // f606
  logic [0:0] f606_wen;
  logic [31:0] f606_wdata;
  logic [0:0] f606_clk;
  logic [0:0] f606_rst;
  logic [31:0] f606_rdata;
  sr_buffer_32_1 f606(.wen(f606_wen), .wdata(f606_wdata), .clk(f606_clk), .rst(f606_rst), .rdata(f606_rdata));
  assign f606_clk = clk;
  assign f606_rst = rst;
  // Bindings to f606

  // f608
  logic [0:0] f608_wen;
  logic [31:0] f608_wdata;
  logic [0:0] f608_clk;
  logic [0:0] f608_rst;
  logic [31:0] f608_rdata;
  sr_buffer_32_1 f608(.wen(f608_wen), .wdata(f608_wdata), .clk(f608_clk), .rst(f608_rst), .rdata(f608_rdata));
  assign f608_clk = clk;
  assign f608_rst = rst;
  // Bindings to f608

  // f610
  logic [0:0] f610_wen;
  logic [31:0] f610_wdata;
  logic [0:0] f610_clk;
  logic [0:0] f610_rst;
  logic [31:0] f610_rdata;
  sr_buffer_32_1 f610(.wen(f610_wen), .wdata(f610_wdata), .clk(f610_clk), .rst(f610_rst), .rdata(f610_rdata));
  assign f610_clk = clk;
  assign f610_rst = rst;
  // Bindings to f610

  // f612
  logic [0:0] f612_wen;
  logic [31:0] f612_wdata;
  logic [0:0] f612_clk;
  logic [0:0] f612_rst;
  logic [31:0] f612_rdata;
  sr_buffer_32_1 f612(.wen(f612_wen), .wdata(f612_wdata), .clk(f612_clk), .rst(f612_rst), .rdata(f612_rdata));
  assign f612_clk = clk;
  assign f612_rst = rst;
  // Bindings to f612

  // f614
  logic [0:0] f614_wen;
  logic [31:0] f614_wdata;
  logic [0:0] f614_clk;
  logic [0:0] f614_rst;
  logic [31:0] f614_rdata;
  sr_buffer_32_1 f614(.wen(f614_wen), .wdata(f614_wdata), .clk(f614_clk), .rst(f614_rst), .rdata(f614_rdata));
  assign f614_clk = clk;
  assign f614_rst = rst;
  // Bindings to f614

  // f616
  logic [0:0] f616_wen;
  logic [31:0] f616_wdata;
  logic [0:0] f616_clk;
  logic [0:0] f616_rst;
  logic [31:0] f616_rdata;
  sr_buffer_32_1 f616(.wen(f616_wen), .wdata(f616_wdata), .clk(f616_clk), .rst(f616_rst), .rdata(f616_rdata));
  assign f616_clk = clk;
  assign f616_rst = rst;
  // Bindings to f616

  // f618
  logic [0:0] f618_wen;
  logic [31:0] f618_wdata;
  logic [0:0] f618_clk;
  logic [0:0] f618_rst;
  logic [31:0] f618_rdata;
  sr_buffer_32_1 f618(.wen(f618_wen), .wdata(f618_wdata), .clk(f618_clk), .rst(f618_rst), .rdata(f618_rdata));
  assign f618_clk = clk;
  assign f618_rst = rst;
  // Bindings to f618

  // f620
  logic [0:0] f620_wen;
  logic [31:0] f620_wdata;
  logic [0:0] f620_clk;
  logic [0:0] f620_rst;
  logic [31:0] f620_rdata;
  sr_buffer_32_1 f620(.wen(f620_wen), .wdata(f620_wdata), .clk(f620_clk), .rst(f620_rst), .rdata(f620_rdata));
  assign f620_clk = clk;
  assign f620_rst = rst;
  // Bindings to f620

  // f622
  logic [0:0] f622_wen;
  logic [31:0] f622_wdata;
  logic [0:0] f622_clk;
  logic [0:0] f622_rst;
  logic [31:0] f622_rdata;
  sr_buffer_32_1 f622(.wen(f622_wen), .wdata(f622_wdata), .clk(f622_clk), .rst(f622_rst), .rdata(f622_rdata));
  assign f622_clk = clk;
  assign f622_rst = rst;
  // Bindings to f622

  // f624
  logic [0:0] f624_wen;
  logic [31:0] f624_wdata;
  logic [0:0] f624_clk;
  logic [0:0] f624_rst;
  logic [31:0] f624_rdata;
  sr_buffer_32_1 f624(.wen(f624_wen), .wdata(f624_wdata), .clk(f624_clk), .rst(f624_rst), .rdata(f624_rdata));
  assign f624_clk = clk;
  assign f624_rst = rst;
  // Bindings to f624

  // f626
  logic [0:0] f626_wen;
  logic [31:0] f626_wdata;
  logic [0:0] f626_clk;
  logic [0:0] f626_rst;
  logic [31:0] f626_rdata;
  sr_buffer_32_1 f626(.wen(f626_wen), .wdata(f626_wdata), .clk(f626_clk), .rst(f626_rst), .rdata(f626_rdata));
  assign f626_clk = clk;
  assign f626_rst = rst;
  // Bindings to f626

  // f628
  logic [0:0] f628_wen;
  logic [31:0] f628_wdata;
  logic [0:0] f628_clk;
  logic [0:0] f628_rst;
  logic [31:0] f628_rdata;
  sr_buffer_32_1 f628(.wen(f628_wen), .wdata(f628_wdata), .clk(f628_clk), .rst(f628_rst), .rdata(f628_rdata));
  assign f628_clk = clk;
  assign f628_rst = rst;
  // Bindings to f628

  // f630
  logic [0:0] f630_wen;
  logic [31:0] f630_wdata;
  logic [0:0] f630_clk;
  logic [0:0] f630_rst;
  logic [31:0] f630_rdata;
  sr_buffer_32_1 f630(.wen(f630_wen), .wdata(f630_wdata), .clk(f630_clk), .rst(f630_rst), .rdata(f630_rdata));
  assign f630_clk = clk;
  assign f630_rst = rst;
  // Bindings to f630

  // f632
  logic [0:0] f632_wen;
  logic [31:0] f632_wdata;
  logic [0:0] f632_clk;
  logic [0:0] f632_rst;
  logic [31:0] f632_rdata;
  sr_buffer_32_1 f632(.wen(f632_wen), .wdata(f632_wdata), .clk(f632_clk), .rst(f632_rst), .rdata(f632_rdata));
  assign f632_clk = clk;
  assign f632_rst = rst;
  // Bindings to f632

  // f634
  logic [0:0] f634_wen;
  logic [31:0] f634_wdata;
  logic [0:0] f634_clk;
  logic [0:0] f634_rst;
  logic [31:0] f634_rdata;
  sr_buffer_32_1 f634(.wen(f634_wen), .wdata(f634_wdata), .clk(f634_clk), .rst(f634_rst), .rdata(f634_rdata));
  assign f634_clk = clk;
  assign f634_rst = rst;
  // Bindings to f634

  // f636
  logic [0:0] f636_wen;
  logic [31:0] f636_wdata;
  logic [0:0] f636_clk;
  logic [0:0] f636_rst;
  logic [31:0] f636_rdata;
  sr_buffer_32_1 f636(.wen(f636_wen), .wdata(f636_wdata), .clk(f636_clk), .rst(f636_rst), .rdata(f636_rdata));
  assign f636_clk = clk;
  assign f636_rst = rst;
  // Bindings to f636

  // f638
  logic [0:0] f638_wen;
  logic [31:0] f638_wdata;
  logic [0:0] f638_clk;
  logic [0:0] f638_rst;
  logic [31:0] f638_rdata;
  sr_buffer_32_1 f638(.wen(f638_wen), .wdata(f638_wdata), .clk(f638_clk), .rst(f638_rst), .rdata(f638_rdata));
  assign f638_clk = clk;
  assign f638_rst = rst;
  // Bindings to f638

  // f640
  logic [0:0] f640_wen;
  logic [31:0] f640_wdata;
  logic [0:0] f640_clk;
  logic [0:0] f640_rst;
  logic [31:0] f640_rdata;
  sr_buffer_32_1 f640(.wen(f640_wen), .wdata(f640_wdata), .clk(f640_clk), .rst(f640_rst), .rdata(f640_rdata));
  assign f640_clk = clk;
  assign f640_rst = rst;
  // Bindings to f640

  // f642
  logic [0:0] f642_wen;
  logic [31:0] f642_wdata;
  logic [0:0] f642_clk;
  logic [0:0] f642_rst;
  logic [31:0] f642_rdata;
  sr_buffer_32_1 f642(.wen(f642_wen), .wdata(f642_wdata), .clk(f642_clk), .rst(f642_rst), .rdata(f642_rdata));
  assign f642_clk = clk;
  assign f642_rst = rst;
  // Bindings to f642

  // f644
  logic [0:0] f644_wen;
  logic [31:0] f644_wdata;
  logic [0:0] f644_clk;
  logic [0:0] f644_rst;
  logic [31:0] f644_rdata;
  sr_buffer_32_1 f644(.wen(f644_wen), .wdata(f644_wdata), .clk(f644_clk), .rst(f644_rst), .rdata(f644_rdata));
  assign f644_clk = clk;
  assign f644_rst = rst;
  // Bindings to f644

  // f646
  logic [0:0] f646_wen;
  logic [31:0] f646_wdata;
  logic [0:0] f646_clk;
  logic [0:0] f646_rst;
  logic [31:0] f646_rdata;
  sr_buffer_32_1 f646(.wen(f646_wen), .wdata(f646_wdata), .clk(f646_clk), .rst(f646_rst), .rdata(f646_rdata));
  assign f646_clk = clk;
  assign f646_rst = rst;
  // Bindings to f646

  // f648
  logic [0:0] f648_wen;
  logic [31:0] f648_wdata;
  logic [0:0] f648_clk;
  logic [0:0] f648_rst;
  logic [31:0] f648_rdata;
  sr_buffer_32_1 f648(.wen(f648_wen), .wdata(f648_wdata), .clk(f648_clk), .rst(f648_rst), .rdata(f648_rdata));
  assign f648_clk = clk;
  assign f648_rst = rst;
  // Bindings to f648

  // f650
  logic [0:0] f650_wen;
  logic [31:0] f650_wdata;
  logic [0:0] f650_clk;
  logic [0:0] f650_rst;
  logic [31:0] f650_rdata;
  sr_buffer_32_1 f650(.wen(f650_wen), .wdata(f650_wdata), .clk(f650_clk), .rst(f650_rst), .rdata(f650_rdata));
  assign f650_clk = clk;
  assign f650_rst = rst;
  // Bindings to f650

  // f652
  logic [0:0] f652_wen;
  logic [31:0] f652_wdata;
  logic [0:0] f652_clk;
  logic [0:0] f652_rst;
  logic [31:0] f652_rdata;
  sr_buffer_32_1 f652(.wen(f652_wen), .wdata(f652_wdata), .clk(f652_clk), .rst(f652_rst), .rdata(f652_rdata));
  assign f652_clk = clk;
  assign f652_rst = rst;
  // Bindings to f652

  // f654
  logic [0:0] f654_wen;
  logic [31:0] f654_wdata;
  logic [0:0] f654_clk;
  logic [0:0] f654_rst;
  logic [31:0] f654_rdata;
  sr_buffer_32_1 f654(.wen(f654_wen), .wdata(f654_wdata), .clk(f654_clk), .rst(f654_rst), .rdata(f654_rdata));
  assign f654_clk = clk;
  assign f654_rst = rst;
  // Bindings to f654

  // f656
  logic [0:0] f656_wen;
  logic [31:0] f656_wdata;
  logic [0:0] f656_clk;
  logic [0:0] f656_rst;
  logic [31:0] f656_rdata;
  sr_buffer_32_1 f656(.wen(f656_wen), .wdata(f656_wdata), .clk(f656_clk), .rst(f656_rst), .rdata(f656_rdata));
  assign f656_clk = clk;
  assign f656_rst = rst;
  // Bindings to f656

  // f658
  logic [0:0] f658_wen;
  logic [31:0] f658_wdata;
  logic [0:0] f658_clk;
  logic [0:0] f658_rst;
  logic [31:0] f658_rdata;
  sr_buffer_32_1 f658(.wen(f658_wen), .wdata(f658_wdata), .clk(f658_clk), .rst(f658_rst), .rdata(f658_rdata));
  assign f658_clk = clk;
  assign f658_rst = rst;
  // Bindings to f658

  // f660
  logic [0:0] f660_wen;
  logic [31:0] f660_wdata;
  logic [0:0] f660_clk;
  logic [0:0] f660_rst;
  logic [31:0] f660_rdata;
  sr_buffer_32_1 f660(.wen(f660_wen), .wdata(f660_wdata), .clk(f660_clk), .rst(f660_rst), .rdata(f660_rdata));
  assign f660_clk = clk;
  assign f660_rst = rst;
  // Bindings to f660

  // f662
  logic [0:0] f662_wen;
  logic [31:0] f662_wdata;
  logic [0:0] f662_clk;
  logic [0:0] f662_rst;
  logic [31:0] f662_rdata;
  sr_buffer_32_1 f662(.wen(f662_wen), .wdata(f662_wdata), .clk(f662_clk), .rst(f662_rst), .rdata(f662_rdata));
  assign f662_clk = clk;
  assign f662_rst = rst;
  // Bindings to f662

  // f664
  logic [0:0] f664_wen;
  logic [31:0] f664_wdata;
  logic [0:0] f664_clk;
  logic [0:0] f664_rst;
  logic [31:0] f664_rdata;
  sr_buffer_32_1 f664(.wen(f664_wen), .wdata(f664_wdata), .clk(f664_clk), .rst(f664_rst), .rdata(f664_rdata));
  assign f664_clk = clk;
  assign f664_rst = rst;
  // Bindings to f664

  // f666
  logic [0:0] f666_wen;
  logic [31:0] f666_wdata;
  logic [0:0] f666_clk;
  logic [0:0] f666_rst;
  logic [31:0] f666_rdata;
  sr_buffer_32_1 f666(.wen(f666_wen), .wdata(f666_wdata), .clk(f666_clk), .rst(f666_rst), .rdata(f666_rdata));
  assign f666_clk = clk;
  assign f666_rst = rst;
  // Bindings to f666

  // f668
  logic [0:0] f668_wen;
  logic [31:0] f668_wdata;
  logic [0:0] f668_clk;
  logic [0:0] f668_rst;
  logic [31:0] f668_rdata;
  sr_buffer_32_1 f668(.wen(f668_wen), .wdata(f668_wdata), .clk(f668_clk), .rst(f668_rst), .rdata(f668_rdata));
  assign f668_clk = clk;
  assign f668_rst = rst;
  // Bindings to f668

  // f670
  logic [0:0] f670_wen;
  logic [31:0] f670_wdata;
  logic [0:0] f670_clk;
  logic [0:0] f670_rst;
  logic [31:0] f670_rdata;
  sr_buffer_32_1 f670(.wen(f670_wen), .wdata(f670_wdata), .clk(f670_clk), .rst(f670_rst), .rdata(f670_rdata));
  assign f670_clk = clk;
  assign f670_rst = rst;
  // Bindings to f670

  // f672
  logic [0:0] f672_wen;
  logic [31:0] f672_wdata;
  logic [0:0] f672_clk;
  logic [0:0] f672_rst;
  logic [31:0] f672_rdata;
  sr_buffer_32_1 f672(.wen(f672_wen), .wdata(f672_wdata), .clk(f672_clk), .rst(f672_rst), .rdata(f672_rdata));
  assign f672_clk = clk;
  assign f672_rst = rst;
  // Bindings to f672

  // f674
  logic [0:0] f674_wen;
  logic [31:0] f674_wdata;
  logic [0:0] f674_clk;
  logic [0:0] f674_rst;
  logic [31:0] f674_rdata;
  sr_buffer_32_1 f674(.wen(f674_wen), .wdata(f674_wdata), .clk(f674_clk), .rst(f674_rst), .rdata(f674_rdata));
  assign f674_clk = clk;
  assign f674_rst = rst;
  // Bindings to f674

  // f676
  logic [0:0] f676_wen;
  logic [31:0] f676_wdata;
  logic [0:0] f676_clk;
  logic [0:0] f676_rst;
  logic [31:0] f676_rdata;
  sr_buffer_32_1 f676(.wen(f676_wen), .wdata(f676_wdata), .clk(f676_clk), .rst(f676_rst), .rdata(f676_rdata));
  assign f676_clk = clk;
  assign f676_rst = rst;
  // Bindings to f676

  // f678
  logic [0:0] f678_wen;
  logic [31:0] f678_wdata;
  logic [0:0] f678_clk;
  logic [0:0] f678_rst;
  logic [31:0] f678_rdata;
  sr_buffer_32_1 f678(.wen(f678_wen), .wdata(f678_wdata), .clk(f678_clk), .rst(f678_rst), .rdata(f678_rdata));
  assign f678_clk = clk;
  assign f678_rst = rst;
  // Bindings to f678

  // f680
  logic [0:0] f680_wen;
  logic [31:0] f680_wdata;
  logic [0:0] f680_clk;
  logic [0:0] f680_rst;
  logic [31:0] f680_rdata;
  sr_buffer_32_1 f680(.wen(f680_wen), .wdata(f680_wdata), .clk(f680_clk), .rst(f680_rst), .rdata(f680_rdata));
  assign f680_clk = clk;
  assign f680_rst = rst;
  // Bindings to f680

  // f682
  logic [0:0] f682_wen;
  logic [31:0] f682_wdata;
  logic [0:0] f682_clk;
  logic [0:0] f682_rst;
  logic [31:0] f682_rdata;
  sr_buffer_32_1 f682(.wen(f682_wen), .wdata(f682_wdata), .clk(f682_clk), .rst(f682_rst), .rdata(f682_rdata));
  assign f682_clk = clk;
  assign f682_rst = rst;
  // Bindings to f682

  // f684
  logic [0:0] f684_wen;
  logic [31:0] f684_wdata;
  logic [0:0] f684_clk;
  logic [0:0] f684_rst;
  logic [31:0] f684_rdata;
  sr_buffer_32_1 f684(.wen(f684_wen), .wdata(f684_wdata), .clk(f684_clk), .rst(f684_rst), .rdata(f684_rdata));
  assign f684_clk = clk;
  assign f684_rst = rst;
  // Bindings to f684

  // f686
  logic [0:0] f686_wen;
  logic [31:0] f686_wdata;
  logic [0:0] f686_clk;
  logic [0:0] f686_rst;
  logic [31:0] f686_rdata;
  sr_buffer_32_1 f686(.wen(f686_wen), .wdata(f686_wdata), .clk(f686_clk), .rst(f686_rst), .rdata(f686_rdata));
  assign f686_clk = clk;
  assign f686_rst = rst;
  // Bindings to f686

  // f688
  logic [0:0] f688_wen;
  logic [31:0] f688_wdata;
  logic [0:0] f688_clk;
  logic [0:0] f688_rst;
  logic [31:0] f688_rdata;
  sr_buffer_32_1 f688(.wen(f688_wen), .wdata(f688_wdata), .clk(f688_clk), .rst(f688_rst), .rdata(f688_rdata));
  assign f688_clk = clk;
  assign f688_rst = rst;
  // Bindings to f688

  // f690
  logic [0:0] f690_wen;
  logic [31:0] f690_wdata;
  logic [0:0] f690_clk;
  logic [0:0] f690_rst;
  logic [31:0] f690_rdata;
  sr_buffer_32_1 f690(.wen(f690_wen), .wdata(f690_wdata), .clk(f690_clk), .rst(f690_rst), .rdata(f690_rdata));
  assign f690_clk = clk;
  assign f690_rst = rst;
  // Bindings to f690

  // f692
  logic [0:0] f692_wen;
  logic [31:0] f692_wdata;
  logic [0:0] f692_clk;
  logic [0:0] f692_rst;
  logic [31:0] f692_rdata;
  sr_buffer_32_1 f692(.wen(f692_wen), .wdata(f692_wdata), .clk(f692_clk), .rst(f692_rst), .rdata(f692_rdata));
  assign f692_clk = clk;
  assign f692_rst = rst;
  // Bindings to f692

  // f694
  logic [0:0] f694_wen;
  logic [31:0] f694_wdata;
  logic [0:0] f694_clk;
  logic [0:0] f694_rst;
  logic [31:0] f694_rdata;
  sr_buffer_32_1 f694(.wen(f694_wen), .wdata(f694_wdata), .clk(f694_clk), .rst(f694_rst), .rdata(f694_rdata));
  assign f694_clk = clk;
  assign f694_rst = rst;
  // Bindings to f694

  // f696
  logic [0:0] f696_wen;
  logic [31:0] f696_wdata;
  logic [0:0] f696_clk;
  logic [0:0] f696_rst;
  logic [31:0] f696_rdata;
  sr_buffer_32_1 f696(.wen(f696_wen), .wdata(f696_wdata), .clk(f696_clk), .rst(f696_rst), .rdata(f696_rdata));
  assign f696_clk = clk;
  assign f696_rst = rst;
  // Bindings to f696

  // f698
  logic [0:0] f698_wen;
  logic [31:0] f698_wdata;
  logic [0:0] f698_clk;
  logic [0:0] f698_rst;
  logic [31:0] f698_rdata;
  sr_buffer_32_1 f698(.wen(f698_wen), .wdata(f698_wdata), .clk(f698_clk), .rst(f698_rst), .rdata(f698_rdata));
  assign f698_clk = clk;
  assign f698_rst = rst;
  // Bindings to f698

  // f700
  logic [0:0] f700_wen;
  logic [31:0] f700_wdata;
  logic [0:0] f700_clk;
  logic [0:0] f700_rst;
  logic [31:0] f700_rdata;
  sr_buffer_32_1 f700(.wen(f700_wen), .wdata(f700_wdata), .clk(f700_clk), .rst(f700_rst), .rdata(f700_rdata));
  assign f700_clk = clk;
  assign f700_rst = rst;
  // Bindings to f700

  // f702
  logic [0:0] f702_wen;
  logic [31:0] f702_wdata;
  logic [0:0] f702_clk;
  logic [0:0] f702_rst;
  logic [31:0] f702_rdata;
  sr_buffer_32_1 f702(.wen(f702_wen), .wdata(f702_wdata), .clk(f702_clk), .rst(f702_rst), .rdata(f702_rdata));
  assign f702_clk = clk;
  assign f702_rst = rst;
  // Bindings to f702

  // f704
  logic [0:0] f704_wen;
  logic [31:0] f704_wdata;
  logic [0:0] f704_clk;
  logic [0:0] f704_rst;
  logic [31:0] f704_rdata;
  sr_buffer_32_1 f704(.wen(f704_wen), .wdata(f704_wdata), .clk(f704_clk), .rst(f704_rst), .rdata(f704_rdata));
  assign f704_clk = clk;
  assign f704_rst = rst;
  // Bindings to f704

  // f706
  logic [0:0] f706_wen;
  logic [31:0] f706_wdata;
  logic [0:0] f706_clk;
  logic [0:0] f706_rst;
  logic [31:0] f706_rdata;
  sr_buffer_32_1 f706(.wen(f706_wen), .wdata(f706_wdata), .clk(f706_clk), .rst(f706_rst), .rdata(f706_rdata));
  assign f706_clk = clk;
  assign f706_rst = rst;
  // Bindings to f706

  // f708
  logic [0:0] f708_wen;
  logic [31:0] f708_wdata;
  logic [0:0] f708_clk;
  logic [0:0] f708_rst;
  logic [31:0] f708_rdata;
  sr_buffer_32_1 f708(.wen(f708_wen), .wdata(f708_wdata), .clk(f708_clk), .rst(f708_rst), .rdata(f708_rdata));
  assign f708_clk = clk;
  assign f708_rst = rst;
  // Bindings to f708

  // f710
  logic [0:0] f710_wen;
  logic [31:0] f710_wdata;
  logic [0:0] f710_clk;
  logic [0:0] f710_rst;
  logic [31:0] f710_rdata;
  sr_buffer_32_1 f710(.wen(f710_wen), .wdata(f710_wdata), .clk(f710_clk), .rst(f710_rst), .rdata(f710_rdata));
  assign f710_clk = clk;
  assign f710_rst = rst;
  // Bindings to f710

  // f712
  logic [0:0] f712_wen;
  logic [31:0] f712_wdata;
  logic [0:0] f712_clk;
  logic [0:0] f712_rst;
  logic [31:0] f712_rdata;
  sr_buffer_32_1 f712(.wen(f712_wen), .wdata(f712_wdata), .clk(f712_clk), .rst(f712_rst), .rdata(f712_rdata));
  assign f712_clk = clk;
  assign f712_rst = rst;
  // Bindings to f712

  // f714
  logic [0:0] f714_wen;
  logic [31:0] f714_wdata;
  logic [0:0] f714_clk;
  logic [0:0] f714_rst;
  logic [31:0] f714_rdata;
  sr_buffer_32_1 f714(.wen(f714_wen), .wdata(f714_wdata), .clk(f714_clk), .rst(f714_rst), .rdata(f714_rdata));
  assign f714_clk = clk;
  assign f714_rst = rst;
  // Bindings to f714

  // f716
  logic [0:0] f716_wen;
  logic [31:0] f716_wdata;
  logic [0:0] f716_clk;
  logic [0:0] f716_rst;
  logic [31:0] f716_rdata;
  sr_buffer_32_1 f716(.wen(f716_wen), .wdata(f716_wdata), .clk(f716_clk), .rst(f716_rst), .rdata(f716_rdata));
  assign f716_clk = clk;
  assign f716_rst = rst;
  // Bindings to f716

  // f718
  logic [0:0] f718_wen;
  logic [31:0] f718_wdata;
  logic [0:0] f718_clk;
  logic [0:0] f718_rst;
  logic [31:0] f718_rdata;
  sr_buffer_32_1 f718(.wen(f718_wen), .wdata(f718_wdata), .clk(f718_clk), .rst(f718_rst), .rdata(f718_rdata));
  assign f718_clk = clk;
  assign f718_rst = rst;
  // Bindings to f718

  // f720
  logic [0:0] f720_wen;
  logic [31:0] f720_wdata;
  logic [0:0] f720_clk;
  logic [0:0] f720_rst;
  logic [31:0] f720_rdata;
  sr_buffer_32_1 f720(.wen(f720_wen), .wdata(f720_wdata), .clk(f720_clk), .rst(f720_rst), .rdata(f720_rdata));
  assign f720_clk = clk;
  assign f720_rst = rst;
  // Bindings to f720

  // f722
  logic [0:0] f722_wen;
  logic [31:0] f722_wdata;
  logic [0:0] f722_clk;
  logic [0:0] f722_rst;
  logic [31:0] f722_rdata;
  sr_buffer_32_1 f722(.wen(f722_wen), .wdata(f722_wdata), .clk(f722_clk), .rst(f722_rst), .rdata(f722_rdata));
  assign f722_clk = clk;
  assign f722_rst = rst;
  // Bindings to f722

  // f724
  logic [0:0] f724_wen;
  logic [31:0] f724_wdata;
  logic [0:0] f724_clk;
  logic [0:0] f724_rst;
  logic [31:0] f724_rdata;
  sr_buffer_32_1 f724(.wen(f724_wen), .wdata(f724_wdata), .clk(f724_clk), .rst(f724_rst), .rdata(f724_rdata));
  assign f724_clk = clk;
  assign f724_rst = rst;
  // Bindings to f724

  // f726
  logic [0:0] f726_wen;
  logic [31:0] f726_wdata;
  logic [0:0] f726_clk;
  logic [0:0] f726_rst;
  logic [31:0] f726_rdata;
  sr_buffer_32_1 f726(.wen(f726_wen), .wdata(f726_wdata), .clk(f726_clk), .rst(f726_rst), .rdata(f726_rdata));
  assign f726_clk = clk;
  assign f726_rst = rst;
  // Bindings to f726

  // f728
  logic [0:0] f728_wen;
  logic [31:0] f728_wdata;
  logic [0:0] f728_clk;
  logic [0:0] f728_rst;
  logic [31:0] f728_rdata;
  sr_buffer_32_1 f728(.wen(f728_wen), .wdata(f728_wdata), .clk(f728_clk), .rst(f728_rst), .rdata(f728_rdata));
  assign f728_clk = clk;
  assign f728_rst = rst;
  // Bindings to f728

  // f730
  logic [0:0] f730_wen;
  logic [31:0] f730_wdata;
  logic [0:0] f730_clk;
  logic [0:0] f730_rst;
  logic [31:0] f730_rdata;
  sr_buffer_32_1 f730(.wen(f730_wen), .wdata(f730_wdata), .clk(f730_clk), .rst(f730_rst), .rdata(f730_rdata));
  assign f730_clk = clk;
  assign f730_rst = rst;
  // Bindings to f730

  // f732
  logic [0:0] f732_wen;
  logic [31:0] f732_wdata;
  logic [0:0] f732_clk;
  logic [0:0] f732_rst;
  logic [31:0] f732_rdata;
  sr_buffer_32_1 f732(.wen(f732_wen), .wdata(f732_wdata), .clk(f732_clk), .rst(f732_rst), .rdata(f732_rdata));
  assign f732_clk = clk;
  assign f732_rst = rst;
  // Bindings to f732

  // f734
  logic [0:0] f734_wen;
  logic [31:0] f734_wdata;
  logic [0:0] f734_clk;
  logic [0:0] f734_rst;
  logic [31:0] f734_rdata;
  sr_buffer_32_1 f734(.wen(f734_wen), .wdata(f734_wdata), .clk(f734_clk), .rst(f734_rst), .rdata(f734_rdata));
  assign f734_clk = clk;
  assign f734_rst = rst;
  // Bindings to f734

  // f736
  logic [0:0] f736_wen;
  logic [31:0] f736_wdata;
  logic [0:0] f736_clk;
  logic [0:0] f736_rst;
  logic [31:0] f736_rdata;
  sr_buffer_32_1 f736(.wen(f736_wen), .wdata(f736_wdata), .clk(f736_clk), .rst(f736_rst), .rdata(f736_rdata));
  assign f736_clk = clk;
  assign f736_rst = rst;
  // Bindings to f736

  // f738
  logic [0:0] f738_wen;
  logic [31:0] f738_wdata;
  logic [0:0] f738_clk;
  logic [0:0] f738_rst;
  logic [31:0] f738_rdata;
  sr_buffer_32_1 f738(.wen(f738_wen), .wdata(f738_wdata), .clk(f738_clk), .rst(f738_rst), .rdata(f738_rdata));
  assign f738_clk = clk;
  assign f738_rst = rst;
  // Bindings to f738

  // f740
  logic [0:0] f740_wen;
  logic [31:0] f740_wdata;
  logic [0:0] f740_clk;
  logic [0:0] f740_rst;
  logic [31:0] f740_rdata;
  sr_buffer_32_1 f740(.wen(f740_wen), .wdata(f740_wdata), .clk(f740_clk), .rst(f740_rst), .rdata(f740_rdata));
  assign f740_clk = clk;
  assign f740_rst = rst;
  // Bindings to f740

  // f742
  logic [0:0] f742_wen;
  logic [31:0] f742_wdata;
  logic [0:0] f742_clk;
  logic [0:0] f742_rst;
  logic [31:0] f742_rdata;
  sr_buffer_32_1 f742(.wen(f742_wen), .wdata(f742_wdata), .clk(f742_clk), .rst(f742_rst), .rdata(f742_rdata));
  assign f742_clk = clk;
  assign f742_rst = rst;
  // Bindings to f742

  // f744
  logic [0:0] f744_wen;
  logic [31:0] f744_wdata;
  logic [0:0] f744_clk;
  logic [0:0] f744_rst;
  logic [31:0] f744_rdata;
  sr_buffer_32_1 f744(.wen(f744_wen), .wdata(f744_wdata), .clk(f744_clk), .rst(f744_rst), .rdata(f744_rdata));
  assign f744_clk = clk;
  assign f744_rst = rst;
  // Bindings to f744

  // f746
  logic [0:0] f746_wen;
  logic [31:0] f746_wdata;
  logic [0:0] f746_clk;
  logic [0:0] f746_rst;
  logic [31:0] f746_rdata;
  sr_buffer_32_1 f746(.wen(f746_wen), .wdata(f746_wdata), .clk(f746_clk), .rst(f746_rst), .rdata(f746_rdata));
  assign f746_clk = clk;
  assign f746_rst = rst;
  // Bindings to f746

  // f748
  logic [0:0] f748_wen;
  logic [31:0] f748_wdata;
  logic [0:0] f748_clk;
  logic [0:0] f748_rst;
  logic [31:0] f748_rdata;
  sr_buffer_32_1 f748(.wen(f748_wen), .wdata(f748_wdata), .clk(f748_clk), .rst(f748_rst), .rdata(f748_rdata));
  assign f748_clk = clk;
  assign f748_rst = rst;
  // Bindings to f748

  // f750
  logic [0:0] f750_wen;
  logic [31:0] f750_wdata;
  logic [0:0] f750_clk;
  logic [0:0] f750_rst;
  logic [31:0] f750_rdata;
  sr_buffer_32_1 f750(.wen(f750_wen), .wdata(f750_wdata), .clk(f750_clk), .rst(f750_rst), .rdata(f750_rdata));
  assign f750_clk = clk;
  assign f750_rst = rst;
  // Bindings to f750

  // f752
  logic [0:0] f752_wen;
  logic [31:0] f752_wdata;
  logic [0:0] f752_clk;
  logic [0:0] f752_rst;
  logic [31:0] f752_rdata;
  sr_buffer_32_1 f752(.wen(f752_wen), .wdata(f752_wdata), .clk(f752_clk), .rst(f752_rst), .rdata(f752_rdata));
  assign f752_clk = clk;
  assign f752_rst = rst;
  // Bindings to f752

  // f754
  logic [0:0] f754_wen;
  logic [31:0] f754_wdata;
  logic [0:0] f754_clk;
  logic [0:0] f754_rst;
  logic [31:0] f754_rdata;
  sr_buffer_32_1 f754(.wen(f754_wen), .wdata(f754_wdata), .clk(f754_clk), .rst(f754_rst), .rdata(f754_rdata));
  assign f754_clk = clk;
  assign f754_rst = rst;
  // Bindings to f754

  // f756
  logic [0:0] f756_wen;
  logic [31:0] f756_wdata;
  logic [0:0] f756_clk;
  logic [0:0] f756_rst;
  logic [31:0] f756_rdata;
  sr_buffer_32_1 f756(.wen(f756_wen), .wdata(f756_wdata), .clk(f756_clk), .rst(f756_rst), .rdata(f756_rdata));
  assign f756_clk = clk;
  assign f756_rst = rst;
  // Bindings to f756

  // f758
  logic [0:0] f758_wen;
  logic [31:0] f758_wdata;
  logic [0:0] f758_clk;
  logic [0:0] f758_rst;
  logic [31:0] f758_rdata;
  sr_buffer_32_1 f758(.wen(f758_wen), .wdata(f758_wdata), .clk(f758_clk), .rst(f758_rst), .rdata(f758_rdata));
  assign f758_clk = clk;
  assign f758_rst = rst;
  // Bindings to f758

  // f760
  logic [0:0] f760_wen;
  logic [31:0] f760_wdata;
  logic [0:0] f760_clk;
  logic [0:0] f760_rst;
  logic [31:0] f760_rdata;
  sr_buffer_32_1 f760(.wen(f760_wen), .wdata(f760_wdata), .clk(f760_clk), .rst(f760_rst), .rdata(f760_rdata));
  assign f760_clk = clk;
  assign f760_rst = rst;
  // Bindings to f760

  // f762
  logic [0:0] f762_wen;
  logic [31:0] f762_wdata;
  logic [0:0] f762_clk;
  logic [0:0] f762_rst;
  logic [31:0] f762_rdata;
  sr_buffer_32_1 f762(.wen(f762_wen), .wdata(f762_wdata), .clk(f762_clk), .rst(f762_rst), .rdata(f762_rdata));
  assign f762_clk = clk;
  assign f762_rst = rst;
  // Bindings to f762

  // f764
  logic [0:0] f764_wen;
  logic [31:0] f764_wdata;
  logic [0:0] f764_clk;
  logic [0:0] f764_rst;
  logic [31:0] f764_rdata;
  sr_buffer_32_1 f764(.wen(f764_wen), .wdata(f764_wdata), .clk(f764_clk), .rst(f764_rst), .rdata(f764_rdata));
  assign f764_clk = clk;
  assign f764_rst = rst;
  // Bindings to f764

  // f766
  logic [0:0] f766_wen;
  logic [31:0] f766_wdata;
  logic [0:0] f766_clk;
  logic [0:0] f766_rst;
  logic [31:0] f766_rdata;
  sr_buffer_32_1 f766(.wen(f766_wen), .wdata(f766_wdata), .clk(f766_clk), .rst(f766_rst), .rdata(f766_rdata));
  assign f766_clk = clk;
  assign f766_rst = rst;
  // Bindings to f766

  // f768
  logic [0:0] f768_wen;
  logic [31:0] f768_wdata;
  logic [0:0] f768_clk;
  logic [0:0] f768_rst;
  logic [31:0] f768_rdata;
  sr_buffer_32_1 f768(.wen(f768_wen), .wdata(f768_wdata), .clk(f768_clk), .rst(f768_rst), .rdata(f768_rdata));
  assign f768_clk = clk;
  assign f768_rst = rst;
  // Bindings to f768

  // f770
  logic [0:0] f770_wen;
  logic [31:0] f770_wdata;
  logic [0:0] f770_clk;
  logic [0:0] f770_rst;
  logic [31:0] f770_rdata;
  sr_buffer_32_1 f770(.wen(f770_wen), .wdata(f770_wdata), .clk(f770_clk), .rst(f770_rst), .rdata(f770_rdata));
  assign f770_clk = clk;
  assign f770_rst = rst;
  // Bindings to f770

  // f772
  logic [0:0] f772_wen;
  logic [31:0] f772_wdata;
  logic [0:0] f772_clk;
  logic [0:0] f772_rst;
  logic [31:0] f772_rdata;
  sr_buffer_32_1 f772(.wen(f772_wen), .wdata(f772_wdata), .clk(f772_clk), .rst(f772_rst), .rdata(f772_rdata));
  assign f772_clk = clk;
  assign f772_rst = rst;
  // Bindings to f772

  // f774
  logic [0:0] f774_wen;
  logic [31:0] f774_wdata;
  logic [0:0] f774_clk;
  logic [0:0] f774_rst;
  logic [31:0] f774_rdata;
  sr_buffer_32_1 f774(.wen(f774_wen), .wdata(f774_wdata), .clk(f774_clk), .rst(f774_rst), .rdata(f774_rdata));
  assign f774_clk = clk;
  assign f774_rst = rst;
  // Bindings to f774

  // f776
  logic [0:0] f776_wen;
  logic [31:0] f776_wdata;
  logic [0:0] f776_clk;
  logic [0:0] f776_rst;
  logic [31:0] f776_rdata;
  sr_buffer_32_1 f776(.wen(f776_wen), .wdata(f776_wdata), .clk(f776_clk), .rst(f776_rst), .rdata(f776_rdata));
  assign f776_clk = clk;
  assign f776_rst = rst;
  // Bindings to f776

  // f778
  logic [0:0] f778_wen;
  logic [31:0] f778_wdata;
  logic [0:0] f778_clk;
  logic [0:0] f778_rst;
  logic [31:0] f778_rdata;
  sr_buffer_32_1 f778(.wen(f778_wen), .wdata(f778_wdata), .clk(f778_clk), .rst(f778_rst), .rdata(f778_rdata));
  assign f778_clk = clk;
  assign f778_rst = rst;
  // Bindings to f778

  // f780
  logic [0:0] f780_wen;
  logic [31:0] f780_wdata;
  logic [0:0] f780_clk;
  logic [0:0] f780_rst;
  logic [31:0] f780_rdata;
  sr_buffer_32_1 f780(.wen(f780_wen), .wdata(f780_wdata), .clk(f780_clk), .rst(f780_rst), .rdata(f780_rdata));
  assign f780_clk = clk;
  assign f780_rst = rst;
  // Bindings to f780

  // f782
  logic [0:0] f782_wen;
  logic [31:0] f782_wdata;
  logic [0:0] f782_clk;
  logic [0:0] f782_rst;
  logic [31:0] f782_rdata;
  sr_buffer_32_1 f782(.wen(f782_wen), .wdata(f782_wdata), .clk(f782_clk), .rst(f782_rst), .rdata(f782_rdata));
  assign f782_clk = clk;
  assign f782_rst = rst;
  // Bindings to f782

  // f784
  logic [0:0] f784_wen;
  logic [31:0] f784_wdata;
  logic [0:0] f784_clk;
  logic [0:0] f784_rst;
  logic [31:0] f784_rdata;
  sr_buffer_32_1 f784(.wen(f784_wen), .wdata(f784_wdata), .clk(f784_clk), .rst(f784_rst), .rdata(f784_rdata));
  assign f784_clk = clk;
  assign f784_rst = rst;
  // Bindings to f784

  // f786
  logic [0:0] f786_wen;
  logic [31:0] f786_wdata;
  logic [0:0] f786_clk;
  logic [0:0] f786_rst;
  logic [31:0] f786_rdata;
  sr_buffer_32_1 f786(.wen(f786_wen), .wdata(f786_wdata), .clk(f786_clk), .rst(f786_rst), .rdata(f786_rdata));
  assign f786_clk = clk;
  assign f786_rst = rst;
  // Bindings to f786

  // f788
  logic [0:0] f788_wen;
  logic [31:0] f788_wdata;
  logic [0:0] f788_clk;
  logic [0:0] f788_rst;
  logic [31:0] f788_rdata;
  sr_buffer_32_1 f788(.wen(f788_wen), .wdata(f788_wdata), .clk(f788_clk), .rst(f788_rst), .rdata(f788_rdata));
  assign f788_clk = clk;
  assign f788_rst = rst;
  // Bindings to f788

  // f790
  logic [0:0] f790_wen;
  logic [31:0] f790_wdata;
  logic [0:0] f790_clk;
  logic [0:0] f790_rst;
  logic [31:0] f790_rdata;
  sr_buffer_32_1 f790(.wen(f790_wen), .wdata(f790_wdata), .clk(f790_clk), .rst(f790_rst), .rdata(f790_rdata));
  assign f790_clk = clk;
  assign f790_rst = rst;
  // Bindings to f790

  // f792
  logic [0:0] f792_wen;
  logic [31:0] f792_wdata;
  logic [0:0] f792_clk;
  logic [0:0] f792_rst;
  logic [31:0] f792_rdata;
  sr_buffer_32_1 f792(.wen(f792_wen), .wdata(f792_wdata), .clk(f792_clk), .rst(f792_rst), .rdata(f792_rdata));
  assign f792_clk = clk;
  assign f792_rst = rst;
  // Bindings to f792

  // f794
  logic [0:0] f794_wen;
  logic [31:0] f794_wdata;
  logic [0:0] f794_clk;
  logic [0:0] f794_rst;
  logic [31:0] f794_rdata;
  sr_buffer_32_1 f794(.wen(f794_wen), .wdata(f794_wdata), .clk(f794_clk), .rst(f794_rst), .rdata(f794_rdata));
  assign f794_clk = clk;
  assign f794_rst = rst;
  // Bindings to f794

  // f796
  logic [0:0] f796_wen;
  logic [31:0] f796_wdata;
  logic [0:0] f796_clk;
  logic [0:0] f796_rst;
  logic [31:0] f796_rdata;
  sr_buffer_32_1 f796(.wen(f796_wen), .wdata(f796_wdata), .clk(f796_clk), .rst(f796_rst), .rdata(f796_rdata));
  assign f796_clk = clk;
  assign f796_rst = rst;
  // Bindings to f796

  // f798
  logic [0:0] f798_wen;
  logic [31:0] f798_wdata;
  logic [0:0] f798_clk;
  logic [0:0] f798_rst;
  logic [31:0] f798_rdata;
  sr_buffer_32_1 f798(.wen(f798_wen), .wdata(f798_wdata), .clk(f798_clk), .rst(f798_rst), .rdata(f798_rdata));
  assign f798_clk = clk;
  assign f798_rst = rst;
  // Bindings to f798

  // f800
  logic [0:0] f800_wen;
  logic [31:0] f800_wdata;
  logic [0:0] f800_clk;
  logic [0:0] f800_rst;
  logic [31:0] f800_rdata;
  sr_buffer_32_1 f800(.wen(f800_wen), .wdata(f800_wdata), .clk(f800_clk), .rst(f800_rst), .rdata(f800_rdata));
  assign f800_clk = clk;
  assign f800_rst = rst;
  // Bindings to f800

  // f802
  logic [0:0] f802_wen;
  logic [31:0] f802_wdata;
  logic [0:0] f802_clk;
  logic [0:0] f802_rst;
  logic [31:0] f802_rdata;
  sr_buffer_32_1 f802(.wen(f802_wen), .wdata(f802_wdata), .clk(f802_clk), .rst(f802_rst), .rdata(f802_rdata));
  assign f802_clk = clk;
  assign f802_rst = rst;
  // Bindings to f802

  // f804
  logic [0:0] f804_wen;
  logic [31:0] f804_wdata;
  logic [0:0] f804_clk;
  logic [0:0] f804_rst;
  logic [31:0] f804_rdata;
  sr_buffer_32_1 f804(.wen(f804_wen), .wdata(f804_wdata), .clk(f804_clk), .rst(f804_rst), .rdata(f804_rdata));
  assign f804_clk = clk;
  assign f804_rst = rst;
  // Bindings to f804

  // f806
  logic [0:0] f806_wen;
  logic [31:0] f806_wdata;
  logic [0:0] f806_clk;
  logic [0:0] f806_rst;
  logic [31:0] f806_rdata;
  sr_buffer_32_1 f806(.wen(f806_wen), .wdata(f806_wdata), .clk(f806_clk), .rst(f806_rst), .rdata(f806_rdata));
  assign f806_clk = clk;
  assign f806_rst = rst;
  // Bindings to f806

  // f808
  logic [0:0] f808_wen;
  logic [31:0] f808_wdata;
  logic [0:0] f808_clk;
  logic [0:0] f808_rst;
  logic [31:0] f808_rdata;
  sr_buffer_32_1 f808(.wen(f808_wen), .wdata(f808_wdata), .clk(f808_clk), .rst(f808_rst), .rdata(f808_rdata));
  assign f808_clk = clk;
  assign f808_rst = rst;
  // Bindings to f808

  // f810
  logic [0:0] f810_wen;
  logic [31:0] f810_wdata;
  logic [0:0] f810_clk;
  logic [0:0] f810_rst;
  logic [31:0] f810_rdata;
  sr_buffer_32_1 f810(.wen(f810_wen), .wdata(f810_wdata), .clk(f810_clk), .rst(f810_rst), .rdata(f810_rdata));
  assign f810_clk = clk;
  assign f810_rst = rst;
  // Bindings to f810

  // f812
  logic [0:0] f812_wen;
  logic [31:0] f812_wdata;
  logic [0:0] f812_clk;
  logic [0:0] f812_rst;
  logic [31:0] f812_rdata;
  sr_buffer_32_1 f812(.wen(f812_wen), .wdata(f812_wdata), .clk(f812_clk), .rst(f812_rst), .rdata(f812_rdata));
  assign f812_clk = clk;
  assign f812_rst = rst;
  // Bindings to f812

  // f814
  logic [0:0] f814_wen;
  logic [31:0] f814_wdata;
  logic [0:0] f814_clk;
  logic [0:0] f814_rst;
  logic [31:0] f814_rdata;
  sr_buffer_32_1 f814(.wen(f814_wen), .wdata(f814_wdata), .clk(f814_clk), .rst(f814_rst), .rdata(f814_rdata));
  assign f814_clk = clk;
  assign f814_rst = rst;
  // Bindings to f814

  // f816
  logic [0:0] f816_wen;
  logic [31:0] f816_wdata;
  logic [0:0] f816_clk;
  logic [0:0] f816_rst;
  logic [31:0] f816_rdata;
  sr_buffer_32_1 f816(.wen(f816_wen), .wdata(f816_wdata), .clk(f816_clk), .rst(f816_rst), .rdata(f816_rdata));
  assign f816_clk = clk;
  assign f816_rst = rst;
  // Bindings to f816

  // f818
  logic [0:0] f818_wen;
  logic [31:0] f818_wdata;
  logic [0:0] f818_clk;
  logic [0:0] f818_rst;
  logic [31:0] f818_rdata;
  sr_buffer_32_1 f818(.wen(f818_wen), .wdata(f818_wdata), .clk(f818_clk), .rst(f818_rst), .rdata(f818_rdata));
  assign f818_clk = clk;
  assign f818_rst = rst;
  // Bindings to f818

  // f820
  logic [0:0] f820_wen;
  logic [31:0] f820_wdata;
  logic [0:0] f820_clk;
  logic [0:0] f820_rst;
  logic [31:0] f820_rdata;
  sr_buffer_32_1 f820(.wen(f820_wen), .wdata(f820_wdata), .clk(f820_clk), .rst(f820_rst), .rdata(f820_rdata));
  assign f820_clk = clk;
  assign f820_rst = rst;
  // Bindings to f820

  // f822
  logic [0:0] f822_wen;
  logic [31:0] f822_wdata;
  logic [0:0] f822_clk;
  logic [0:0] f822_rst;
  logic [31:0] f822_rdata;
  sr_buffer_32_1 f822(.wen(f822_wen), .wdata(f822_wdata), .clk(f822_clk), .rst(f822_rst), .rdata(f822_rdata));
  assign f822_clk = clk;
  assign f822_rst = rst;
  // Bindings to f822

  // f824
  logic [0:0] f824_wen;
  logic [31:0] f824_wdata;
  logic [0:0] f824_clk;
  logic [0:0] f824_rst;
  logic [31:0] f824_rdata;
  sr_buffer_32_1 f824(.wen(f824_wen), .wdata(f824_wdata), .clk(f824_clk), .rst(f824_rst), .rdata(f824_rdata));
  assign f824_clk = clk;
  assign f824_rst = rst;
  // Bindings to f824

  // f826
  logic [0:0] f826_wen;
  logic [31:0] f826_wdata;
  logic [0:0] f826_clk;
  logic [0:0] f826_rst;
  logic [31:0] f826_rdata;
  sr_buffer_32_1 f826(.wen(f826_wen), .wdata(f826_wdata), .clk(f826_clk), .rst(f826_rst), .rdata(f826_rdata));
  assign f826_clk = clk;
  assign f826_rst = rst;
  // Bindings to f826

  // f828
  logic [0:0] f828_wen;
  logic [31:0] f828_wdata;
  logic [0:0] f828_clk;
  logic [0:0] f828_rst;
  logic [31:0] f828_rdata;
  sr_buffer_32_1 f828(.wen(f828_wen), .wdata(f828_wdata), .clk(f828_clk), .rst(f828_rst), .rdata(f828_rdata));
  assign f828_clk = clk;
  assign f828_rst = rst;
  // Bindings to f828

  // f830
  logic [0:0] f830_wen;
  logic [31:0] f830_wdata;
  logic [0:0] f830_clk;
  logic [0:0] f830_rst;
  logic [31:0] f830_rdata;
  sr_buffer_32_1 f830(.wen(f830_wen), .wdata(f830_wdata), .clk(f830_clk), .rst(f830_rst), .rdata(f830_rdata));
  assign f830_clk = clk;
  assign f830_rst = rst;
  // Bindings to f830

  // f832
  logic [0:0] f832_wen;
  logic [31:0] f832_wdata;
  logic [0:0] f832_clk;
  logic [0:0] f832_rst;
  logic [31:0] f832_rdata;
  sr_buffer_32_1 f832(.wen(f832_wen), .wdata(f832_wdata), .clk(f832_clk), .rst(f832_rst), .rdata(f832_rdata));
  assign f832_clk = clk;
  assign f832_rst = rst;
  // Bindings to f832

  // f834
  logic [0:0] f834_wen;
  logic [31:0] f834_wdata;
  logic [0:0] f834_clk;
  logic [0:0] f834_rst;
  logic [31:0] f834_rdata;
  sr_buffer_32_1 f834(.wen(f834_wen), .wdata(f834_wdata), .clk(f834_clk), .rst(f834_rst), .rdata(f834_rdata));
  assign f834_clk = clk;
  assign f834_rst = rst;
  // Bindings to f834

  // f836
  logic [0:0] f836_wen;
  logic [31:0] f836_wdata;
  logic [0:0] f836_clk;
  logic [0:0] f836_rst;
  logic [31:0] f836_rdata;
  sr_buffer_32_1 f836(.wen(f836_wen), .wdata(f836_wdata), .clk(f836_clk), .rst(f836_rst), .rdata(f836_rdata));
  assign f836_clk = clk;
  assign f836_rst = rst;
  // Bindings to f836

  // f838
  logic [0:0] f838_wen;
  logic [31:0] f838_wdata;
  logic [0:0] f838_clk;
  logic [0:0] f838_rst;
  logic [31:0] f838_rdata;
  sr_buffer_32_1 f838(.wen(f838_wen), .wdata(f838_wdata), .clk(f838_clk), .rst(f838_rst), .rdata(f838_rdata));
  assign f838_clk = clk;
  assign f838_rst = rst;
  // Bindings to f838

  // f840
  logic [0:0] f840_wen;
  logic [31:0] f840_wdata;
  logic [0:0] f840_clk;
  logic [0:0] f840_rst;
  logic [31:0] f840_rdata;
  sr_buffer_32_1 f840(.wen(f840_wen), .wdata(f840_wdata), .clk(f840_clk), .rst(f840_rst), .rdata(f840_rdata));
  assign f840_clk = clk;
  assign f840_rst = rst;
  // Bindings to f840

  // f842
  logic [0:0] f842_wen;
  logic [31:0] f842_wdata;
  logic [0:0] f842_clk;
  logic [0:0] f842_rst;
  logic [31:0] f842_rdata;
  sr_buffer_32_1 f842(.wen(f842_wen), .wdata(f842_wdata), .clk(f842_clk), .rst(f842_rst), .rdata(f842_rdata));
  assign f842_clk = clk;
  assign f842_rst = rst;
  // Bindings to f842

  // f844
  logic [0:0] f844_wen;
  logic [31:0] f844_wdata;
  logic [0:0] f844_clk;
  logic [0:0] f844_rst;
  logic [31:0] f844_rdata;
  sr_buffer_32_1 f844(.wen(f844_wen), .wdata(f844_wdata), .clk(f844_clk), .rst(f844_rst), .rdata(f844_rdata));
  assign f844_clk = clk;
  assign f844_rst = rst;
  // Bindings to f844

  // f846
  logic [0:0] f846_wen;
  logic [31:0] f846_wdata;
  logic [0:0] f846_clk;
  logic [0:0] f846_rst;
  logic [31:0] f846_rdata;
  sr_buffer_32_1 f846(.wen(f846_wen), .wdata(f846_wdata), .clk(f846_clk), .rst(f846_rst), .rdata(f846_rdata));
  assign f846_clk = clk;
  assign f846_rst = rst;
  // Bindings to f846

  // f848
  logic [0:0] f848_wen;
  logic [31:0] f848_wdata;
  logic [0:0] f848_clk;
  logic [0:0] f848_rst;
  logic [31:0] f848_rdata;
  sr_buffer_32_1 f848(.wen(f848_wen), .wdata(f848_wdata), .clk(f848_clk), .rst(f848_rst), .rdata(f848_rdata));
  assign f848_clk = clk;
  assign f848_rst = rst;
  // Bindings to f848

  // f850
  logic [0:0] f850_wen;
  logic [31:0] f850_wdata;
  logic [0:0] f850_clk;
  logic [0:0] f850_rst;
  logic [31:0] f850_rdata;
  sr_buffer_32_1 f850(.wen(f850_wen), .wdata(f850_wdata), .clk(f850_clk), .rst(f850_rst), .rdata(f850_rdata));
  assign f850_clk = clk;
  assign f850_rst = rst;
  // Bindings to f850

  // f852
  logic [0:0] f852_wen;
  logic [31:0] f852_wdata;
  logic [0:0] f852_clk;
  logic [0:0] f852_rst;
  logic [31:0] f852_rdata;
  sr_buffer_32_1 f852(.wen(f852_wen), .wdata(f852_wdata), .clk(f852_clk), .rst(f852_rst), .rdata(f852_rdata));
  assign f852_clk = clk;
  assign f852_rst = rst;
  // Bindings to f852

  // f854
  logic [0:0] f854_wen;
  logic [31:0] f854_wdata;
  logic [0:0] f854_clk;
  logic [0:0] f854_rst;
  logic [31:0] f854_rdata;
  sr_buffer_32_1 f854(.wen(f854_wen), .wdata(f854_wdata), .clk(f854_clk), .rst(f854_rst), .rdata(f854_rdata));
  assign f854_clk = clk;
  assign f854_rst = rst;
  // Bindings to f854

  // f856
  logic [0:0] f856_wen;
  logic [31:0] f856_wdata;
  logic [0:0] f856_clk;
  logic [0:0] f856_rst;
  logic [31:0] f856_rdata;
  sr_buffer_32_1 f856(.wen(f856_wen), .wdata(f856_wdata), .clk(f856_clk), .rst(f856_rst), .rdata(f856_rdata));
  assign f856_clk = clk;
  assign f856_rst = rst;
  // Bindings to f856

  // f858
  logic [0:0] f858_wen;
  logic [31:0] f858_wdata;
  logic [0:0] f858_clk;
  logic [0:0] f858_rst;
  logic [31:0] f858_rdata;
  sr_buffer_32_1 f858(.wen(f858_wen), .wdata(f858_wdata), .clk(f858_clk), .rst(f858_rst), .rdata(f858_rdata));
  assign f858_clk = clk;
  assign f858_rst = rst;
  // Bindings to f858

  // f860
  logic [0:0] f860_wen;
  logic [31:0] f860_wdata;
  logic [0:0] f860_clk;
  logic [0:0] f860_rst;
  logic [31:0] f860_rdata;
  sr_buffer_32_1 f860(.wen(f860_wen), .wdata(f860_wdata), .clk(f860_clk), .rst(f860_rst), .rdata(f860_rdata));
  assign f860_clk = clk;
  assign f860_rst = rst;
  // Bindings to f860

  // f862
  logic [0:0] f862_wen;
  logic [31:0] f862_wdata;
  logic [0:0] f862_clk;
  logic [0:0] f862_rst;
  logic [31:0] f862_rdata;
  sr_buffer_32_1 f862(.wen(f862_wen), .wdata(f862_wdata), .clk(f862_clk), .rst(f862_rst), .rdata(f862_rdata));
  assign f862_clk = clk;
  assign f862_rst = rst;
  // Bindings to f862

  // f864
  logic [0:0] f864_wen;
  logic [31:0] f864_wdata;
  logic [0:0] f864_clk;
  logic [0:0] f864_rst;
  logic [31:0] f864_rdata;
  sr_buffer_32_1 f864(.wen(f864_wen), .wdata(f864_wdata), .clk(f864_clk), .rst(f864_rst), .rdata(f864_rdata));
  assign f864_clk = clk;
  assign f864_rst = rst;
  // Bindings to f864

  // f866
  logic [0:0] f866_wen;
  logic [31:0] f866_wdata;
  logic [0:0] f866_clk;
  logic [0:0] f866_rst;
  logic [31:0] f866_rdata;
  sr_buffer_32_1 f866(.wen(f866_wen), .wdata(f866_wdata), .clk(f866_clk), .rst(f866_rst), .rdata(f866_rdata));
  assign f866_clk = clk;
  assign f866_rst = rst;
  // Bindings to f866

  // f868
  logic [0:0] f868_wen;
  logic [31:0] f868_wdata;
  logic [0:0] f868_clk;
  logic [0:0] f868_rst;
  logic [31:0] f868_rdata;
  sr_buffer_32_1 f868(.wen(f868_wen), .wdata(f868_wdata), .clk(f868_clk), .rst(f868_rst), .rdata(f868_rdata));
  assign f868_clk = clk;
  assign f868_rst = rst;
  // Bindings to f868

  // f870
  logic [0:0] f870_wen;
  logic [31:0] f870_wdata;
  logic [0:0] f870_clk;
  logic [0:0] f870_rst;
  logic [31:0] f870_rdata;
  sr_buffer_32_1 f870(.wen(f870_wen), .wdata(f870_wdata), .clk(f870_clk), .rst(f870_rst), .rdata(f870_rdata));
  assign f870_clk = clk;
  assign f870_rst = rst;
  // Bindings to f870

  // f872
  logic [0:0] f872_wen;
  logic [31:0] f872_wdata;
  logic [0:0] f872_clk;
  logic [0:0] f872_rst;
  logic [31:0] f872_rdata;
  sr_buffer_32_1 f872(.wen(f872_wen), .wdata(f872_wdata), .clk(f872_clk), .rst(f872_rst), .rdata(f872_rdata));
  assign f872_clk = clk;
  assign f872_rst = rst;
  // Bindings to f872

  // f874
  logic [0:0] f874_wen;
  logic [31:0] f874_wdata;
  logic [0:0] f874_clk;
  logic [0:0] f874_rst;
  logic [31:0] f874_rdata;
  sr_buffer_32_1 f874(.wen(f874_wen), .wdata(f874_wdata), .clk(f874_clk), .rst(f874_rst), .rdata(f874_rdata));
  assign f874_clk = clk;
  assign f874_rst = rst;
  // Bindings to f874

  // f876
  logic [0:0] f876_wen;
  logic [31:0] f876_wdata;
  logic [0:0] f876_clk;
  logic [0:0] f876_rst;
  logic [31:0] f876_rdata;
  sr_buffer_32_1 f876(.wen(f876_wen), .wdata(f876_wdata), .clk(f876_clk), .rst(f876_rst), .rdata(f876_rdata));
  assign f876_clk = clk;
  assign f876_rst = rst;
  // Bindings to f876

  // f878
  logic [0:0] f878_wen;
  logic [31:0] f878_wdata;
  logic [0:0] f878_clk;
  logic [0:0] f878_rst;
  logic [31:0] f878_rdata;
  sr_buffer_32_1 f878(.wen(f878_wen), .wdata(f878_wdata), .clk(f878_clk), .rst(f878_rst), .rdata(f878_rdata));
  assign f878_clk = clk;
  assign f878_rst = rst;
  // Bindings to f878

  // f880
  logic [0:0] f880_wen;
  logic [31:0] f880_wdata;
  logic [0:0] f880_clk;
  logic [0:0] f880_rst;
  logic [31:0] f880_rdata;
  sr_buffer_32_1 f880(.wen(f880_wen), .wdata(f880_wdata), .clk(f880_clk), .rst(f880_rst), .rdata(f880_rdata));
  assign f880_clk = clk;
  assign f880_rst = rst;
  // Bindings to f880

  // f882
  logic [0:0] f882_wen;
  logic [31:0] f882_wdata;
  logic [0:0] f882_clk;
  logic [0:0] f882_rst;
  logic [31:0] f882_rdata;
  sr_buffer_32_1 f882(.wen(f882_wen), .wdata(f882_wdata), .clk(f882_clk), .rst(f882_rst), .rdata(f882_rdata));
  assign f882_clk = clk;
  assign f882_rst = rst;
  // Bindings to f882

  // f884
  logic [0:0] f884_wen;
  logic [31:0] f884_wdata;
  logic [0:0] f884_clk;
  logic [0:0] f884_rst;
  logic [31:0] f884_rdata;
  sr_buffer_32_1 f884(.wen(f884_wen), .wdata(f884_wdata), .clk(f884_clk), .rst(f884_rst), .rdata(f884_rdata));
  assign f884_clk = clk;
  assign f884_rst = rst;
  // Bindings to f884

  // f886
  logic [0:0] f886_wen;
  logic [31:0] f886_wdata;
  logic [0:0] f886_clk;
  logic [0:0] f886_rst;
  logic [31:0] f886_rdata;
  sr_buffer_32_1 f886(.wen(f886_wen), .wdata(f886_wdata), .clk(f886_clk), .rst(f886_rst), .rdata(f886_rdata));
  assign f886_clk = clk;
  assign f886_rst = rst;
  // Bindings to f886

  // f888
  logic [0:0] f888_wen;
  logic [31:0] f888_wdata;
  logic [0:0] f888_clk;
  logic [0:0] f888_rst;
  logic [31:0] f888_rdata;
  sr_buffer_32_1 f888(.wen(f888_wen), .wdata(f888_wdata), .clk(f888_clk), .rst(f888_rst), .rdata(f888_rdata));
  assign f888_clk = clk;
  assign f888_rst = rst;
  // Bindings to f888

  // f890
  logic [0:0] f890_wen;
  logic [31:0] f890_wdata;
  logic [0:0] f890_clk;
  logic [0:0] f890_rst;
  logic [31:0] f890_rdata;
  sr_buffer_32_1 f890(.wen(f890_wen), .wdata(f890_wdata), .clk(f890_clk), .rst(f890_rst), .rdata(f890_rdata));
  assign f890_clk = clk;
  assign f890_rst = rst;
  // Bindings to f890

  // f892
  logic [0:0] f892_wen;
  logic [31:0] f892_wdata;
  logic [0:0] f892_clk;
  logic [0:0] f892_rst;
  logic [31:0] f892_rdata;
  sr_buffer_32_1 f892(.wen(f892_wen), .wdata(f892_wdata), .clk(f892_clk), .rst(f892_rst), .rdata(f892_rdata));
  assign f892_clk = clk;
  assign f892_rst = rst;
  // Bindings to f892

  // f894
  logic [0:0] f894_wen;
  logic [31:0] f894_wdata;
  logic [0:0] f894_clk;
  logic [0:0] f894_rst;
  logic [31:0] f894_rdata;
  sr_buffer_32_1 f894(.wen(f894_wen), .wdata(f894_wdata), .clk(f894_clk), .rst(f894_rst), .rdata(f894_rdata));
  assign f894_clk = clk;
  assign f894_rst = rst;
  // Bindings to f894

  // f896
  logic [0:0] f896_wen;
  logic [31:0] f896_wdata;
  logic [0:0] f896_clk;
  logic [0:0] f896_rst;
  logic [31:0] f896_rdata;
  sr_buffer_32_1 f896(.wen(f896_wen), .wdata(f896_wdata), .clk(f896_clk), .rst(f896_rst), .rdata(f896_rdata));
  assign f896_clk = clk;
  assign f896_rst = rst;
  // Bindings to f896

  // f898
  logic [0:0] f898_wen;
  logic [31:0] f898_wdata;
  logic [0:0] f898_clk;
  logic [0:0] f898_rst;
  logic [31:0] f898_rdata;
  sr_buffer_32_1 f898(.wen(f898_wen), .wdata(f898_wdata), .clk(f898_clk), .rst(f898_rst), .rdata(f898_rdata));
  assign f898_clk = clk;
  assign f898_rst = rst;
  // Bindings to f898

  // f900
  logic [0:0] f900_wen;
  logic [31:0] f900_wdata;
  logic [0:0] f900_clk;
  logic [0:0] f900_rst;
  logic [31:0] f900_rdata;
  sr_buffer_32_1 f900(.wen(f900_wen), .wdata(f900_wdata), .clk(f900_clk), .rst(f900_rst), .rdata(f900_rdata));
  assign f900_clk = clk;
  assign f900_rst = rst;
  // Bindings to f900

  // f902
  logic [0:0] f902_wen;
  logic [31:0] f902_wdata;
  logic [0:0] f902_clk;
  logic [0:0] f902_rst;
  logic [31:0] f902_rdata;
  sr_buffer_32_1 f902(.wen(f902_wen), .wdata(f902_wdata), .clk(f902_clk), .rst(f902_rst), .rdata(f902_rdata));
  assign f902_clk = clk;
  assign f902_rst = rst;
  // Bindings to f902

  // f904
  logic [0:0] f904_wen;
  logic [31:0] f904_wdata;
  logic [0:0] f904_clk;
  logic [0:0] f904_rst;
  logic [31:0] f904_rdata;
  sr_buffer_32_1 f904(.wen(f904_wen), .wdata(f904_wdata), .clk(f904_clk), .rst(f904_rst), .rdata(f904_rdata));
  assign f904_clk = clk;
  assign f904_rst = rst;
  // Bindings to f904

  // f906
  logic [0:0] f906_wen;
  logic [31:0] f906_wdata;
  logic [0:0] f906_clk;
  logic [0:0] f906_rst;
  logic [31:0] f906_rdata;
  sr_buffer_32_1 f906(.wen(f906_wen), .wdata(f906_wdata), .clk(f906_clk), .rst(f906_rst), .rdata(f906_rdata));
  assign f906_clk = clk;
  assign f906_rst = rst;
  // Bindings to f906

  // f908
  logic [0:0] f908_wen;
  logic [31:0] f908_wdata;
  logic [0:0] f908_clk;
  logic [0:0] f908_rst;
  logic [31:0] f908_rdata;
  sr_buffer_32_1 f908(.wen(f908_wen), .wdata(f908_wdata), .clk(f908_clk), .rst(f908_rst), .rdata(f908_rdata));
  assign f908_clk = clk;
  assign f908_rst = rst;
  // Bindings to f908

  // f910
  logic [0:0] f910_wen;
  logic [31:0] f910_wdata;
  logic [0:0] f910_clk;
  logic [0:0] f910_rst;
  logic [31:0] f910_rdata;
  sr_buffer_32_1 f910(.wen(f910_wen), .wdata(f910_wdata), .clk(f910_clk), .rst(f910_rst), .rdata(f910_rdata));
  assign f910_clk = clk;
  assign f910_rst = rst;
  // Bindings to f910

  // f912
  logic [0:0] f912_wen;
  logic [31:0] f912_wdata;
  logic [0:0] f912_clk;
  logic [0:0] f912_rst;
  logic [31:0] f912_rdata;
  sr_buffer_32_1 f912(.wen(f912_wen), .wdata(f912_wdata), .clk(f912_clk), .rst(f912_rst), .rdata(f912_rdata));
  assign f912_clk = clk;
  assign f912_rst = rst;
  // Bindings to f912

  // f914
  logic [0:0] f914_wen;
  logic [31:0] f914_wdata;
  logic [0:0] f914_clk;
  logic [0:0] f914_rst;
  logic [31:0] f914_rdata;
  sr_buffer_32_1 f914(.wen(f914_wen), .wdata(f914_wdata), .clk(f914_clk), .rst(f914_rst), .rdata(f914_rdata));
  assign f914_clk = clk;
  assign f914_rst = rst;
  // Bindings to f914

  // f916
  logic [0:0] f916_wen;
  logic [31:0] f916_wdata;
  logic [0:0] f916_clk;
  logic [0:0] f916_rst;
  logic [31:0] f916_rdata;
  sr_buffer_32_1 f916(.wen(f916_wen), .wdata(f916_wdata), .clk(f916_clk), .rst(f916_rst), .rdata(f916_rdata));
  assign f916_clk = clk;
  assign f916_rst = rst;
  // Bindings to f916

  // f918
  logic [0:0] f918_wen;
  logic [31:0] f918_wdata;
  logic [0:0] f918_clk;
  logic [0:0] f918_rst;
  logic [31:0] f918_rdata;
  sr_buffer_32_1 f918(.wen(f918_wen), .wdata(f918_wdata), .clk(f918_clk), .rst(f918_rst), .rdata(f918_rdata));
  assign f918_clk = clk;
  assign f918_rst = rst;
  // Bindings to f918

  // f920
  logic [0:0] f920_wen;
  logic [31:0] f920_wdata;
  logic [0:0] f920_clk;
  logic [0:0] f920_rst;
  logic [31:0] f920_rdata;
  sr_buffer_32_1 f920(.wen(f920_wen), .wdata(f920_wdata), .clk(f920_clk), .rst(f920_rst), .rdata(f920_rdata));
  assign f920_clk = clk;
  assign f920_rst = rst;
  // Bindings to f920

  // f922
  logic [0:0] f922_wen;
  logic [31:0] f922_wdata;
  logic [0:0] f922_clk;
  logic [0:0] f922_rst;
  logic [31:0] f922_rdata;
  sr_buffer_32_1 f922(.wen(f922_wen), .wdata(f922_wdata), .clk(f922_clk), .rst(f922_rst), .rdata(f922_rdata));
  assign f922_clk = clk;
  assign f922_rst = rst;
  // Bindings to f922

  // f924
  logic [0:0] f924_wen;
  logic [31:0] f924_wdata;
  logic [0:0] f924_clk;
  logic [0:0] f924_rst;
  logic [31:0] f924_rdata;
  sr_buffer_32_1 f924(.wen(f924_wen), .wdata(f924_wdata), .clk(f924_clk), .rst(f924_rst), .rdata(f924_rdata));
  assign f924_clk = clk;
  assign f924_rst = rst;
  // Bindings to f924

  // f926
  logic [0:0] f926_wen;
  logic [31:0] f926_wdata;
  logic [0:0] f926_clk;
  logic [0:0] f926_rst;
  logic [31:0] f926_rdata;
  sr_buffer_32_1 f926(.wen(f926_wen), .wdata(f926_wdata), .clk(f926_clk), .rst(f926_rst), .rdata(f926_rdata));
  assign f926_clk = clk;
  assign f926_rst = rst;
  // Bindings to f926

  // f928
  logic [0:0] f928_wen;
  logic [31:0] f928_wdata;
  logic [0:0] f928_clk;
  logic [0:0] f928_rst;
  logic [31:0] f928_rdata;
  sr_buffer_32_1 f928(.wen(f928_wen), .wdata(f928_wdata), .clk(f928_clk), .rst(f928_rst), .rdata(f928_rdata));
  assign f928_clk = clk;
  assign f928_rst = rst;
  // Bindings to f928

  // f930
  logic [0:0] f930_wen;
  logic [31:0] f930_wdata;
  logic [0:0] f930_clk;
  logic [0:0] f930_rst;
  logic [31:0] f930_rdata;
  sr_buffer_32_1 f930(.wen(f930_wen), .wdata(f930_wdata), .clk(f930_clk), .rst(f930_rst), .rdata(f930_rdata));
  assign f930_clk = clk;
  assign f930_rst = rst;
  // Bindings to f930

  // f932
  logic [0:0] f932_wen;
  logic [31:0] f932_wdata;
  logic [0:0] f932_clk;
  logic [0:0] f932_rst;
  logic [31:0] f932_rdata;
  sr_buffer_32_1 f932(.wen(f932_wen), .wdata(f932_wdata), .clk(f932_clk), .rst(f932_rst), .rdata(f932_rdata));
  assign f932_clk = clk;
  assign f932_rst = rst;
  // Bindings to f932

  // f934
  logic [0:0] f934_wen;
  logic [31:0] f934_wdata;
  logic [0:0] f934_clk;
  logic [0:0] f934_rst;
  logic [31:0] f934_rdata;
  sr_buffer_32_1 f934(.wen(f934_wen), .wdata(f934_wdata), .clk(f934_clk), .rst(f934_rst), .rdata(f934_rdata));
  assign f934_clk = clk;
  assign f934_rst = rst;
  // Bindings to f934

  // f936
  logic [0:0] f936_wen;
  logic [31:0] f936_wdata;
  logic [0:0] f936_clk;
  logic [0:0] f936_rst;
  logic [31:0] f936_rdata;
  sr_buffer_32_1 f936(.wen(f936_wen), .wdata(f936_wdata), .clk(f936_clk), .rst(f936_rst), .rdata(f936_rdata));
  assign f936_clk = clk;
  assign f936_rst = rst;
  // Bindings to f936

  // f938
  logic [0:0] f938_wen;
  logic [31:0] f938_wdata;
  logic [0:0] f938_clk;
  logic [0:0] f938_rst;
  logic [31:0] f938_rdata;
  sr_buffer_32_1 f938(.wen(f938_wen), .wdata(f938_wdata), .clk(f938_clk), .rst(f938_rst), .rdata(f938_rdata));
  assign f938_clk = clk;
  assign f938_rst = rst;
  // Bindings to f938

  // f940
  logic [0:0] f940_wen;
  logic [31:0] f940_wdata;
  logic [0:0] f940_clk;
  logic [0:0] f940_rst;
  logic [31:0] f940_rdata;
  sr_buffer_32_1 f940(.wen(f940_wen), .wdata(f940_wdata), .clk(f940_clk), .rst(f940_rst), .rdata(f940_rdata));
  assign f940_clk = clk;
  assign f940_rst = rst;
  // Bindings to f940

  // f942
  logic [0:0] f942_wen;
  logic [31:0] f942_wdata;
  logic [0:0] f942_clk;
  logic [0:0] f942_rst;
  logic [31:0] f942_rdata;
  sr_buffer_32_1 f942(.wen(f942_wen), .wdata(f942_wdata), .clk(f942_clk), .rst(f942_rst), .rdata(f942_rdata));
  assign f942_clk = clk;
  assign f942_rst = rst;
  // Bindings to f942

  // f944
  logic [0:0] f944_wen;
  logic [31:0] f944_wdata;
  logic [0:0] f944_clk;
  logic [0:0] f944_rst;
  logic [31:0] f944_rdata;
  sr_buffer_32_1 f944(.wen(f944_wen), .wdata(f944_wdata), .clk(f944_clk), .rst(f944_rst), .rdata(f944_rdata));
  assign f944_clk = clk;
  assign f944_rst = rst;
  // Bindings to f944

  // f946
  logic [0:0] f946_wen;
  logic [31:0] f946_wdata;
  logic [0:0] f946_clk;
  logic [0:0] f946_rst;
  logic [31:0] f946_rdata;
  sr_buffer_32_1 f946(.wen(f946_wen), .wdata(f946_wdata), .clk(f946_clk), .rst(f946_rst), .rdata(f946_rdata));
  assign f946_clk = clk;
  assign f946_rst = rst;
  // Bindings to f946

  // f948
  logic [0:0] f948_wen;
  logic [31:0] f948_wdata;
  logic [0:0] f948_clk;
  logic [0:0] f948_rst;
  logic [31:0] f948_rdata;
  sr_buffer_32_1 f948(.wen(f948_wen), .wdata(f948_wdata), .clk(f948_clk), .rst(f948_rst), .rdata(f948_rdata));
  assign f948_clk = clk;
  assign f948_rst = rst;
  // Bindings to f948

  // f950
  logic [0:0] f950_wen;
  logic [31:0] f950_wdata;
  logic [0:0] f950_clk;
  logic [0:0] f950_rst;
  logic [31:0] f950_rdata;
  sr_buffer_32_1 f950(.wen(f950_wen), .wdata(f950_wdata), .clk(f950_clk), .rst(f950_rst), .rdata(f950_rdata));
  assign f950_clk = clk;
  assign f950_rst = rst;
  // Bindings to f950

  // f952
  logic [0:0] f952_wen;
  logic [31:0] f952_wdata;
  logic [0:0] f952_clk;
  logic [0:0] f952_rst;
  logic [31:0] f952_rdata;
  sr_buffer_32_1 f952(.wen(f952_wen), .wdata(f952_wdata), .clk(f952_clk), .rst(f952_rst), .rdata(f952_rdata));
  assign f952_clk = clk;
  assign f952_rst = rst;
  // Bindings to f952

  // f954
  logic [0:0] f954_wen;
  logic [31:0] f954_wdata;
  logic [0:0] f954_clk;
  logic [0:0] f954_rst;
  logic [31:0] f954_rdata;
  sr_buffer_32_1 f954(.wen(f954_wen), .wdata(f954_wdata), .clk(f954_clk), .rst(f954_rst), .rdata(f954_rdata));
  assign f954_clk = clk;
  assign f954_rst = rst;
  // Bindings to f954

  // f956
  logic [0:0] f956_wen;
  logic [31:0] f956_wdata;
  logic [0:0] f956_clk;
  logic [0:0] f956_rst;
  logic [31:0] f956_rdata;
  sr_buffer_32_1 f956(.wen(f956_wen), .wdata(f956_wdata), .clk(f956_clk), .rst(f956_rst), .rdata(f956_rdata));
  assign f956_clk = clk;
  assign f956_rst = rst;
  // Bindings to f956

  // f958
  logic [0:0] f958_wen;
  logic [31:0] f958_wdata;
  logic [0:0] f958_clk;
  logic [0:0] f958_rst;
  logic [31:0] f958_rdata;
  sr_buffer_32_1 f958(.wen(f958_wen), .wdata(f958_wdata), .clk(f958_clk), .rst(f958_rst), .rdata(f958_rdata));
  assign f958_clk = clk;
  assign f958_rst = rst;
  // Bindings to f958

  // f960
  logic [0:0] f960_wen;
  logic [31:0] f960_wdata;
  logic [0:0] f960_clk;
  logic [0:0] f960_rst;
  logic [31:0] f960_rdata;
  sr_buffer_32_1 f960(.wen(f960_wen), .wdata(f960_wdata), .clk(f960_clk), .rst(f960_rst), .rdata(f960_rdata));
  assign f960_clk = clk;
  assign f960_rst = rst;
  // Bindings to f960

  // f962
  logic [0:0] f962_wen;
  logic [31:0] f962_wdata;
  logic [0:0] f962_clk;
  logic [0:0] f962_rst;
  logic [31:0] f962_rdata;
  sr_buffer_32_1 f962(.wen(f962_wen), .wdata(f962_wdata), .clk(f962_clk), .rst(f962_rst), .rdata(f962_rdata));
  assign f962_clk = clk;
  assign f962_rst = rst;
  // Bindings to f962

  // f964
  logic [0:0] f964_wen;
  logic [31:0] f964_wdata;
  logic [0:0] f964_clk;
  logic [0:0] f964_rst;
  logic [31:0] f964_rdata;
  sr_buffer_32_1 f964(.wen(f964_wen), .wdata(f964_wdata), .clk(f964_clk), .rst(f964_rst), .rdata(f964_rdata));
  assign f964_clk = clk;
  assign f964_rst = rst;
  // Bindings to f964

  // f966
  logic [0:0] f966_wen;
  logic [31:0] f966_wdata;
  logic [0:0] f966_clk;
  logic [0:0] f966_rst;
  logic [31:0] f966_rdata;
  sr_buffer_32_1 f966(.wen(f966_wen), .wdata(f966_wdata), .clk(f966_clk), .rst(f966_rst), .rdata(f966_rdata));
  assign f966_clk = clk;
  assign f966_rst = rst;
  // Bindings to f966

  // f968
  logic [0:0] f968_wen;
  logic [31:0] f968_wdata;
  logic [0:0] f968_clk;
  logic [0:0] f968_rst;
  logic [31:0] f968_rdata;
  sr_buffer_32_1 f968(.wen(f968_wen), .wdata(f968_wdata), .clk(f968_clk), .rst(f968_rst), .rdata(f968_rdata));
  assign f968_clk = clk;
  assign f968_rst = rst;
  // Bindings to f968

  // f970
  logic [0:0] f970_wen;
  logic [31:0] f970_wdata;
  logic [0:0] f970_clk;
  logic [0:0] f970_rst;
  logic [31:0] f970_rdata;
  sr_buffer_32_1 f970(.wen(f970_wen), .wdata(f970_wdata), .clk(f970_clk), .rst(f970_rst), .rdata(f970_rdata));
  assign f970_clk = clk;
  assign f970_rst = rst;
  // Bindings to f970

  // f972
  logic [0:0] f972_wen;
  logic [31:0] f972_wdata;
  logic [0:0] f972_clk;
  logic [0:0] f972_rst;
  logic [31:0] f972_rdata;
  sr_buffer_32_1 f972(.wen(f972_wen), .wdata(f972_wdata), .clk(f972_clk), .rst(f972_rst), .rdata(f972_rdata));
  assign f972_clk = clk;
  assign f972_rst = rst;
  // Bindings to f972

  // f974
  logic [0:0] f974_wen;
  logic [31:0] f974_wdata;
  logic [0:0] f974_clk;
  logic [0:0] f974_rst;
  logic [31:0] f974_rdata;
  sr_buffer_32_1 f974(.wen(f974_wen), .wdata(f974_wdata), .clk(f974_clk), .rst(f974_rst), .rdata(f974_rdata));
  assign f974_clk = clk;
  assign f974_rst = rst;
  // Bindings to f974

  // f976
  logic [0:0] f976_wen;
  logic [31:0] f976_wdata;
  logic [0:0] f976_clk;
  logic [0:0] f976_rst;
  logic [31:0] f976_rdata;
  sr_buffer_32_1 f976(.wen(f976_wen), .wdata(f976_wdata), .clk(f976_clk), .rst(f976_rst), .rdata(f976_rdata));
  assign f976_clk = clk;
  assign f976_rst = rst;
  // Bindings to f976

  // f978
  logic [0:0] f978_wen;
  logic [31:0] f978_wdata;
  logic [0:0] f978_clk;
  logic [0:0] f978_rst;
  logic [31:0] f978_rdata;
  sr_buffer_32_1 f978(.wen(f978_wen), .wdata(f978_wdata), .clk(f978_clk), .rst(f978_rst), .rdata(f978_rdata));
  assign f978_clk = clk;
  assign f978_rst = rst;
  // Bindings to f978

  // f980
  logic [0:0] f980_wen;
  logic [31:0] f980_wdata;
  logic [0:0] f980_clk;
  logic [0:0] f980_rst;
  logic [31:0] f980_rdata;
  sr_buffer_32_1 f980(.wen(f980_wen), .wdata(f980_wdata), .clk(f980_clk), .rst(f980_rst), .rdata(f980_rdata));
  assign f980_clk = clk;
  assign f980_rst = rst;
  // Bindings to f980

  // f982
  logic [0:0] f982_wen;
  logic [31:0] f982_wdata;
  logic [0:0] f982_clk;
  logic [0:0] f982_rst;
  logic [31:0] f982_rdata;
  sr_buffer_32_1 f982(.wen(f982_wen), .wdata(f982_wdata), .clk(f982_clk), .rst(f982_rst), .rdata(f982_rdata));
  assign f982_clk = clk;
  assign f982_rst = rst;
  // Bindings to f982

  // f984
  logic [0:0] f984_wen;
  logic [31:0] f984_wdata;
  logic [0:0] f984_clk;
  logic [0:0] f984_rst;
  logic [31:0] f984_rdata;
  sr_buffer_32_1 f984(.wen(f984_wen), .wdata(f984_wdata), .clk(f984_clk), .rst(f984_rst), .rdata(f984_rdata));
  assign f984_clk = clk;
  assign f984_rst = rst;
  // Bindings to f984

  // f986
  logic [0:0] f986_wen;
  logic [31:0] f986_wdata;
  logic [0:0] f986_clk;
  logic [0:0] f986_rst;
  logic [31:0] f986_rdata;
  sr_buffer_32_1 f986(.wen(f986_wen), .wdata(f986_wdata), .clk(f986_clk), .rst(f986_rst), .rdata(f986_rdata));
  assign f986_clk = clk;
  assign f986_rst = rst;
  // Bindings to f986

  // f988
  logic [0:0] f988_wen;
  logic [31:0] f988_wdata;
  logic [0:0] f988_clk;
  logic [0:0] f988_rst;
  logic [31:0] f988_rdata;
  sr_buffer_32_1 f988(.wen(f988_wen), .wdata(f988_wdata), .clk(f988_clk), .rst(f988_rst), .rdata(f988_rdata));
  assign f988_clk = clk;
  assign f988_rst = rst;
  // Bindings to f988

  // f990
  logic [0:0] f990_wen;
  logic [31:0] f990_wdata;
  logic [0:0] f990_clk;
  logic [0:0] f990_rst;
  logic [31:0] f990_rdata;
  sr_buffer_32_1 f990(.wen(f990_wen), .wdata(f990_wdata), .clk(f990_clk), .rst(f990_rst), .rdata(f990_rdata));
  assign f990_clk = clk;
  assign f990_rst = rst;
  // Bindings to f990

  // f992
  logic [0:0] f992_wen;
  logic [31:0] f992_wdata;
  logic [0:0] f992_clk;
  logic [0:0] f992_rst;
  logic [31:0] f992_rdata;
  sr_buffer_32_1 f992(.wen(f992_wen), .wdata(f992_wdata), .clk(f992_clk), .rst(f992_rst), .rdata(f992_rdata));
  assign f992_clk = clk;
  assign f992_rst = rst;
  // Bindings to f992

  // f994
  logic [0:0] f994_wen;
  logic [31:0] f994_wdata;
  logic [0:0] f994_clk;
  logic [0:0] f994_rst;
  logic [31:0] f994_rdata;
  sr_buffer_32_1 f994(.wen(f994_wen), .wdata(f994_wdata), .clk(f994_clk), .rst(f994_rst), .rdata(f994_rdata));
  assign f994_clk = clk;
  assign f994_rst = rst;
  // Bindings to f994

  // f996
  logic [0:0] f996_wen;
  logic [31:0] f996_wdata;
  logic [0:0] f996_clk;
  logic [0:0] f996_rst;
  logic [31:0] f996_rdata;
  sr_buffer_32_1 f996(.wen(f996_wen), .wdata(f996_wdata), .clk(f996_clk), .rst(f996_rst), .rdata(f996_rdata));
  assign f996_clk = clk;
  assign f996_rst = rst;
  // Bindings to f996

  // f998
  logic [0:0] f998_wen;
  logic [31:0] f998_wdata;
  logic [0:0] f998_clk;
  logic [0:0] f998_rst;
  logic [31:0] f998_rdata;
  sr_buffer_32_1 f998(.wen(f998_wen), .wdata(f998_wdata), .clk(f998_clk), .rst(f998_rst), .rdata(f998_rdata));
  assign f998_clk = clk;
  assign f998_rst = rst;
  // Bindings to f998

  // f1000
  logic [0:0] f1000_wen;
  logic [31:0] f1000_wdata;
  logic [0:0] f1000_clk;
  logic [0:0] f1000_rst;
  logic [31:0] f1000_rdata;
  sr_buffer_32_1 f1000(.wen(f1000_wen), .wdata(f1000_wdata), .clk(f1000_clk), .rst(f1000_rst), .rdata(f1000_rdata));
  assign f1000_clk = clk;
  assign f1000_rst = rst;
  // Bindings to f1000

  // f1002
  logic [0:0] f1002_wen;
  logic [31:0] f1002_wdata;
  logic [0:0] f1002_clk;
  logic [0:0] f1002_rst;
  logic [31:0] f1002_rdata;
  sr_buffer_32_1 f1002(.wen(f1002_wen), .wdata(f1002_wdata), .clk(f1002_clk), .rst(f1002_rst), .rdata(f1002_rdata));
  assign f1002_clk = clk;
  assign f1002_rst = rst;
  // Bindings to f1002

  // f1004
  logic [0:0] f1004_wen;
  logic [31:0] f1004_wdata;
  logic [0:0] f1004_clk;
  logic [0:0] f1004_rst;
  logic [31:0] f1004_rdata;
  sr_buffer_32_1 f1004(.wen(f1004_wen), .wdata(f1004_wdata), .clk(f1004_clk), .rst(f1004_rst), .rdata(f1004_rdata));
  assign f1004_clk = clk;
  assign f1004_rst = rst;
  // Bindings to f1004

  // f1006
  logic [0:0] f1006_wen;
  logic [31:0] f1006_wdata;
  logic [0:0] f1006_clk;
  logic [0:0] f1006_rst;
  logic [31:0] f1006_rdata;
  sr_buffer_32_1 f1006(.wen(f1006_wen), .wdata(f1006_wdata), .clk(f1006_clk), .rst(f1006_rst), .rdata(f1006_rdata));
  assign f1006_clk = clk;
  assign f1006_rst = rst;
  // Bindings to f1006

  // f1008
  logic [0:0] f1008_wen;
  logic [31:0] f1008_wdata;
  logic [0:0] f1008_clk;
  logic [0:0] f1008_rst;
  logic [31:0] f1008_rdata;
  sr_buffer_32_1 f1008(.wen(f1008_wen), .wdata(f1008_wdata), .clk(f1008_clk), .rst(f1008_rst), .rdata(f1008_rdata));
  assign f1008_clk = clk;
  assign f1008_rst = rst;
  // Bindings to f1008

  // f1010
  logic [0:0] f1010_wen;
  logic [31:0] f1010_wdata;
  logic [0:0] f1010_clk;
  logic [0:0] f1010_rst;
  logic [31:0] f1010_rdata;
  sr_buffer_32_1 f1010(.wen(f1010_wen), .wdata(f1010_wdata), .clk(f1010_clk), .rst(f1010_rst), .rdata(f1010_rdata));
  assign f1010_clk = clk;
  assign f1010_rst = rst;
  // Bindings to f1010

  // f1012
  logic [0:0] f1012_wen;
  logic [31:0] f1012_wdata;
  logic [0:0] f1012_clk;
  logic [0:0] f1012_rst;
  logic [31:0] f1012_rdata;
  sr_buffer_32_1 f1012(.wen(f1012_wen), .wdata(f1012_wdata), .clk(f1012_clk), .rst(f1012_rst), .rdata(f1012_rdata));
  assign f1012_clk = clk;
  assign f1012_rst = rst;
  // Bindings to f1012

  // f1014
  logic [0:0] f1014_wen;
  logic [31:0] f1014_wdata;
  logic [0:0] f1014_clk;
  logic [0:0] f1014_rst;
  logic [31:0] f1014_rdata;
  sr_buffer_32_1 f1014(.wen(f1014_wen), .wdata(f1014_wdata), .clk(f1014_clk), .rst(f1014_rst), .rdata(f1014_rdata));
  assign f1014_clk = clk;
  assign f1014_rst = rst;
  // Bindings to f1014

  // f1016
  logic [0:0] f1016_wen;
  logic [31:0] f1016_wdata;
  logic [0:0] f1016_clk;
  logic [0:0] f1016_rst;
  logic [31:0] f1016_rdata;
  sr_buffer_32_1 f1016(.wen(f1016_wen), .wdata(f1016_wdata), .clk(f1016_clk), .rst(f1016_rst), .rdata(f1016_rdata));
  assign f1016_clk = clk;
  assign f1016_rst = rst;
  // Bindings to f1016

  // f1018
  logic [0:0] f1018_wen;
  logic [31:0] f1018_wdata;
  logic [0:0] f1018_clk;
  logic [0:0] f1018_rst;
  logic [31:0] f1018_rdata;
  sr_buffer_32_1 f1018(.wen(f1018_wen), .wdata(f1018_wdata), .clk(f1018_clk), .rst(f1018_rst), .rdata(f1018_rdata));
  assign f1018_clk = clk;
  assign f1018_rst = rst;
  // Bindings to f1018

  // f1020
  logic [0:0] f1020_wen;
  logic [31:0] f1020_wdata;
  logic [0:0] f1020_clk;
  logic [0:0] f1020_rst;
  logic [31:0] f1020_rdata;
  sr_buffer_32_1 f1020(.wen(f1020_wen), .wdata(f1020_wdata), .clk(f1020_clk), .rst(f1020_rst), .rdata(f1020_rdata));
  assign f1020_clk = clk;
  assign f1020_rst = rst;
  // Bindings to f1020

  // f1022
  logic [0:0] f1022_wen;
  logic [31:0] f1022_wdata;
  logic [0:0] f1022_clk;
  logic [0:0] f1022_rst;
  logic [31:0] f1022_rdata;
  sr_buffer_32_1 f1022(.wen(f1022_wen), .wdata(f1022_wdata), .clk(f1022_clk), .rst(f1022_rst), .rdata(f1022_rdata));
  assign f1022_clk = clk;
  assign f1022_rst = rst;
  // Bindings to f1022

  // f1024
  logic [0:0] f1024_wen;
  logic [31:0] f1024_wdata;
  logic [0:0] f1024_clk;
  logic [0:0] f1024_rst;
  logic [31:0] f1024_rdata;
  sr_buffer_32_1 f1024(.wen(f1024_wen), .wdata(f1024_wdata), .clk(f1024_clk), .rst(f1024_rst), .rdata(f1024_rdata));
  assign f1024_clk = clk;
  assign f1024_rst = rst;
  // Bindings to f1024

  // f1026
  logic [0:0] f1026_wen;
  logic [31:0] f1026_wdata;
  logic [0:0] f1026_clk;
  logic [0:0] f1026_rst;
  logic [31:0] f1026_rdata;
  sr_buffer_32_1 f1026(.wen(f1026_wen), .wdata(f1026_wdata), .clk(f1026_clk), .rst(f1026_rst), .rdata(f1026_rdata));
  assign f1026_clk = clk;
  assign f1026_rst = rst;
  // Bindings to f1026

  // f1028
  logic [0:0] f1028_wen;
  logic [31:0] f1028_wdata;
  logic [0:0] f1028_clk;
  logic [0:0] f1028_rst;
  logic [31:0] f1028_rdata;
  sr_buffer_32_1 f1028(.wen(f1028_wen), .wdata(f1028_wdata), .clk(f1028_clk), .rst(f1028_rst), .rdata(f1028_rdata));
  assign f1028_clk = clk;
  assign f1028_rst = rst;
  // Bindings to f1028

  // f1030
  logic [0:0] f1030_wen;
  logic [31:0] f1030_wdata;
  logic [0:0] f1030_clk;
  logic [0:0] f1030_rst;
  logic [31:0] f1030_rdata;
  sr_buffer_32_1 f1030(.wen(f1030_wen), .wdata(f1030_wdata), .clk(f1030_clk), .rst(f1030_rst), .rdata(f1030_rdata));
  assign f1030_clk = clk;
  assign f1030_rst = rst;
  // Bindings to f1030

  // f1032
  logic [0:0] f1032_wen;
  logic [31:0] f1032_wdata;
  logic [0:0] f1032_clk;
  logic [0:0] f1032_rst;
  logic [31:0] f1032_rdata;
  sr_buffer_32_1 f1032(.wen(f1032_wen), .wdata(f1032_wdata), .clk(f1032_clk), .rst(f1032_rst), .rdata(f1032_rdata));
  assign f1032_clk = clk;
  assign f1032_rst = rst;
  // Bindings to f1032

  // f1034
  logic [0:0] f1034_wen;
  logic [31:0] f1034_wdata;
  logic [0:0] f1034_clk;
  logic [0:0] f1034_rst;
  logic [31:0] f1034_rdata;
  sr_buffer_32_1 f1034(.wen(f1034_wen), .wdata(f1034_wdata), .clk(f1034_clk), .rst(f1034_rst), .rdata(f1034_rdata));
  assign f1034_clk = clk;
  assign f1034_rst = rst;
  // Bindings to f1034

  // f1036
  logic [0:0] f1036_wen;
  logic [31:0] f1036_wdata;
  logic [0:0] f1036_clk;
  logic [0:0] f1036_rst;
  logic [31:0] f1036_rdata;
  sr_buffer_32_1 f1036(.wen(f1036_wen), .wdata(f1036_wdata), .clk(f1036_clk), .rst(f1036_rst), .rdata(f1036_rdata));
  assign f1036_clk = clk;
  assign f1036_rst = rst;
  // Bindings to f1036

  // f1038
  logic [0:0] f1038_wen;
  logic [31:0] f1038_wdata;
  logic [0:0] f1038_clk;
  logic [0:0] f1038_rst;
  logic [31:0] f1038_rdata;
  sr_buffer_32_1 f1038(.wen(f1038_wen), .wdata(f1038_wdata), .clk(f1038_clk), .rst(f1038_rst), .rdata(f1038_rdata));
  assign f1038_clk = clk;
  assign f1038_rst = rst;
  // Bindings to f1038

  // f1040
  logic [0:0] f1040_wen;
  logic [31:0] f1040_wdata;
  logic [0:0] f1040_clk;
  logic [0:0] f1040_rst;
  logic [31:0] f1040_rdata;
  sr_buffer_32_1 f1040(.wen(f1040_wen), .wdata(f1040_wdata), .clk(f1040_clk), .rst(f1040_rst), .rdata(f1040_rdata));
  assign f1040_clk = clk;
  assign f1040_rst = rst;
  // Bindings to f1040

  // f1042
  logic [0:0] f1042_wen;
  logic [31:0] f1042_wdata;
  logic [0:0] f1042_clk;
  logic [0:0] f1042_rst;
  logic [31:0] f1042_rdata;
  sr_buffer_32_1 f1042(.wen(f1042_wen), .wdata(f1042_wdata), .clk(f1042_clk), .rst(f1042_rst), .rdata(f1042_rdata));
  assign f1042_clk = clk;
  assign f1042_rst = rst;
  // Bindings to f1042

  // f1044
  logic [0:0] f1044_wen;
  logic [31:0] f1044_wdata;
  logic [0:0] f1044_clk;
  logic [0:0] f1044_rst;
  logic [31:0] f1044_rdata;
  sr_buffer_32_1 f1044(.wen(f1044_wen), .wdata(f1044_wdata), .clk(f1044_clk), .rst(f1044_rst), .rdata(f1044_rdata));
  assign f1044_clk = clk;
  assign f1044_rst = rst;
  // Bindings to f1044

  // f1046
  logic [0:0] f1046_wen;
  logic [31:0] f1046_wdata;
  logic [0:0] f1046_clk;
  logic [0:0] f1046_rst;
  logic [31:0] f1046_rdata;
  sr_buffer_32_1 f1046(.wen(f1046_wen), .wdata(f1046_wdata), .clk(f1046_clk), .rst(f1046_rst), .rdata(f1046_rdata));
  assign f1046_clk = clk;
  assign f1046_rst = rst;
  // Bindings to f1046

  // f1048
  logic [0:0] f1048_wen;
  logic [31:0] f1048_wdata;
  logic [0:0] f1048_clk;
  logic [0:0] f1048_rst;
  logic [31:0] f1048_rdata;
  sr_buffer_32_1 f1048(.wen(f1048_wen), .wdata(f1048_wdata), .clk(f1048_clk), .rst(f1048_rst), .rdata(f1048_rdata));
  assign f1048_clk = clk;
  assign f1048_rst = rst;
  // Bindings to f1048

  // f1050
  logic [0:0] f1050_wen;
  logic [31:0] f1050_wdata;
  logic [0:0] f1050_clk;
  logic [0:0] f1050_rst;
  logic [31:0] f1050_rdata;
  sr_buffer_32_1 f1050(.wen(f1050_wen), .wdata(f1050_wdata), .clk(f1050_clk), .rst(f1050_rst), .rdata(f1050_rdata));
  assign f1050_clk = clk;
  assign f1050_rst = rst;
  // Bindings to f1050

  // f1052
  logic [0:0] f1052_wen;
  logic [31:0] f1052_wdata;
  logic [0:0] f1052_clk;
  logic [0:0] f1052_rst;
  logic [31:0] f1052_rdata;
  sr_buffer_32_1 f1052(.wen(f1052_wen), .wdata(f1052_wdata), .clk(f1052_clk), .rst(f1052_rst), .rdata(f1052_rdata));
  assign f1052_clk = clk;
  assign f1052_rst = rst;
  // Bindings to f1052

  // f1054
  logic [0:0] f1054_wen;
  logic [31:0] f1054_wdata;
  logic [0:0] f1054_clk;
  logic [0:0] f1054_rst;
  logic [31:0] f1054_rdata;
  sr_buffer_32_1 f1054(.wen(f1054_wen), .wdata(f1054_wdata), .clk(f1054_clk), .rst(f1054_rst), .rdata(f1054_rdata));
  assign f1054_clk = clk;
  assign f1054_rst = rst;
  // Bindings to f1054

  // f1056
  logic [0:0] f1056_wen;
  logic [31:0] f1056_wdata;
  logic [0:0] f1056_clk;
  logic [0:0] f1056_rst;
  logic [31:0] f1056_rdata;
  sr_buffer_32_1 f1056(.wen(f1056_wen), .wdata(f1056_wdata), .clk(f1056_clk), .rst(f1056_rst), .rdata(f1056_rdata));
  assign f1056_clk = clk;
  assign f1056_rst = rst;
  // Bindings to f1056

  // f1058
  logic [0:0] f1058_wen;
  logic [31:0] f1058_wdata;
  logic [0:0] f1058_clk;
  logic [0:0] f1058_rst;
  logic [31:0] f1058_rdata;
  sr_buffer_32_1 f1058(.wen(f1058_wen), .wdata(f1058_wdata), .clk(f1058_clk), .rst(f1058_rst), .rdata(f1058_rdata));
  assign f1058_clk = clk;
  assign f1058_rst = rst;
  // Bindings to f1058

  // f1060
  logic [0:0] f1060_wen;
  logic [31:0] f1060_wdata;
  logic [0:0] f1060_clk;
  logic [0:0] f1060_rst;
  logic [31:0] f1060_rdata;
  sr_buffer_32_1 f1060(.wen(f1060_wen), .wdata(f1060_wdata), .clk(f1060_clk), .rst(f1060_rst), .rdata(f1060_rdata));
  assign f1060_clk = clk;
  assign f1060_rst = rst;
  // Bindings to f1060

  // f1062
  logic [0:0] f1062_wen;
  logic [31:0] f1062_wdata;
  logic [0:0] f1062_clk;
  logic [0:0] f1062_rst;
  logic [31:0] f1062_rdata;
  sr_buffer_32_1 f1062(.wen(f1062_wen), .wdata(f1062_wdata), .clk(f1062_clk), .rst(f1062_rst), .rdata(f1062_rdata));
  assign f1062_clk = clk;
  assign f1062_rst = rst;
  // Bindings to f1062

  // f1064
  logic [0:0] f1064_wen;
  logic [31:0] f1064_wdata;
  logic [0:0] f1064_clk;
  logic [0:0] f1064_rst;
  logic [31:0] f1064_rdata;
  sr_buffer_32_1 f1064(.wen(f1064_wen), .wdata(f1064_wdata), .clk(f1064_clk), .rst(f1064_rst), .rdata(f1064_rdata));
  assign f1064_clk = clk;
  assign f1064_rst = rst;
  // Bindings to f1064

  // f1066
  logic [0:0] f1066_wen;
  logic [31:0] f1066_wdata;
  logic [0:0] f1066_clk;
  logic [0:0] f1066_rst;
  logic [31:0] f1066_rdata;
  sr_buffer_32_1 f1066(.wen(f1066_wen), .wdata(f1066_wdata), .clk(f1066_clk), .rst(f1066_rst), .rdata(f1066_rdata));
  assign f1066_clk = clk;
  assign f1066_rst = rst;
  // Bindings to f1066

  // f1068
  logic [0:0] f1068_wen;
  logic [31:0] f1068_wdata;
  logic [0:0] f1068_clk;
  logic [0:0] f1068_rst;
  logic [31:0] f1068_rdata;
  sr_buffer_32_1 f1068(.wen(f1068_wen), .wdata(f1068_wdata), .clk(f1068_clk), .rst(f1068_rst), .rdata(f1068_rdata));
  assign f1068_clk = clk;
  assign f1068_rst = rst;
  // Bindings to f1068

  // f1070
  logic [0:0] f1070_wen;
  logic [31:0] f1070_wdata;
  logic [0:0] f1070_clk;
  logic [0:0] f1070_rst;
  logic [31:0] f1070_rdata;
  sr_buffer_32_1 f1070(.wen(f1070_wen), .wdata(f1070_wdata), .clk(f1070_clk), .rst(f1070_rst), .rdata(f1070_rdata));
  assign f1070_clk = clk;
  assign f1070_rst = rst;
  // Bindings to f1070

  // f1072
  logic [0:0] f1072_wen;
  logic [31:0] f1072_wdata;
  logic [0:0] f1072_clk;
  logic [0:0] f1072_rst;
  logic [31:0] f1072_rdata;
  sr_buffer_32_1 f1072(.wen(f1072_wen), .wdata(f1072_wdata), .clk(f1072_clk), .rst(f1072_rst), .rdata(f1072_rdata));
  assign f1072_clk = clk;
  assign f1072_rst = rst;
  // Bindings to f1072

  // f1074
  logic [0:0] f1074_wen;
  logic [31:0] f1074_wdata;
  logic [0:0] f1074_clk;
  logic [0:0] f1074_rst;
  logic [31:0] f1074_rdata;
  sr_buffer_32_1 f1074(.wen(f1074_wen), .wdata(f1074_wdata), .clk(f1074_clk), .rst(f1074_rst), .rdata(f1074_rdata));
  assign f1074_clk = clk;
  assign f1074_rst = rst;
  // Bindings to f1074

  // f1076
  logic [0:0] f1076_wen;
  logic [31:0] f1076_wdata;
  logic [0:0] f1076_clk;
  logic [0:0] f1076_rst;
  logic [31:0] f1076_rdata;
  sr_buffer_32_1 f1076(.wen(f1076_wen), .wdata(f1076_wdata), .clk(f1076_clk), .rst(f1076_rst), .rdata(f1076_rdata));
  assign f1076_clk = clk;
  assign f1076_rst = rst;
  // Bindings to f1076

  // f1078
  logic [0:0] f1078_wen;
  logic [31:0] f1078_wdata;
  logic [0:0] f1078_clk;
  logic [0:0] f1078_rst;
  logic [31:0] f1078_rdata;
  sr_buffer_32_1 f1078(.wen(f1078_wen), .wdata(f1078_wdata), .clk(f1078_clk), .rst(f1078_rst), .rdata(f1078_rdata));
  assign f1078_clk = clk;
  assign f1078_rst = rst;
  // Bindings to f1078

  // f1080
  logic [0:0] f1080_wen;
  logic [31:0] f1080_wdata;
  logic [0:0] f1080_clk;
  logic [0:0] f1080_rst;
  logic [31:0] f1080_rdata;
  sr_buffer_32_1 f1080(.wen(f1080_wen), .wdata(f1080_wdata), .clk(f1080_clk), .rst(f1080_rst), .rdata(f1080_rdata));
  assign f1080_clk = clk;
  assign f1080_rst = rst;
  // Bindings to f1080

  // f1082
  logic [0:0] f1082_wen;
  logic [31:0] f1082_wdata;
  logic [0:0] f1082_clk;
  logic [0:0] f1082_rst;
  logic [31:0] f1082_rdata;
  sr_buffer_32_1 f1082(.wen(f1082_wen), .wdata(f1082_wdata), .clk(f1082_clk), .rst(f1082_rst), .rdata(f1082_rdata));
  assign f1082_clk = clk;
  assign f1082_rst = rst;
  // Bindings to f1082

  // f1084
  logic [0:0] f1084_wen;
  logic [31:0] f1084_wdata;
  logic [0:0] f1084_clk;
  logic [0:0] f1084_rst;
  logic [31:0] f1084_rdata;
  sr_buffer_32_1 f1084(.wen(f1084_wen), .wdata(f1084_wdata), .clk(f1084_clk), .rst(f1084_rst), .rdata(f1084_rdata));
  assign f1084_clk = clk;
  assign f1084_rst = rst;
  // Bindings to f1084

  // f1086
  logic [0:0] f1086_wen;
  logic [31:0] f1086_wdata;
  logic [0:0] f1086_clk;
  logic [0:0] f1086_rst;
  logic [31:0] f1086_rdata;
  sr_buffer_32_1 f1086(.wen(f1086_wen), .wdata(f1086_wdata), .clk(f1086_clk), .rst(f1086_rst), .rdata(f1086_rdata));
  assign f1086_clk = clk;
  assign f1086_rst = rst;
  // Bindings to f1086

  // f1088
  logic [0:0] f1088_wen;
  logic [31:0] f1088_wdata;
  logic [0:0] f1088_clk;
  logic [0:0] f1088_rst;
  logic [31:0] f1088_rdata;
  sr_buffer_32_1 f1088(.wen(f1088_wen), .wdata(f1088_wdata), .clk(f1088_clk), .rst(f1088_rst), .rdata(f1088_rdata));
  assign f1088_clk = clk;
  assign f1088_rst = rst;
  // Bindings to f1088

  // f1090
  logic [0:0] f1090_wen;
  logic [31:0] f1090_wdata;
  logic [0:0] f1090_clk;
  logic [0:0] f1090_rst;
  logic [31:0] f1090_rdata;
  sr_buffer_32_1 f1090(.wen(f1090_wen), .wdata(f1090_wdata), .clk(f1090_clk), .rst(f1090_rst), .rdata(f1090_rdata));
  assign f1090_clk = clk;
  assign f1090_rst = rst;
  // Bindings to f1090

  // f1092
  logic [0:0] f1092_wen;
  logic [31:0] f1092_wdata;
  logic [0:0] f1092_clk;
  logic [0:0] f1092_rst;
  logic [31:0] f1092_rdata;
  sr_buffer_32_1 f1092(.wen(f1092_wen), .wdata(f1092_wdata), .clk(f1092_clk), .rst(f1092_rst), .rdata(f1092_rdata));
  assign f1092_clk = clk;
  assign f1092_rst = rst;
  // Bindings to f1092

  // f1094
  logic [0:0] f1094_wen;
  logic [31:0] f1094_wdata;
  logic [0:0] f1094_clk;
  logic [0:0] f1094_rst;
  logic [31:0] f1094_rdata;
  sr_buffer_32_1 f1094(.wen(f1094_wen), .wdata(f1094_wdata), .clk(f1094_clk), .rst(f1094_rst), .rdata(f1094_rdata));
  assign f1094_clk = clk;
  assign f1094_rst = rst;
  // Bindings to f1094

  // f1096
  logic [0:0] f1096_wen;
  logic [31:0] f1096_wdata;
  logic [0:0] f1096_clk;
  logic [0:0] f1096_rst;
  logic [31:0] f1096_rdata;
  sr_buffer_32_1 f1096(.wen(f1096_wen), .wdata(f1096_wdata), .clk(f1096_clk), .rst(f1096_rst), .rdata(f1096_rdata));
  assign f1096_clk = clk;
  assign f1096_rst = rst;
  // Bindings to f1096

  // f1098
  logic [0:0] f1098_wen;
  logic [31:0] f1098_wdata;
  logic [0:0] f1098_clk;
  logic [0:0] f1098_rst;
  logic [31:0] f1098_rdata;
  sr_buffer_32_1 f1098(.wen(f1098_wen), .wdata(f1098_wdata), .clk(f1098_clk), .rst(f1098_rst), .rdata(f1098_rdata));
  assign f1098_clk = clk;
  assign f1098_rst = rst;
  // Bindings to f1098

  // f1100
  logic [0:0] f1100_wen;
  logic [31:0] f1100_wdata;
  logic [0:0] f1100_clk;
  logic [0:0] f1100_rst;
  logic [31:0] f1100_rdata;
  sr_buffer_32_1 f1100(.wen(f1100_wen), .wdata(f1100_wdata), .clk(f1100_clk), .rst(f1100_rst), .rdata(f1100_rdata));
  assign f1100_clk = clk;
  assign f1100_rst = rst;
  // Bindings to f1100

  // f1102
  logic [0:0] f1102_wen;
  logic [31:0] f1102_wdata;
  logic [0:0] f1102_clk;
  logic [0:0] f1102_rst;
  logic [31:0] f1102_rdata;
  sr_buffer_32_1 f1102(.wen(f1102_wen), .wdata(f1102_wdata), .clk(f1102_clk), .rst(f1102_rst), .rdata(f1102_rdata));
  assign f1102_clk = clk;
  assign f1102_rst = rst;
  // Bindings to f1102

  // f1104
  logic [0:0] f1104_wen;
  logic [31:0] f1104_wdata;
  logic [0:0] f1104_clk;
  logic [0:0] f1104_rst;
  logic [31:0] f1104_rdata;
  sr_buffer_32_1 f1104(.wen(f1104_wen), .wdata(f1104_wdata), .clk(f1104_clk), .rst(f1104_rst), .rdata(f1104_rdata));
  assign f1104_clk = clk;
  assign f1104_rst = rst;
  // Bindings to f1104

  // f1106
  logic [0:0] f1106_wen;
  logic [31:0] f1106_wdata;
  logic [0:0] f1106_clk;
  logic [0:0] f1106_rst;
  logic [31:0] f1106_rdata;
  sr_buffer_32_1 f1106(.wen(f1106_wen), .wdata(f1106_wdata), .clk(f1106_clk), .rst(f1106_rst), .rdata(f1106_rdata));
  assign f1106_clk = clk;
  assign f1106_rst = rst;
  // Bindings to f1106

  // f1108
  logic [0:0] f1108_wen;
  logic [31:0] f1108_wdata;
  logic [0:0] f1108_clk;
  logic [0:0] f1108_rst;
  logic [31:0] f1108_rdata;
  sr_buffer_32_1 f1108(.wen(f1108_wen), .wdata(f1108_wdata), .clk(f1108_clk), .rst(f1108_rst), .rdata(f1108_rdata));
  assign f1108_clk = clk;
  assign f1108_rst = rst;
  // Bindings to f1108

  // f1110
  logic [0:0] f1110_wen;
  logic [31:0] f1110_wdata;
  logic [0:0] f1110_clk;
  logic [0:0] f1110_rst;
  logic [31:0] f1110_rdata;
  sr_buffer_32_1 f1110(.wen(f1110_wen), .wdata(f1110_wdata), .clk(f1110_clk), .rst(f1110_rst), .rdata(f1110_rdata));
  assign f1110_clk = clk;
  assign f1110_rst = rst;
  // Bindings to f1110

  // f1112
  logic [0:0] f1112_wen;
  logic [31:0] f1112_wdata;
  logic [0:0] f1112_clk;
  logic [0:0] f1112_rst;
  logic [31:0] f1112_rdata;
  sr_buffer_32_1 f1112(.wen(f1112_wen), .wdata(f1112_wdata), .clk(f1112_clk), .rst(f1112_rst), .rdata(f1112_rdata));
  assign f1112_clk = clk;
  assign f1112_rst = rst;
  // Bindings to f1112

  // f1114
  logic [0:0] f1114_wen;
  logic [31:0] f1114_wdata;
  logic [0:0] f1114_clk;
  logic [0:0] f1114_rst;
  logic [31:0] f1114_rdata;
  sr_buffer_32_1 f1114(.wen(f1114_wen), .wdata(f1114_wdata), .clk(f1114_clk), .rst(f1114_rst), .rdata(f1114_rdata));
  assign f1114_clk = clk;
  assign f1114_rst = rst;
  // Bindings to f1114

  // f1116
  logic [0:0] f1116_wen;
  logic [31:0] f1116_wdata;
  logic [0:0] f1116_clk;
  logic [0:0] f1116_rst;
  logic [31:0] f1116_rdata;
  sr_buffer_32_1 f1116(.wen(f1116_wen), .wdata(f1116_wdata), .clk(f1116_clk), .rst(f1116_rst), .rdata(f1116_rdata));
  assign f1116_clk = clk;
  assign f1116_rst = rst;
  // Bindings to f1116

  // f1118
  logic [0:0] f1118_wen;
  logic [31:0] f1118_wdata;
  logic [0:0] f1118_clk;
  logic [0:0] f1118_rst;
  logic [31:0] f1118_rdata;
  sr_buffer_32_1 f1118(.wen(f1118_wen), .wdata(f1118_wdata), .clk(f1118_clk), .rst(f1118_rst), .rdata(f1118_rdata));
  assign f1118_clk = clk;
  assign f1118_rst = rst;
  // Bindings to f1118

  // f1120
  logic [0:0] f1120_wen;
  logic [31:0] f1120_wdata;
  logic [0:0] f1120_clk;
  logic [0:0] f1120_rst;
  logic [31:0] f1120_rdata;
  sr_buffer_32_1 f1120(.wen(f1120_wen), .wdata(f1120_wdata), .clk(f1120_clk), .rst(f1120_rst), .rdata(f1120_rdata));
  assign f1120_clk = clk;
  assign f1120_rst = rst;
  // Bindings to f1120

  // f1122
  logic [0:0] f1122_wen;
  logic [31:0] f1122_wdata;
  logic [0:0] f1122_clk;
  logic [0:0] f1122_rst;
  logic [31:0] f1122_rdata;
  sr_buffer_32_1 f1122(.wen(f1122_wen), .wdata(f1122_wdata), .clk(f1122_clk), .rst(f1122_rst), .rdata(f1122_rdata));
  assign f1122_clk = clk;
  assign f1122_rst = rst;
  // Bindings to f1122

  // f1124
  logic [0:0] f1124_wen;
  logic [31:0] f1124_wdata;
  logic [0:0] f1124_clk;
  logic [0:0] f1124_rst;
  logic [31:0] f1124_rdata;
  sr_buffer_32_1 f1124(.wen(f1124_wen), .wdata(f1124_wdata), .clk(f1124_clk), .rst(f1124_rst), .rdata(f1124_rdata));
  assign f1124_clk = clk;
  assign f1124_rst = rst;
  // Bindings to f1124

  // f1126
  logic [0:0] f1126_wen;
  logic [31:0] f1126_wdata;
  logic [0:0] f1126_clk;
  logic [0:0] f1126_rst;
  logic [31:0] f1126_rdata;
  sr_buffer_32_1 f1126(.wen(f1126_wen), .wdata(f1126_wdata), .clk(f1126_clk), .rst(f1126_rst), .rdata(f1126_rdata));
  assign f1126_clk = clk;
  assign f1126_rst = rst;
  // Bindings to f1126

  // f1128
  logic [0:0] f1128_wen;
  logic [31:0] f1128_wdata;
  logic [0:0] f1128_clk;
  logic [0:0] f1128_rst;
  logic [31:0] f1128_rdata;
  sr_buffer_32_1 f1128(.wen(f1128_wen), .wdata(f1128_wdata), .clk(f1128_clk), .rst(f1128_rst), .rdata(f1128_rdata));
  assign f1128_clk = clk;
  assign f1128_rst = rst;
  // Bindings to f1128

  // f1130
  logic [0:0] f1130_wen;
  logic [31:0] f1130_wdata;
  logic [0:0] f1130_clk;
  logic [0:0] f1130_rst;
  logic [31:0] f1130_rdata;
  sr_buffer_32_1 f1130(.wen(f1130_wen), .wdata(f1130_wdata), .clk(f1130_clk), .rst(f1130_rst), .rdata(f1130_rdata));
  assign f1130_clk = clk;
  assign f1130_rst = rst;
  // Bindings to f1130

  // f1132
  logic [0:0] f1132_wen;
  logic [31:0] f1132_wdata;
  logic [0:0] f1132_clk;
  logic [0:0] f1132_rst;
  logic [31:0] f1132_rdata;
  sr_buffer_32_1 f1132(.wen(f1132_wen), .wdata(f1132_wdata), .clk(f1132_clk), .rst(f1132_rst), .rdata(f1132_rdata));
  assign f1132_clk = clk;
  assign f1132_rst = rst;
  // Bindings to f1132

  // f1134
  logic [0:0] f1134_wen;
  logic [31:0] f1134_wdata;
  logic [0:0] f1134_clk;
  logic [0:0] f1134_rst;
  logic [31:0] f1134_rdata;
  sr_buffer_32_1 f1134(.wen(f1134_wen), .wdata(f1134_wdata), .clk(f1134_clk), .rst(f1134_rst), .rdata(f1134_rdata));
  assign f1134_clk = clk;
  assign f1134_rst = rst;
  // Bindings to f1134

  // f1136
  logic [0:0] f1136_wen;
  logic [31:0] f1136_wdata;
  logic [0:0] f1136_clk;
  logic [0:0] f1136_rst;
  logic [31:0] f1136_rdata;
  sr_buffer_32_1 f1136(.wen(f1136_wen), .wdata(f1136_wdata), .clk(f1136_clk), .rst(f1136_rst), .rdata(f1136_rdata));
  assign f1136_clk = clk;
  assign f1136_rst = rst;
  // Bindings to f1136

  // f1138
  logic [0:0] f1138_wen;
  logic [31:0] f1138_wdata;
  logic [0:0] f1138_clk;
  logic [0:0] f1138_rst;
  logic [31:0] f1138_rdata;
  sr_buffer_32_1 f1138(.wen(f1138_wen), .wdata(f1138_wdata), .clk(f1138_clk), .rst(f1138_rst), .rdata(f1138_rdata));
  assign f1138_clk = clk;
  assign f1138_rst = rst;
  // Bindings to f1138

  // f1140
  logic [0:0] f1140_wen;
  logic [31:0] f1140_wdata;
  logic [0:0] f1140_clk;
  logic [0:0] f1140_rst;
  logic [31:0] f1140_rdata;
  sr_buffer_32_1 f1140(.wen(f1140_wen), .wdata(f1140_wdata), .clk(f1140_clk), .rst(f1140_rst), .rdata(f1140_rdata));
  assign f1140_clk = clk;
  assign f1140_rst = rst;
  // Bindings to f1140

  // f1142
  logic [0:0] f1142_wen;
  logic [31:0] f1142_wdata;
  logic [0:0] f1142_clk;
  logic [0:0] f1142_rst;
  logic [31:0] f1142_rdata;
  sr_buffer_32_1 f1142(.wen(f1142_wen), .wdata(f1142_wdata), .clk(f1142_clk), .rst(f1142_rst), .rdata(f1142_rdata));
  assign f1142_clk = clk;
  assign f1142_rst = rst;
  // Bindings to f1142

  // f1144
  logic [0:0] f1144_wen;
  logic [31:0] f1144_wdata;
  logic [0:0] f1144_clk;
  logic [0:0] f1144_rst;
  logic [31:0] f1144_rdata;
  sr_buffer_32_1 f1144(.wen(f1144_wen), .wdata(f1144_wdata), .clk(f1144_clk), .rst(f1144_rst), .rdata(f1144_rdata));
  assign f1144_clk = clk;
  assign f1144_rst = rst;
  // Bindings to f1144

  // f1146
  logic [0:0] f1146_wen;
  logic [31:0] f1146_wdata;
  logic [0:0] f1146_clk;
  logic [0:0] f1146_rst;
  logic [31:0] f1146_rdata;
  sr_buffer_32_1 f1146(.wen(f1146_wen), .wdata(f1146_wdata), .clk(f1146_clk), .rst(f1146_rst), .rdata(f1146_rdata));
  assign f1146_clk = clk;
  assign f1146_rst = rst;
  // Bindings to f1146

  // f1148
  logic [0:0] f1148_wen;
  logic [31:0] f1148_wdata;
  logic [0:0] f1148_clk;
  logic [0:0] f1148_rst;
  logic [31:0] f1148_rdata;
  sr_buffer_32_1 f1148(.wen(f1148_wen), .wdata(f1148_wdata), .clk(f1148_clk), .rst(f1148_rst), .rdata(f1148_rdata));
  assign f1148_clk = clk;
  assign f1148_rst = rst;
  // Bindings to f1148

  // f1150
  logic [0:0] f1150_wen;
  logic [31:0] f1150_wdata;
  logic [0:0] f1150_clk;
  logic [0:0] f1150_rst;
  logic [31:0] f1150_rdata;
  sr_buffer_32_1 f1150(.wen(f1150_wen), .wdata(f1150_wdata), .clk(f1150_clk), .rst(f1150_rst), .rdata(f1150_rdata));
  assign f1150_clk = clk;
  assign f1150_rst = rst;
  // Bindings to f1150

  // f1152
  logic [0:0] f1152_wen;
  logic [31:0] f1152_wdata;
  logic [0:0] f1152_clk;
  logic [0:0] f1152_rst;
  logic [31:0] f1152_rdata;
  sr_buffer_32_1 f1152(.wen(f1152_wen), .wdata(f1152_wdata), .clk(f1152_clk), .rst(f1152_rst), .rdata(f1152_rdata));
  assign f1152_clk = clk;
  assign f1152_rst = rst;
  // Bindings to f1152

  // f1154
  logic [0:0] f1154_wen;
  logic [31:0] f1154_wdata;
  logic [0:0] f1154_clk;
  logic [0:0] f1154_rst;
  logic [31:0] f1154_rdata;
  sr_buffer_32_1 f1154(.wen(f1154_wen), .wdata(f1154_wdata), .clk(f1154_clk), .rst(f1154_rst), .rdata(f1154_rdata));
  assign f1154_clk = clk;
  assign f1154_rst = rst;
  // Bindings to f1154

  // f1156
  logic [0:0] f1156_wen;
  logic [31:0] f1156_wdata;
  logic [0:0] f1156_clk;
  logic [0:0] f1156_rst;
  logic [31:0] f1156_rdata;
  sr_buffer_32_1 f1156(.wen(f1156_wen), .wdata(f1156_wdata), .clk(f1156_clk), .rst(f1156_rst), .rdata(f1156_rdata));
  assign f1156_clk = clk;
  assign f1156_rst = rst;
  // Bindings to f1156

  // f1158
  logic [0:0] f1158_wen;
  logic [31:0] f1158_wdata;
  logic [0:0] f1158_clk;
  logic [0:0] f1158_rst;
  logic [31:0] f1158_rdata;
  sr_buffer_32_1 f1158(.wen(f1158_wen), .wdata(f1158_wdata), .clk(f1158_clk), .rst(f1158_rst), .rdata(f1158_rdata));
  assign f1158_clk = clk;
  assign f1158_rst = rst;
  // Bindings to f1158

  // f1160
  logic [0:0] f1160_wen;
  logic [31:0] f1160_wdata;
  logic [0:0] f1160_clk;
  logic [0:0] f1160_rst;
  logic [31:0] f1160_rdata;
  sr_buffer_32_1 f1160(.wen(f1160_wen), .wdata(f1160_wdata), .clk(f1160_clk), .rst(f1160_rst), .rdata(f1160_rdata));
  assign f1160_clk = clk;
  assign f1160_rst = rst;
  // Bindings to f1160

  // f1162
  logic [0:0] f1162_wen;
  logic [31:0] f1162_wdata;
  logic [0:0] f1162_clk;
  logic [0:0] f1162_rst;
  logic [31:0] f1162_rdata;
  sr_buffer_32_1 f1162(.wen(f1162_wen), .wdata(f1162_wdata), .clk(f1162_clk), .rst(f1162_rst), .rdata(f1162_rdata));
  assign f1162_clk = clk;
  assign f1162_rst = rst;
  // Bindings to f1162

  // f1164
  logic [0:0] f1164_wen;
  logic [31:0] f1164_wdata;
  logic [0:0] f1164_clk;
  logic [0:0] f1164_rst;
  logic [31:0] f1164_rdata;
  sr_buffer_32_1 f1164(.wen(f1164_wen), .wdata(f1164_wdata), .clk(f1164_clk), .rst(f1164_rst), .rdata(f1164_rdata));
  assign f1164_clk = clk;
  assign f1164_rst = rst;
  // Bindings to f1164

  // f1166
  logic [0:0] f1166_wen;
  logic [31:0] f1166_wdata;
  logic [0:0] f1166_clk;
  logic [0:0] f1166_rst;
  logic [31:0] f1166_rdata;
  sr_buffer_32_1 f1166(.wen(f1166_wen), .wdata(f1166_wdata), .clk(f1166_clk), .rst(f1166_rst), .rdata(f1166_rdata));
  assign f1166_clk = clk;
  assign f1166_rst = rst;
  // Bindings to f1166

  // f1168
  logic [0:0] f1168_wen;
  logic [31:0] f1168_wdata;
  logic [0:0] f1168_clk;
  logic [0:0] f1168_rst;
  logic [31:0] f1168_rdata;
  sr_buffer_32_1 f1168(.wen(f1168_wen), .wdata(f1168_wdata), .clk(f1168_clk), .rst(f1168_rst), .rdata(f1168_rdata));
  assign f1168_clk = clk;
  assign f1168_rst = rst;
  // Bindings to f1168

  // f1170
  logic [0:0] f1170_wen;
  logic [31:0] f1170_wdata;
  logic [0:0] f1170_clk;
  logic [0:0] f1170_rst;
  logic [31:0] f1170_rdata;
  sr_buffer_32_1 f1170(.wen(f1170_wen), .wdata(f1170_wdata), .clk(f1170_clk), .rst(f1170_rst), .rdata(f1170_rdata));
  assign f1170_clk = clk;
  assign f1170_rst = rst;
  // Bindings to f1170

  // f1172
  logic [0:0] f1172_wen;
  logic [31:0] f1172_wdata;
  logic [0:0] f1172_clk;
  logic [0:0] f1172_rst;
  logic [31:0] f1172_rdata;
  sr_buffer_32_1 f1172(.wen(f1172_wen), .wdata(f1172_wdata), .clk(f1172_clk), .rst(f1172_rst), .rdata(f1172_rdata));
  assign f1172_clk = clk;
  assign f1172_rst = rst;
  // Bindings to f1172

  // f1174
  logic [0:0] f1174_wen;
  logic [31:0] f1174_wdata;
  logic [0:0] f1174_clk;
  logic [0:0] f1174_rst;
  logic [31:0] f1174_rdata;
  sr_buffer_32_1 f1174(.wen(f1174_wen), .wdata(f1174_wdata), .clk(f1174_clk), .rst(f1174_rst), .rdata(f1174_rdata));
  assign f1174_clk = clk;
  assign f1174_rst = rst;
  // Bindings to f1174

  // f1176
  logic [0:0] f1176_wen;
  logic [31:0] f1176_wdata;
  logic [0:0] f1176_clk;
  logic [0:0] f1176_rst;
  logic [31:0] f1176_rdata;
  sr_buffer_32_1 f1176(.wen(f1176_wen), .wdata(f1176_wdata), .clk(f1176_clk), .rst(f1176_rst), .rdata(f1176_rdata));
  assign f1176_clk = clk;
  assign f1176_rst = rst;
  // Bindings to f1176

  // f1178
  logic [0:0] f1178_wen;
  logic [31:0] f1178_wdata;
  logic [0:0] f1178_clk;
  logic [0:0] f1178_rst;
  logic [31:0] f1178_rdata;
  sr_buffer_32_1 f1178(.wen(f1178_wen), .wdata(f1178_wdata), .clk(f1178_clk), .rst(f1178_rst), .rdata(f1178_rdata));
  assign f1178_clk = clk;
  assign f1178_rst = rst;
  // Bindings to f1178

  // f1180
  logic [0:0] f1180_wen;
  logic [31:0] f1180_wdata;
  logic [0:0] f1180_clk;
  logic [0:0] f1180_rst;
  logic [31:0] f1180_rdata;
  sr_buffer_32_1 f1180(.wen(f1180_wen), .wdata(f1180_wdata), .clk(f1180_clk), .rst(f1180_rst), .rdata(f1180_rdata));
  assign f1180_clk = clk;
  assign f1180_rst = rst;
  // Bindings to f1180

  // f1182
  logic [0:0] f1182_wen;
  logic [31:0] f1182_wdata;
  logic [0:0] f1182_clk;
  logic [0:0] f1182_rst;
  logic [31:0] f1182_rdata;
  sr_buffer_32_1 f1182(.wen(f1182_wen), .wdata(f1182_wdata), .clk(f1182_clk), .rst(f1182_rst), .rdata(f1182_rdata));
  assign f1182_clk = clk;
  assign f1182_rst = rst;
  // Bindings to f1182

  // f1184
  logic [0:0] f1184_wen;
  logic [31:0] f1184_wdata;
  logic [0:0] f1184_clk;
  logic [0:0] f1184_rst;
  logic [31:0] f1184_rdata;
  sr_buffer_32_1 f1184(.wen(f1184_wen), .wdata(f1184_wdata), .clk(f1184_clk), .rst(f1184_rst), .rdata(f1184_rdata));
  assign f1184_clk = clk;
  assign f1184_rst = rst;
  // Bindings to f1184

  // f1186
  logic [0:0] f1186_wen;
  logic [31:0] f1186_wdata;
  logic [0:0] f1186_clk;
  logic [0:0] f1186_rst;
  logic [31:0] f1186_rdata;
  sr_buffer_32_1 f1186(.wen(f1186_wen), .wdata(f1186_wdata), .clk(f1186_clk), .rst(f1186_rst), .rdata(f1186_rdata));
  assign f1186_clk = clk;
  assign f1186_rst = rst;
  // Bindings to f1186

  // f1188
  logic [0:0] f1188_wen;
  logic [31:0] f1188_wdata;
  logic [0:0] f1188_clk;
  logic [0:0] f1188_rst;
  logic [31:0] f1188_rdata;
  sr_buffer_32_1 f1188(.wen(f1188_wen), .wdata(f1188_wdata), .clk(f1188_clk), .rst(f1188_rst), .rdata(f1188_rdata));
  assign f1188_clk = clk;
  assign f1188_rst = rst;
  // Bindings to f1188

  // f1190
  logic [0:0] f1190_wen;
  logic [31:0] f1190_wdata;
  logic [0:0] f1190_clk;
  logic [0:0] f1190_rst;
  logic [31:0] f1190_rdata;
  sr_buffer_32_1 f1190(.wen(f1190_wen), .wdata(f1190_wdata), .clk(f1190_clk), .rst(f1190_rst), .rdata(f1190_rdata));
  assign f1190_clk = clk;
  assign f1190_rst = rst;
  // Bindings to f1190

  // f1192
  logic [0:0] f1192_wen;
  logic [31:0] f1192_wdata;
  logic [0:0] f1192_clk;
  logic [0:0] f1192_rst;
  logic [31:0] f1192_rdata;
  sr_buffer_32_1 f1192(.wen(f1192_wen), .wdata(f1192_wdata), .clk(f1192_clk), .rst(f1192_rst), .rdata(f1192_rdata));
  assign f1192_clk = clk;
  assign f1192_rst = rst;
  // Bindings to f1192

  // f1194
  logic [0:0] f1194_wen;
  logic [31:0] f1194_wdata;
  logic [0:0] f1194_clk;
  logic [0:0] f1194_rst;
  logic [31:0] f1194_rdata;
  sr_buffer_32_1 f1194(.wen(f1194_wen), .wdata(f1194_wdata), .clk(f1194_clk), .rst(f1194_rst), .rdata(f1194_rdata));
  assign f1194_clk = clk;
  assign f1194_rst = rst;
  // Bindings to f1194

  // f1196
  logic [0:0] f1196_wen;
  logic [31:0] f1196_wdata;
  logic [0:0] f1196_clk;
  logic [0:0] f1196_rst;
  logic [31:0] f1196_rdata;
  sr_buffer_32_1 f1196(.wen(f1196_wen), .wdata(f1196_wdata), .clk(f1196_clk), .rst(f1196_rst), .rdata(f1196_rdata));
  assign f1196_clk = clk;
  assign f1196_rst = rst;
  // Bindings to f1196

  // f1198
  logic [0:0] f1198_wen;
  logic [31:0] f1198_wdata;
  logic [0:0] f1198_clk;
  logic [0:0] f1198_rst;
  logic [31:0] f1198_rdata;
  sr_buffer_32_1 f1198(.wen(f1198_wen), .wdata(f1198_wdata), .clk(f1198_clk), .rst(f1198_rst), .rdata(f1198_rdata));
  assign f1198_clk = clk;
  assign f1198_rst = rst;
  // Bindings to f1198

  // f1200
  logic [0:0] f1200_wen;
  logic [31:0] f1200_wdata;
  logic [0:0] f1200_clk;
  logic [0:0] f1200_rst;
  logic [31:0] f1200_rdata;
  sr_buffer_32_1 f1200(.wen(f1200_wen), .wdata(f1200_wdata), .clk(f1200_clk), .rst(f1200_rst), .rdata(f1200_rdata));
  assign f1200_clk = clk;
  assign f1200_rst = rst;
  // Bindings to f1200

  // f1202
  logic [0:0] f1202_wen;
  logic [31:0] f1202_wdata;
  logic [0:0] f1202_clk;
  logic [0:0] f1202_rst;
  logic [31:0] f1202_rdata;
  sr_buffer_32_1 f1202(.wen(f1202_wen), .wdata(f1202_wdata), .clk(f1202_clk), .rst(f1202_rst), .rdata(f1202_rdata));
  assign f1202_clk = clk;
  assign f1202_rst = rst;
  // Bindings to f1202

  // f1204
  logic [0:0] f1204_wen;
  logic [31:0] f1204_wdata;
  logic [0:0] f1204_clk;
  logic [0:0] f1204_rst;
  logic [31:0] f1204_rdata;
  sr_buffer_32_1 f1204(.wen(f1204_wen), .wdata(f1204_wdata), .clk(f1204_clk), .rst(f1204_rst), .rdata(f1204_rdata));
  assign f1204_clk = clk;
  assign f1204_rst = rst;
  // Bindings to f1204

  // f1206
  logic [0:0] f1206_wen;
  logic [31:0] f1206_wdata;
  logic [0:0] f1206_clk;
  logic [0:0] f1206_rst;
  logic [31:0] f1206_rdata;
  sr_buffer_32_1 f1206(.wen(f1206_wen), .wdata(f1206_wdata), .clk(f1206_clk), .rst(f1206_rst), .rdata(f1206_rdata));
  assign f1206_clk = clk;
  assign f1206_rst = rst;
  // Bindings to f1206

  // f1208
  logic [0:0] f1208_wen;
  logic [31:0] f1208_wdata;
  logic [0:0] f1208_clk;
  logic [0:0] f1208_rst;
  logic [31:0] f1208_rdata;
  sr_buffer_32_1 f1208(.wen(f1208_wen), .wdata(f1208_wdata), .clk(f1208_clk), .rst(f1208_rst), .rdata(f1208_rdata));
  assign f1208_clk = clk;
  assign f1208_rst = rst;
  // Bindings to f1208

  // f1210
  logic [0:0] f1210_wen;
  logic [31:0] f1210_wdata;
  logic [0:0] f1210_clk;
  logic [0:0] f1210_rst;
  logic [31:0] f1210_rdata;
  sr_buffer_32_1 f1210(.wen(f1210_wen), .wdata(f1210_wdata), .clk(f1210_clk), .rst(f1210_rst), .rdata(f1210_rdata));
  assign f1210_clk = clk;
  assign f1210_rst = rst;
  // Bindings to f1210

  // f1212
  logic [0:0] f1212_wen;
  logic [31:0] f1212_wdata;
  logic [0:0] f1212_clk;
  logic [0:0] f1212_rst;
  logic [31:0] f1212_rdata;
  sr_buffer_32_1 f1212(.wen(f1212_wen), .wdata(f1212_wdata), .clk(f1212_clk), .rst(f1212_rst), .rdata(f1212_rdata));
  assign f1212_clk = clk;
  assign f1212_rst = rst;
  // Bindings to f1212

  // f1214
  logic [0:0] f1214_wen;
  logic [31:0] f1214_wdata;
  logic [0:0] f1214_clk;
  logic [0:0] f1214_rst;
  logic [31:0] f1214_rdata;
  sr_buffer_32_1 f1214(.wen(f1214_wen), .wdata(f1214_wdata), .clk(f1214_clk), .rst(f1214_rst), .rdata(f1214_rdata));
  assign f1214_clk = clk;
  assign f1214_rst = rst;
  // Bindings to f1214

  // f1216
  logic [0:0] f1216_wen;
  logic [31:0] f1216_wdata;
  logic [0:0] f1216_clk;
  logic [0:0] f1216_rst;
  logic [31:0] f1216_rdata;
  sr_buffer_32_1 f1216(.wen(f1216_wen), .wdata(f1216_wdata), .clk(f1216_clk), .rst(f1216_rst), .rdata(f1216_rdata));
  assign f1216_clk = clk;
  assign f1216_rst = rst;
  // Bindings to f1216

  // f1218
  logic [0:0] f1218_wen;
  logic [31:0] f1218_wdata;
  logic [0:0] f1218_clk;
  logic [0:0] f1218_rst;
  logic [31:0] f1218_rdata;
  sr_buffer_32_1 f1218(.wen(f1218_wen), .wdata(f1218_wdata), .clk(f1218_clk), .rst(f1218_rst), .rdata(f1218_rdata));
  assign f1218_clk = clk;
  assign f1218_rst = rst;
  // Bindings to f1218

  // f1220
  logic [0:0] f1220_wen;
  logic [31:0] f1220_wdata;
  logic [0:0] f1220_clk;
  logic [0:0] f1220_rst;
  logic [31:0] f1220_rdata;
  sr_buffer_32_1 f1220(.wen(f1220_wen), .wdata(f1220_wdata), .clk(f1220_clk), .rst(f1220_rst), .rdata(f1220_rdata));
  assign f1220_clk = clk;
  assign f1220_rst = rst;
  // Bindings to f1220

  // f1222
  logic [0:0] f1222_wen;
  logic [31:0] f1222_wdata;
  logic [0:0] f1222_clk;
  logic [0:0] f1222_rst;
  logic [31:0] f1222_rdata;
  sr_buffer_32_1 f1222(.wen(f1222_wen), .wdata(f1222_wdata), .clk(f1222_clk), .rst(f1222_rst), .rdata(f1222_rdata));
  assign f1222_clk = clk;
  assign f1222_rst = rst;
  // Bindings to f1222

  // f1224
  logic [0:0] f1224_wen;
  logic [31:0] f1224_wdata;
  logic [0:0] f1224_clk;
  logic [0:0] f1224_rst;
  logic [31:0] f1224_rdata;
  sr_buffer_32_1 f1224(.wen(f1224_wen), .wdata(f1224_wdata), .clk(f1224_clk), .rst(f1224_rst), .rdata(f1224_rdata));
  assign f1224_clk = clk;
  assign f1224_rst = rst;
  // Bindings to f1224

  // f1226
  logic [0:0] f1226_wen;
  logic [31:0] f1226_wdata;
  logic [0:0] f1226_clk;
  logic [0:0] f1226_rst;
  logic [31:0] f1226_rdata;
  sr_buffer_32_1 f1226(.wen(f1226_wen), .wdata(f1226_wdata), .clk(f1226_clk), .rst(f1226_rst), .rdata(f1226_rdata));
  assign f1226_clk = clk;
  assign f1226_rst = rst;
  // Bindings to f1226

  // f1228
  logic [0:0] f1228_wen;
  logic [31:0] f1228_wdata;
  logic [0:0] f1228_clk;
  logic [0:0] f1228_rst;
  logic [31:0] f1228_rdata;
  sr_buffer_32_1 f1228(.wen(f1228_wen), .wdata(f1228_wdata), .clk(f1228_clk), .rst(f1228_rst), .rdata(f1228_rdata));
  assign f1228_clk = clk;
  assign f1228_rst = rst;
  // Bindings to f1228

  // f1230
  logic [0:0] f1230_wen;
  logic [31:0] f1230_wdata;
  logic [0:0] f1230_clk;
  logic [0:0] f1230_rst;
  logic [31:0] f1230_rdata;
  sr_buffer_32_1 f1230(.wen(f1230_wen), .wdata(f1230_wdata), .clk(f1230_clk), .rst(f1230_rst), .rdata(f1230_rdata));
  assign f1230_clk = clk;
  assign f1230_rst = rst;
  // Bindings to f1230

  // f1232
  logic [0:0] f1232_wen;
  logic [31:0] f1232_wdata;
  logic [0:0] f1232_clk;
  logic [0:0] f1232_rst;
  logic [31:0] f1232_rdata;
  sr_buffer_32_1 f1232(.wen(f1232_wen), .wdata(f1232_wdata), .clk(f1232_clk), .rst(f1232_rst), .rdata(f1232_rdata));
  assign f1232_clk = clk;
  assign f1232_rst = rst;
  // Bindings to f1232

  // f1234
  logic [0:0] f1234_wen;
  logic [31:0] f1234_wdata;
  logic [0:0] f1234_clk;
  logic [0:0] f1234_rst;
  logic [31:0] f1234_rdata;
  sr_buffer_32_1 f1234(.wen(f1234_wen), .wdata(f1234_wdata), .clk(f1234_clk), .rst(f1234_rst), .rdata(f1234_rdata));
  assign f1234_clk = clk;
  assign f1234_rst = rst;
  // Bindings to f1234

  // f1236
  logic [0:0] f1236_wen;
  logic [31:0] f1236_wdata;
  logic [0:0] f1236_clk;
  logic [0:0] f1236_rst;
  logic [31:0] f1236_rdata;
  sr_buffer_32_1 f1236(.wen(f1236_wen), .wdata(f1236_wdata), .clk(f1236_clk), .rst(f1236_rst), .rdata(f1236_rdata));
  assign f1236_clk = clk;
  assign f1236_rst = rst;
  // Bindings to f1236

  // f1238
  logic [0:0] f1238_wen;
  logic [31:0] f1238_wdata;
  logic [0:0] f1238_clk;
  logic [0:0] f1238_rst;
  logic [31:0] f1238_rdata;
  sr_buffer_32_1 f1238(.wen(f1238_wen), .wdata(f1238_wdata), .clk(f1238_clk), .rst(f1238_rst), .rdata(f1238_rdata));
  assign f1238_clk = clk;
  assign f1238_rst = rst;
  // Bindings to f1238

  // f1240
  logic [0:0] f1240_wen;
  logic [31:0] f1240_wdata;
  logic [0:0] f1240_clk;
  logic [0:0] f1240_rst;
  logic [31:0] f1240_rdata;
  sr_buffer_32_1 f1240(.wen(f1240_wen), .wdata(f1240_wdata), .clk(f1240_clk), .rst(f1240_rst), .rdata(f1240_rdata));
  assign f1240_clk = clk;
  assign f1240_rst = rst;
  // Bindings to f1240

  // f1242
  logic [0:0] f1242_wen;
  logic [31:0] f1242_wdata;
  logic [0:0] f1242_clk;
  logic [0:0] f1242_rst;
  logic [31:0] f1242_rdata;
  sr_buffer_32_1 f1242(.wen(f1242_wen), .wdata(f1242_wdata), .clk(f1242_clk), .rst(f1242_rst), .rdata(f1242_rdata));
  assign f1242_clk = clk;
  assign f1242_rst = rst;
  // Bindings to f1242

  // f1244
  logic [0:0] f1244_wen;
  logic [31:0] f1244_wdata;
  logic [0:0] f1244_clk;
  logic [0:0] f1244_rst;
  logic [31:0] f1244_rdata;
  sr_buffer_32_1 f1244(.wen(f1244_wen), .wdata(f1244_wdata), .clk(f1244_clk), .rst(f1244_rst), .rdata(f1244_rdata));
  assign f1244_clk = clk;
  assign f1244_rst = rst;
  // Bindings to f1244

  // f1246
  logic [0:0] f1246_wen;
  logic [31:0] f1246_wdata;
  logic [0:0] f1246_clk;
  logic [0:0] f1246_rst;
  logic [31:0] f1246_rdata;
  sr_buffer_32_1 f1246(.wen(f1246_wen), .wdata(f1246_wdata), .clk(f1246_clk), .rst(f1246_rst), .rdata(f1246_rdata));
  assign f1246_clk = clk;
  assign f1246_rst = rst;
  // Bindings to f1246

  // f1248
  logic [0:0] f1248_wen;
  logic [31:0] f1248_wdata;
  logic [0:0] f1248_clk;
  logic [0:0] f1248_rst;
  logic [31:0] f1248_rdata;
  sr_buffer_32_1 f1248(.wen(f1248_wen), .wdata(f1248_wdata), .clk(f1248_clk), .rst(f1248_rst), .rdata(f1248_rdata));
  assign f1248_clk = clk;
  assign f1248_rst = rst;
  // Bindings to f1248

  // f1250
  logic [0:0] f1250_wen;
  logic [31:0] f1250_wdata;
  logic [0:0] f1250_clk;
  logic [0:0] f1250_rst;
  logic [31:0] f1250_rdata;
  sr_buffer_32_1 f1250(.wen(f1250_wen), .wdata(f1250_wdata), .clk(f1250_clk), .rst(f1250_rst), .rdata(f1250_rdata));
  assign f1250_clk = clk;
  assign f1250_rst = rst;
  // Bindings to f1250

  // f1252
  logic [0:0] f1252_wen;
  logic [31:0] f1252_wdata;
  logic [0:0] f1252_clk;
  logic [0:0] f1252_rst;
  logic [31:0] f1252_rdata;
  sr_buffer_32_1 f1252(.wen(f1252_wen), .wdata(f1252_wdata), .clk(f1252_clk), .rst(f1252_rst), .rdata(f1252_rdata));
  assign f1252_clk = clk;
  assign f1252_rst = rst;
  // Bindings to f1252

  // f1254
  logic [0:0] f1254_wen;
  logic [31:0] f1254_wdata;
  logic [0:0] f1254_clk;
  logic [0:0] f1254_rst;
  logic [31:0] f1254_rdata;
  sr_buffer_32_1 f1254(.wen(f1254_wen), .wdata(f1254_wdata), .clk(f1254_clk), .rst(f1254_rst), .rdata(f1254_rdata));
  assign f1254_clk = clk;
  assign f1254_rst = rst;
  // Bindings to f1254

  // f1256
  logic [0:0] f1256_wen;
  logic [31:0] f1256_wdata;
  logic [0:0] f1256_clk;
  logic [0:0] f1256_rst;
  logic [31:0] f1256_rdata;
  sr_buffer_32_1 f1256(.wen(f1256_wen), .wdata(f1256_wdata), .clk(f1256_clk), .rst(f1256_rst), .rdata(f1256_rdata));
  assign f1256_clk = clk;
  assign f1256_rst = rst;
  // Bindings to f1256

  // f1258
  logic [0:0] f1258_wen;
  logic [31:0] f1258_wdata;
  logic [0:0] f1258_clk;
  logic [0:0] f1258_rst;
  logic [31:0] f1258_rdata;
  sr_buffer_32_1 f1258(.wen(f1258_wen), .wdata(f1258_wdata), .clk(f1258_clk), .rst(f1258_rst), .rdata(f1258_rdata));
  assign f1258_clk = clk;
  assign f1258_rst = rst;
  // Bindings to f1258

  // f1260
  logic [0:0] f1260_wen;
  logic [31:0] f1260_wdata;
  logic [0:0] f1260_clk;
  logic [0:0] f1260_rst;
  logic [31:0] f1260_rdata;
  sr_buffer_32_1 f1260(.wen(f1260_wen), .wdata(f1260_wdata), .clk(f1260_clk), .rst(f1260_rst), .rdata(f1260_rdata));
  assign f1260_clk = clk;
  assign f1260_rst = rst;
  // Bindings to f1260

  // f1262
  logic [0:0] f1262_wen;
  logic [31:0] f1262_wdata;
  logic [0:0] f1262_clk;
  logic [0:0] f1262_rst;
  logic [31:0] f1262_rdata;
  sr_buffer_32_1 f1262(.wen(f1262_wen), .wdata(f1262_wdata), .clk(f1262_clk), .rst(f1262_rst), .rdata(f1262_rdata));
  assign f1262_clk = clk;
  assign f1262_rst = rst;
  // Bindings to f1262

  // f1264
  logic [0:0] f1264_wen;
  logic [31:0] f1264_wdata;
  logic [0:0] f1264_clk;
  logic [0:0] f1264_rst;
  logic [31:0] f1264_rdata;
  sr_buffer_32_1 f1264(.wen(f1264_wen), .wdata(f1264_wdata), .clk(f1264_clk), .rst(f1264_rst), .rdata(f1264_rdata));
  assign f1264_clk = clk;
  assign f1264_rst = rst;
  // Bindings to f1264

  // f1266
  logic [0:0] f1266_wen;
  logic [31:0] f1266_wdata;
  logic [0:0] f1266_clk;
  logic [0:0] f1266_rst;
  logic [31:0] f1266_rdata;
  sr_buffer_32_1 f1266(.wen(f1266_wen), .wdata(f1266_wdata), .clk(f1266_clk), .rst(f1266_rst), .rdata(f1266_rdata));
  assign f1266_clk = clk;
  assign f1266_rst = rst;
  // Bindings to f1266

  // f1268
  logic [0:0] f1268_wen;
  logic [31:0] f1268_wdata;
  logic [0:0] f1268_clk;
  logic [0:0] f1268_rst;
  logic [31:0] f1268_rdata;
  sr_buffer_32_1 f1268(.wen(f1268_wen), .wdata(f1268_wdata), .clk(f1268_clk), .rst(f1268_rst), .rdata(f1268_rdata));
  assign f1268_clk = clk;
  assign f1268_rst = rst;
  // Bindings to f1268

  // f1270
  logic [0:0] f1270_wen;
  logic [31:0] f1270_wdata;
  logic [0:0] f1270_clk;
  logic [0:0] f1270_rst;
  logic [31:0] f1270_rdata;
  sr_buffer_32_1 f1270(.wen(f1270_wen), .wdata(f1270_wdata), .clk(f1270_clk), .rst(f1270_rst), .rdata(f1270_rdata));
  assign f1270_clk = clk;
  assign f1270_rst = rst;
  // Bindings to f1270

  // f1272
  logic [0:0] f1272_wen;
  logic [31:0] f1272_wdata;
  logic [0:0] f1272_clk;
  logic [0:0] f1272_rst;
  logic [31:0] f1272_rdata;
  sr_buffer_32_1 f1272(.wen(f1272_wen), .wdata(f1272_wdata), .clk(f1272_clk), .rst(f1272_rst), .rdata(f1272_rdata));
  assign f1272_clk = clk;
  assign f1272_rst = rst;
  // Bindings to f1272

  // f1274
  logic [0:0] f1274_wen;
  logic [31:0] f1274_wdata;
  logic [0:0] f1274_clk;
  logic [0:0] f1274_rst;
  logic [31:0] f1274_rdata;
  sr_buffer_32_1 f1274(.wen(f1274_wen), .wdata(f1274_wdata), .clk(f1274_clk), .rst(f1274_rst), .rdata(f1274_rdata));
  assign f1274_clk = clk;
  assign f1274_rst = rst;
  // Bindings to f1274

  // f1276
  logic [0:0] f1276_wen;
  logic [31:0] f1276_wdata;
  logic [0:0] f1276_clk;
  logic [0:0] f1276_rst;
  logic [31:0] f1276_rdata;
  sr_buffer_32_1 f1276(.wen(f1276_wen), .wdata(f1276_wdata), .clk(f1276_clk), .rst(f1276_rst), .rdata(f1276_rdata));
  assign f1276_clk = clk;
  assign f1276_rst = rst;
  // Bindings to f1276

  // f1278
  logic [0:0] f1278_wen;
  logic [31:0] f1278_wdata;
  logic [0:0] f1278_clk;
  logic [0:0] f1278_rst;
  logic [31:0] f1278_rdata;
  sr_buffer_32_1 f1278(.wen(f1278_wen), .wdata(f1278_wdata), .clk(f1278_clk), .rst(f1278_rst), .rdata(f1278_rdata));
  assign f1278_clk = clk;
  assign f1278_rst = rst;
  // Bindings to f1278

  // f1280
  logic [0:0] f1280_wen;
  logic [31:0] f1280_wdata;
  logic [0:0] f1280_clk;
  logic [0:0] f1280_rst;
  logic [31:0] f1280_rdata;
  sr_buffer_32_1 f1280(.wen(f1280_wen), .wdata(f1280_wdata), .clk(f1280_clk), .rst(f1280_rst), .rdata(f1280_rdata));
  assign f1280_clk = clk;
  assign f1280_rst = rst;
  // Bindings to f1280

  // f1282
  logic [0:0] f1282_wen;
  logic [31:0] f1282_wdata;
  logic [0:0] f1282_clk;
  logic [0:0] f1282_rst;
  logic [31:0] f1282_rdata;
  sr_buffer_32_1 f1282(.wen(f1282_wen), .wdata(f1282_wdata), .clk(f1282_clk), .rst(f1282_rst), .rdata(f1282_rdata));
  assign f1282_clk = clk;
  assign f1282_rst = rst;
  // Bindings to f1282

  // f1284
  logic [0:0] f1284_wen;
  logic [31:0] f1284_wdata;
  logic [0:0] f1284_clk;
  logic [0:0] f1284_rst;
  logic [31:0] f1284_rdata;
  sr_buffer_32_1 f1284(.wen(f1284_wen), .wdata(f1284_wdata), .clk(f1284_clk), .rst(f1284_rst), .rdata(f1284_rdata));
  assign f1284_clk = clk;
  assign f1284_rst = rst;
  // Bindings to f1284

  // f1286
  logic [0:0] f1286_wen;
  logic [31:0] f1286_wdata;
  logic [0:0] f1286_clk;
  logic [0:0] f1286_rst;
  logic [31:0] f1286_rdata;
  sr_buffer_32_1 f1286(.wen(f1286_wen), .wdata(f1286_wdata), .clk(f1286_clk), .rst(f1286_rst), .rdata(f1286_rdata));
  assign f1286_clk = clk;
  assign f1286_rst = rst;
  // Bindings to f1286

  // f1288
  logic [0:0] f1288_wen;
  logic [31:0] f1288_wdata;
  logic [0:0] f1288_clk;
  logic [0:0] f1288_rst;
  logic [31:0] f1288_rdata;
  sr_buffer_32_1 f1288(.wen(f1288_wen), .wdata(f1288_wdata), .clk(f1288_clk), .rst(f1288_rst), .rdata(f1288_rdata));
  assign f1288_clk = clk;
  assign f1288_rst = rst;
  // Bindings to f1288

  // f1290
  logic [0:0] f1290_wen;
  logic [31:0] f1290_wdata;
  logic [0:0] f1290_clk;
  logic [0:0] f1290_rst;
  logic [31:0] f1290_rdata;
  sr_buffer_32_1 f1290(.wen(f1290_wen), .wdata(f1290_wdata), .clk(f1290_clk), .rst(f1290_rst), .rdata(f1290_rdata));
  assign f1290_clk = clk;
  assign f1290_rst = rst;
  // Bindings to f1290

  // f1292
  logic [0:0] f1292_wen;
  logic [31:0] f1292_wdata;
  logic [0:0] f1292_clk;
  logic [0:0] f1292_rst;
  logic [31:0] f1292_rdata;
  sr_buffer_32_1 f1292(.wen(f1292_wen), .wdata(f1292_wdata), .clk(f1292_clk), .rst(f1292_rst), .rdata(f1292_rdata));
  assign f1292_clk = clk;
  assign f1292_rst = rst;
  // Bindings to f1292

  // f1294
  logic [0:0] f1294_wen;
  logic [31:0] f1294_wdata;
  logic [0:0] f1294_clk;
  logic [0:0] f1294_rst;
  logic [31:0] f1294_rdata;
  sr_buffer_32_1 f1294(.wen(f1294_wen), .wdata(f1294_wdata), .clk(f1294_clk), .rst(f1294_rst), .rdata(f1294_rdata));
  assign f1294_clk = clk;
  assign f1294_rst = rst;
  // Bindings to f1294

  // f1296
  logic [0:0] f1296_wen;
  logic [31:0] f1296_wdata;
  logic [0:0] f1296_clk;
  logic [0:0] f1296_rst;
  logic [31:0] f1296_rdata;
  sr_buffer_32_1 f1296(.wen(f1296_wen), .wdata(f1296_wdata), .clk(f1296_clk), .rst(f1296_rst), .rdata(f1296_rdata));
  assign f1296_clk = clk;
  assign f1296_rst = rst;
  // Bindings to f1296

  // f1298
  logic [0:0] f1298_wen;
  logic [31:0] f1298_wdata;
  logic [0:0] f1298_clk;
  logic [0:0] f1298_rst;
  logic [31:0] f1298_rdata;
  sr_buffer_32_1 f1298(.wen(f1298_wen), .wdata(f1298_wdata), .clk(f1298_clk), .rst(f1298_rst), .rdata(f1298_rdata));
  assign f1298_clk = clk;
  assign f1298_rst = rst;
  // Bindings to f1298

  // f1300
  logic [0:0] f1300_wen;
  logic [31:0] f1300_wdata;
  logic [0:0] f1300_clk;
  logic [0:0] f1300_rst;
  logic [31:0] f1300_rdata;
  sr_buffer_32_1 f1300(.wen(f1300_wen), .wdata(f1300_wdata), .clk(f1300_clk), .rst(f1300_rst), .rdata(f1300_rdata));
  assign f1300_clk = clk;
  assign f1300_rst = rst;
  // Bindings to f1300

  // f1302
  logic [0:0] f1302_wen;
  logic [31:0] f1302_wdata;
  logic [0:0] f1302_clk;
  logic [0:0] f1302_rst;
  logic [31:0] f1302_rdata;
  sr_buffer_32_1 f1302(.wen(f1302_wen), .wdata(f1302_wdata), .clk(f1302_clk), .rst(f1302_rst), .rdata(f1302_rdata));
  assign f1302_clk = clk;
  assign f1302_rst = rst;
  // Bindings to f1302

  // f1304
  logic [0:0] f1304_wen;
  logic [31:0] f1304_wdata;
  logic [0:0] f1304_clk;
  logic [0:0] f1304_rst;
  logic [31:0] f1304_rdata;
  sr_buffer_32_1 f1304(.wen(f1304_wen), .wdata(f1304_wdata), .clk(f1304_clk), .rst(f1304_rst), .rdata(f1304_rdata));
  assign f1304_clk = clk;
  assign f1304_rst = rst;
  // Bindings to f1304

  // f1306
  logic [0:0] f1306_wen;
  logic [31:0] f1306_wdata;
  logic [0:0] f1306_clk;
  logic [0:0] f1306_rst;
  logic [31:0] f1306_rdata;
  sr_buffer_32_1 f1306(.wen(f1306_wen), .wdata(f1306_wdata), .clk(f1306_clk), .rst(f1306_rst), .rdata(f1306_rdata));
  assign f1306_clk = clk;
  assign f1306_rst = rst;
  // Bindings to f1306

  // f1308
  logic [0:0] f1308_wen;
  logic [31:0] f1308_wdata;
  logic [0:0] f1308_clk;
  logic [0:0] f1308_rst;
  logic [31:0] f1308_rdata;
  sr_buffer_32_1 f1308(.wen(f1308_wen), .wdata(f1308_wdata), .clk(f1308_clk), .rst(f1308_rst), .rdata(f1308_rdata));
  assign f1308_clk = clk;
  assign f1308_rst = rst;
  // Bindings to f1308

  // f1310
  logic [0:0] f1310_wen;
  logic [31:0] f1310_wdata;
  logic [0:0] f1310_clk;
  logic [0:0] f1310_rst;
  logic [31:0] f1310_rdata;
  sr_buffer_32_1 f1310(.wen(f1310_wen), .wdata(f1310_wdata), .clk(f1310_clk), .rst(f1310_rst), .rdata(f1310_rdata));
  assign f1310_clk = clk;
  assign f1310_rst = rst;
  // Bindings to f1310

  // f1312
  logic [0:0] f1312_wen;
  logic [31:0] f1312_wdata;
  logic [0:0] f1312_clk;
  logic [0:0] f1312_rst;
  logic [31:0] f1312_rdata;
  sr_buffer_32_1 f1312(.wen(f1312_wen), .wdata(f1312_wdata), .clk(f1312_clk), .rst(f1312_rst), .rdata(f1312_rdata));
  assign f1312_clk = clk;
  assign f1312_rst = rst;
  // Bindings to f1312

  // f1314
  logic [0:0] f1314_wen;
  logic [31:0] f1314_wdata;
  logic [0:0] f1314_clk;
  logic [0:0] f1314_rst;
  logic [31:0] f1314_rdata;
  sr_buffer_32_1 f1314(.wen(f1314_wen), .wdata(f1314_wdata), .clk(f1314_clk), .rst(f1314_rst), .rdata(f1314_rdata));
  assign f1314_clk = clk;
  assign f1314_rst = rst;
  // Bindings to f1314

  // f1316
  logic [0:0] f1316_wen;
  logic [31:0] f1316_wdata;
  logic [0:0] f1316_clk;
  logic [0:0] f1316_rst;
  logic [31:0] f1316_rdata;
  sr_buffer_32_1 f1316(.wen(f1316_wen), .wdata(f1316_wdata), .clk(f1316_clk), .rst(f1316_rst), .rdata(f1316_rdata));
  assign f1316_clk = clk;
  assign f1316_rst = rst;
  // Bindings to f1316

  // f1318
  logic [0:0] f1318_wen;
  logic [31:0] f1318_wdata;
  logic [0:0] f1318_clk;
  logic [0:0] f1318_rst;
  logic [31:0] f1318_rdata;
  sr_buffer_32_1 f1318(.wen(f1318_wen), .wdata(f1318_wdata), .clk(f1318_clk), .rst(f1318_rst), .rdata(f1318_rdata));
  assign f1318_clk = clk;
  assign f1318_rst = rst;
  // Bindings to f1318

  // f1320
  logic [0:0] f1320_wen;
  logic [31:0] f1320_wdata;
  logic [0:0] f1320_clk;
  logic [0:0] f1320_rst;
  logic [31:0] f1320_rdata;
  sr_buffer_32_1 f1320(.wen(f1320_wen), .wdata(f1320_wdata), .clk(f1320_clk), .rst(f1320_rst), .rdata(f1320_rdata));
  assign f1320_clk = clk;
  assign f1320_rst = rst;
  // Bindings to f1320

  // f1322
  logic [0:0] f1322_wen;
  logic [31:0] f1322_wdata;
  logic [0:0] f1322_clk;
  logic [0:0] f1322_rst;
  logic [31:0] f1322_rdata;
  sr_buffer_32_1 f1322(.wen(f1322_wen), .wdata(f1322_wdata), .clk(f1322_clk), .rst(f1322_rst), .rdata(f1322_rdata));
  assign f1322_clk = clk;
  assign f1322_rst = rst;
  // Bindings to f1322

  // f1324
  logic [0:0] f1324_wen;
  logic [31:0] f1324_wdata;
  logic [0:0] f1324_clk;
  logic [0:0] f1324_rst;
  logic [31:0] f1324_rdata;
  sr_buffer_32_1 f1324(.wen(f1324_wen), .wdata(f1324_wdata), .clk(f1324_clk), .rst(f1324_rst), .rdata(f1324_rdata));
  assign f1324_clk = clk;
  assign f1324_rst = rst;
  // Bindings to f1324

  // f1326
  logic [0:0] f1326_wen;
  logic [31:0] f1326_wdata;
  logic [0:0] f1326_clk;
  logic [0:0] f1326_rst;
  logic [31:0] f1326_rdata;
  sr_buffer_32_1 f1326(.wen(f1326_wen), .wdata(f1326_wdata), .clk(f1326_clk), .rst(f1326_rst), .rdata(f1326_rdata));
  assign f1326_clk = clk;
  assign f1326_rst = rst;
  // Bindings to f1326

  // f1328
  logic [0:0] f1328_wen;
  logic [31:0] f1328_wdata;
  logic [0:0] f1328_clk;
  logic [0:0] f1328_rst;
  logic [31:0] f1328_rdata;
  sr_buffer_32_1 f1328(.wen(f1328_wen), .wdata(f1328_wdata), .clk(f1328_clk), .rst(f1328_rst), .rdata(f1328_rdata));
  assign f1328_clk = clk;
  assign f1328_rst = rst;
  // Bindings to f1328

  // f1330
  logic [0:0] f1330_wen;
  logic [31:0] f1330_wdata;
  logic [0:0] f1330_clk;
  logic [0:0] f1330_rst;
  logic [31:0] f1330_rdata;
  sr_buffer_32_1 f1330(.wen(f1330_wen), .wdata(f1330_wdata), .clk(f1330_clk), .rst(f1330_rst), .rdata(f1330_rdata));
  assign f1330_clk = clk;
  assign f1330_rst = rst;
  // Bindings to f1330

  // f1332
  logic [0:0] f1332_wen;
  logic [31:0] f1332_wdata;
  logic [0:0] f1332_clk;
  logic [0:0] f1332_rst;
  logic [31:0] f1332_rdata;
  sr_buffer_32_1 f1332(.wen(f1332_wen), .wdata(f1332_wdata), .clk(f1332_clk), .rst(f1332_rst), .rdata(f1332_rdata));
  assign f1332_clk = clk;
  assign f1332_rst = rst;
  // Bindings to f1332

  // f1334
  logic [0:0] f1334_wen;
  logic [31:0] f1334_wdata;
  logic [0:0] f1334_clk;
  logic [0:0] f1334_rst;
  logic [31:0] f1334_rdata;
  sr_buffer_32_1 f1334(.wen(f1334_wen), .wdata(f1334_wdata), .clk(f1334_clk), .rst(f1334_rst), .rdata(f1334_rdata));
  assign f1334_clk = clk;
  assign f1334_rst = rst;
  // Bindings to f1334

  // f1336
  logic [0:0] f1336_wen;
  logic [31:0] f1336_wdata;
  logic [0:0] f1336_clk;
  logic [0:0] f1336_rst;
  logic [31:0] f1336_rdata;
  sr_buffer_32_1 f1336(.wen(f1336_wen), .wdata(f1336_wdata), .clk(f1336_clk), .rst(f1336_rst), .rdata(f1336_rdata));
  assign f1336_clk = clk;
  assign f1336_rst = rst;
  // Bindings to f1336

  // f1338
  logic [0:0] f1338_wen;
  logic [31:0] f1338_wdata;
  logic [0:0] f1338_clk;
  logic [0:0] f1338_rst;
  logic [31:0] f1338_rdata;
  sr_buffer_32_1 f1338(.wen(f1338_wen), .wdata(f1338_wdata), .clk(f1338_clk), .rst(f1338_rst), .rdata(f1338_rdata));
  assign f1338_clk = clk;
  assign f1338_rst = rst;
  // Bindings to f1338

  // f1340
  logic [0:0] f1340_wen;
  logic [31:0] f1340_wdata;
  logic [0:0] f1340_clk;
  logic [0:0] f1340_rst;
  logic [31:0] f1340_rdata;
  sr_buffer_32_1 f1340(.wen(f1340_wen), .wdata(f1340_wdata), .clk(f1340_clk), .rst(f1340_rst), .rdata(f1340_rdata));
  assign f1340_clk = clk;
  assign f1340_rst = rst;
  // Bindings to f1340

  // f1342
  logic [0:0] f1342_wen;
  logic [31:0] f1342_wdata;
  logic [0:0] f1342_clk;
  logic [0:0] f1342_rst;
  logic [31:0] f1342_rdata;
  sr_buffer_32_1 f1342(.wen(f1342_wen), .wdata(f1342_wdata), .clk(f1342_clk), .rst(f1342_rst), .rdata(f1342_rdata));
  assign f1342_clk = clk;
  assign f1342_rst = rst;
  // Bindings to f1342

  // f1344
  logic [0:0] f1344_wen;
  logic [31:0] f1344_wdata;
  logic [0:0] f1344_clk;
  logic [0:0] f1344_rst;
  logic [31:0] f1344_rdata;
  sr_buffer_32_1 f1344(.wen(f1344_wen), .wdata(f1344_wdata), .clk(f1344_clk), .rst(f1344_rst), .rdata(f1344_rdata));
  assign f1344_clk = clk;
  assign f1344_rst = rst;
  // Bindings to f1344

  // f1346
  logic [0:0] f1346_wen;
  logic [31:0] f1346_wdata;
  logic [0:0] f1346_clk;
  logic [0:0] f1346_rst;
  logic [31:0] f1346_rdata;
  sr_buffer_32_1 f1346(.wen(f1346_wen), .wdata(f1346_wdata), .clk(f1346_clk), .rst(f1346_rst), .rdata(f1346_rdata));
  assign f1346_clk = clk;
  assign f1346_rst = rst;
  // Bindings to f1346

  // f1348
  logic [0:0] f1348_wen;
  logic [31:0] f1348_wdata;
  logic [0:0] f1348_clk;
  logic [0:0] f1348_rst;
  logic [31:0] f1348_rdata;
  sr_buffer_32_1 f1348(.wen(f1348_wen), .wdata(f1348_wdata), .clk(f1348_clk), .rst(f1348_rst), .rdata(f1348_rdata));
  assign f1348_clk = clk;
  assign f1348_rst = rst;
  // Bindings to f1348

  // f1350
  logic [0:0] f1350_wen;
  logic [31:0] f1350_wdata;
  logic [0:0] f1350_clk;
  logic [0:0] f1350_rst;
  logic [31:0] f1350_rdata;
  sr_buffer_32_1 f1350(.wen(f1350_wen), .wdata(f1350_wdata), .clk(f1350_clk), .rst(f1350_rst), .rdata(f1350_rdata));
  assign f1350_clk = clk;
  assign f1350_rst = rst;
  // Bindings to f1350

  // f1352
  logic [0:0] f1352_wen;
  logic [31:0] f1352_wdata;
  logic [0:0] f1352_clk;
  logic [0:0] f1352_rst;
  logic [31:0] f1352_rdata;
  sr_buffer_32_1 f1352(.wen(f1352_wen), .wdata(f1352_wdata), .clk(f1352_clk), .rst(f1352_rst), .rdata(f1352_rdata));
  assign f1352_clk = clk;
  assign f1352_rst = rst;
  // Bindings to f1352

  // f1354
  logic [0:0] f1354_wen;
  logic [31:0] f1354_wdata;
  logic [0:0] f1354_clk;
  logic [0:0] f1354_rst;
  logic [31:0] f1354_rdata;
  sr_buffer_32_1 f1354(.wen(f1354_wen), .wdata(f1354_wdata), .clk(f1354_clk), .rst(f1354_rst), .rdata(f1354_rdata));
  assign f1354_clk = clk;
  assign f1354_rst = rst;
  // Bindings to f1354

  // f1356
  logic [0:0] f1356_wen;
  logic [31:0] f1356_wdata;
  logic [0:0] f1356_clk;
  logic [0:0] f1356_rst;
  logic [31:0] f1356_rdata;
  sr_buffer_32_1 f1356(.wen(f1356_wen), .wdata(f1356_wdata), .clk(f1356_clk), .rst(f1356_rst), .rdata(f1356_rdata));
  assign f1356_clk = clk;
  assign f1356_rst = rst;
  // Bindings to f1356

  // f1358
  logic [0:0] f1358_wen;
  logic [31:0] f1358_wdata;
  logic [0:0] f1358_clk;
  logic [0:0] f1358_rst;
  logic [31:0] f1358_rdata;
  sr_buffer_32_1 f1358(.wen(f1358_wen), .wdata(f1358_wdata), .clk(f1358_clk), .rst(f1358_rst), .rdata(f1358_rdata));
  assign f1358_clk = clk;
  assign f1358_rst = rst;
  // Bindings to f1358

  // f1360
  logic [0:0] f1360_wen;
  logic [31:0] f1360_wdata;
  logic [0:0] f1360_clk;
  logic [0:0] f1360_rst;
  logic [31:0] f1360_rdata;
  sr_buffer_32_1 f1360(.wen(f1360_wen), .wdata(f1360_wdata), .clk(f1360_clk), .rst(f1360_rst), .rdata(f1360_rdata));
  assign f1360_clk = clk;
  assign f1360_rst = rst;
  // Bindings to f1360

  // f1362
  logic [0:0] f1362_wen;
  logic [31:0] f1362_wdata;
  logic [0:0] f1362_clk;
  logic [0:0] f1362_rst;
  logic [31:0] f1362_rdata;
  sr_buffer_32_1 f1362(.wen(f1362_wen), .wdata(f1362_wdata), .clk(f1362_clk), .rst(f1362_rst), .rdata(f1362_rdata));
  assign f1362_clk = clk;
  assign f1362_rst = rst;
  // Bindings to f1362

  // f1364
  logic [0:0] f1364_wen;
  logic [31:0] f1364_wdata;
  logic [0:0] f1364_clk;
  logic [0:0] f1364_rst;
  logic [31:0] f1364_rdata;
  sr_buffer_32_1 f1364(.wen(f1364_wen), .wdata(f1364_wdata), .clk(f1364_clk), .rst(f1364_rst), .rdata(f1364_rdata));
  assign f1364_clk = clk;
  assign f1364_rst = rst;
  // Bindings to f1364

  // f1366
  logic [0:0] f1366_wen;
  logic [31:0] f1366_wdata;
  logic [0:0] f1366_clk;
  logic [0:0] f1366_rst;
  logic [31:0] f1366_rdata;
  sr_buffer_32_1 f1366(.wen(f1366_wen), .wdata(f1366_wdata), .clk(f1366_clk), .rst(f1366_rst), .rdata(f1366_rdata));
  assign f1366_clk = clk;
  assign f1366_rst = rst;
  // Bindings to f1366

  // f1368
  logic [0:0] f1368_wen;
  logic [31:0] f1368_wdata;
  logic [0:0] f1368_clk;
  logic [0:0] f1368_rst;
  logic [31:0] f1368_rdata;
  sr_buffer_32_1 f1368(.wen(f1368_wen), .wdata(f1368_wdata), .clk(f1368_clk), .rst(f1368_rst), .rdata(f1368_rdata));
  assign f1368_clk = clk;
  assign f1368_rst = rst;
  // Bindings to f1368

  // f1370
  logic [0:0] f1370_wen;
  logic [31:0] f1370_wdata;
  logic [0:0] f1370_clk;
  logic [0:0] f1370_rst;
  logic [31:0] f1370_rdata;
  sr_buffer_32_1 f1370(.wen(f1370_wen), .wdata(f1370_wdata), .clk(f1370_clk), .rst(f1370_rst), .rdata(f1370_rdata));
  assign f1370_clk = clk;
  assign f1370_rst = rst;
  // Bindings to f1370

  // f1372
  logic [0:0] f1372_wen;
  logic [31:0] f1372_wdata;
  logic [0:0] f1372_clk;
  logic [0:0] f1372_rst;
  logic [31:0] f1372_rdata;
  sr_buffer_32_1 f1372(.wen(f1372_wen), .wdata(f1372_wdata), .clk(f1372_clk), .rst(f1372_rst), .rdata(f1372_rdata));
  assign f1372_clk = clk;
  assign f1372_rst = rst;
  // Bindings to f1372

  // f1374
  logic [0:0] f1374_wen;
  logic [31:0] f1374_wdata;
  logic [0:0] f1374_clk;
  logic [0:0] f1374_rst;
  logic [31:0] f1374_rdata;
  sr_buffer_32_1 f1374(.wen(f1374_wen), .wdata(f1374_wdata), .clk(f1374_clk), .rst(f1374_rst), .rdata(f1374_rdata));
  assign f1374_clk = clk;
  assign f1374_rst = rst;
  // Bindings to f1374

  // f1376
  logic [0:0] f1376_wen;
  logic [31:0] f1376_wdata;
  logic [0:0] f1376_clk;
  logic [0:0] f1376_rst;
  logic [31:0] f1376_rdata;
  sr_buffer_32_1 f1376(.wen(f1376_wen), .wdata(f1376_wdata), .clk(f1376_clk), .rst(f1376_rst), .rdata(f1376_rdata));
  assign f1376_clk = clk;
  assign f1376_rst = rst;
  // Bindings to f1376

  // f1378
  logic [0:0] f1378_wen;
  logic [31:0] f1378_wdata;
  logic [0:0] f1378_clk;
  logic [0:0] f1378_rst;
  logic [31:0] f1378_rdata;
  sr_buffer_32_1 f1378(.wen(f1378_wen), .wdata(f1378_wdata), .clk(f1378_clk), .rst(f1378_rst), .rdata(f1378_rdata));
  assign f1378_clk = clk;
  assign f1378_rst = rst;
  // Bindings to f1378

  // f1380
  logic [0:0] f1380_wen;
  logic [31:0] f1380_wdata;
  logic [0:0] f1380_clk;
  logic [0:0] f1380_rst;
  logic [31:0] f1380_rdata;
  sr_buffer_32_1 f1380(.wen(f1380_wen), .wdata(f1380_wdata), .clk(f1380_clk), .rst(f1380_rst), .rdata(f1380_rdata));
  assign f1380_clk = clk;
  assign f1380_rst = rst;
  // Bindings to f1380

  // f1382
  logic [0:0] f1382_wen;
  logic [31:0] f1382_wdata;
  logic [0:0] f1382_clk;
  logic [0:0] f1382_rst;
  logic [31:0] f1382_rdata;
  sr_buffer_32_1 f1382(.wen(f1382_wen), .wdata(f1382_wdata), .clk(f1382_clk), .rst(f1382_rst), .rdata(f1382_rdata));
  assign f1382_clk = clk;
  assign f1382_rst = rst;
  // Bindings to f1382

  // f1384
  logic [0:0] f1384_wen;
  logic [31:0] f1384_wdata;
  logic [0:0] f1384_clk;
  logic [0:0] f1384_rst;
  logic [31:0] f1384_rdata;
  sr_buffer_32_1 f1384(.wen(f1384_wen), .wdata(f1384_wdata), .clk(f1384_clk), .rst(f1384_rst), .rdata(f1384_rdata));
  assign f1384_clk = clk;
  assign f1384_rst = rst;
  // Bindings to f1384

  // f1386
  logic [0:0] f1386_wen;
  logic [31:0] f1386_wdata;
  logic [0:0] f1386_clk;
  logic [0:0] f1386_rst;
  logic [31:0] f1386_rdata;
  sr_buffer_32_1 f1386(.wen(f1386_wen), .wdata(f1386_wdata), .clk(f1386_clk), .rst(f1386_rst), .rdata(f1386_rdata));
  assign f1386_clk = clk;
  assign f1386_rst = rst;
  // Bindings to f1386

  // f1388
  logic [0:0] f1388_wen;
  logic [31:0] f1388_wdata;
  logic [0:0] f1388_clk;
  logic [0:0] f1388_rst;
  logic [31:0] f1388_rdata;
  sr_buffer_32_1 f1388(.wen(f1388_wen), .wdata(f1388_wdata), .clk(f1388_clk), .rst(f1388_rst), .rdata(f1388_rdata));
  assign f1388_clk = clk;
  assign f1388_rst = rst;
  // Bindings to f1388

  // f1390
  logic [0:0] f1390_wen;
  logic [31:0] f1390_wdata;
  logic [0:0] f1390_clk;
  logic [0:0] f1390_rst;
  logic [31:0] f1390_rdata;
  sr_buffer_32_1 f1390(.wen(f1390_wen), .wdata(f1390_wdata), .clk(f1390_clk), .rst(f1390_rst), .rdata(f1390_rdata));
  assign f1390_clk = clk;
  assign f1390_rst = rst;
  // Bindings to f1390

  // f1392
  logic [0:0] f1392_wen;
  logic [31:0] f1392_wdata;
  logic [0:0] f1392_clk;
  logic [0:0] f1392_rst;
  logic [31:0] f1392_rdata;
  sr_buffer_32_1 f1392(.wen(f1392_wen), .wdata(f1392_wdata), .clk(f1392_clk), .rst(f1392_rst), .rdata(f1392_rdata));
  assign f1392_clk = clk;
  assign f1392_rst = rst;
  // Bindings to f1392

  // f1394
  logic [0:0] f1394_wen;
  logic [31:0] f1394_wdata;
  logic [0:0] f1394_clk;
  logic [0:0] f1394_rst;
  logic [31:0] f1394_rdata;
  sr_buffer_32_1 f1394(.wen(f1394_wen), .wdata(f1394_wdata), .clk(f1394_clk), .rst(f1394_rst), .rdata(f1394_rdata));
  assign f1394_clk = clk;
  assign f1394_rst = rst;
  // Bindings to f1394

  // f1396
  logic [0:0] f1396_wen;
  logic [31:0] f1396_wdata;
  logic [0:0] f1396_clk;
  logic [0:0] f1396_rst;
  logic [31:0] f1396_rdata;
  sr_buffer_32_1 f1396(.wen(f1396_wen), .wdata(f1396_wdata), .clk(f1396_clk), .rst(f1396_rst), .rdata(f1396_rdata));
  assign f1396_clk = clk;
  assign f1396_rst = rst;
  // Bindings to f1396

  // f1398
  logic [0:0] f1398_wen;
  logic [31:0] f1398_wdata;
  logic [0:0] f1398_clk;
  logic [0:0] f1398_rst;
  logic [31:0] f1398_rdata;
  sr_buffer_32_1 f1398(.wen(f1398_wen), .wdata(f1398_wdata), .clk(f1398_clk), .rst(f1398_rst), .rdata(f1398_rdata));
  assign f1398_clk = clk;
  assign f1398_rst = rst;
  // Bindings to f1398

  // f1400
  logic [0:0] f1400_wen;
  logic [31:0] f1400_wdata;
  logic [0:0] f1400_clk;
  logic [0:0] f1400_rst;
  logic [31:0] f1400_rdata;
  sr_buffer_32_1 f1400(.wen(f1400_wen), .wdata(f1400_wdata), .clk(f1400_clk), .rst(f1400_rst), .rdata(f1400_rdata));
  assign f1400_clk = clk;
  assign f1400_rst = rst;
  // Bindings to f1400

  // f1402
  logic [0:0] f1402_wen;
  logic [31:0] f1402_wdata;
  logic [0:0] f1402_clk;
  logic [0:0] f1402_rst;
  logic [31:0] f1402_rdata;
  sr_buffer_32_1 f1402(.wen(f1402_wen), .wdata(f1402_wdata), .clk(f1402_clk), .rst(f1402_rst), .rdata(f1402_rdata));
  assign f1402_clk = clk;
  assign f1402_rst = rst;
  // Bindings to f1402

  // f1404
  logic [0:0] f1404_wen;
  logic [31:0] f1404_wdata;
  logic [0:0] f1404_clk;
  logic [0:0] f1404_rst;
  logic [31:0] f1404_rdata;
  sr_buffer_32_1 f1404(.wen(f1404_wen), .wdata(f1404_wdata), .clk(f1404_clk), .rst(f1404_rst), .rdata(f1404_rdata));
  assign f1404_clk = clk;
  assign f1404_rst = rst;
  // Bindings to f1404

  // f1406
  logic [0:0] f1406_wen;
  logic [31:0] f1406_wdata;
  logic [0:0] f1406_clk;
  logic [0:0] f1406_rst;
  logic [31:0] f1406_rdata;
  sr_buffer_32_1 f1406(.wen(f1406_wen), .wdata(f1406_wdata), .clk(f1406_clk), .rst(f1406_rst), .rdata(f1406_rdata));
  assign f1406_clk = clk;
  assign f1406_rst = rst;
  // Bindings to f1406

  // f1408
  logic [0:0] f1408_wen;
  logic [31:0] f1408_wdata;
  logic [0:0] f1408_clk;
  logic [0:0] f1408_rst;
  logic [31:0] f1408_rdata;
  sr_buffer_32_1 f1408(.wen(f1408_wen), .wdata(f1408_wdata), .clk(f1408_clk), .rst(f1408_rst), .rdata(f1408_rdata));
  assign f1408_clk = clk;
  assign f1408_rst = rst;
  // Bindings to f1408

  // f1410
  logic [0:0] f1410_wen;
  logic [31:0] f1410_wdata;
  logic [0:0] f1410_clk;
  logic [0:0] f1410_rst;
  logic [31:0] f1410_rdata;
  sr_buffer_32_1 f1410(.wen(f1410_wen), .wdata(f1410_wdata), .clk(f1410_clk), .rst(f1410_rst), .rdata(f1410_rdata));
  assign f1410_clk = clk;
  assign f1410_rst = rst;
  // Bindings to f1410

  // f1412
  logic [0:0] f1412_wen;
  logic [31:0] f1412_wdata;
  logic [0:0] f1412_clk;
  logic [0:0] f1412_rst;
  logic [31:0] f1412_rdata;
  sr_buffer_32_1 f1412(.wen(f1412_wen), .wdata(f1412_wdata), .clk(f1412_clk), .rst(f1412_rst), .rdata(f1412_rdata));
  assign f1412_clk = clk;
  assign f1412_rst = rst;
  // Bindings to f1412

  // f1414
  logic [0:0] f1414_wen;
  logic [31:0] f1414_wdata;
  logic [0:0] f1414_clk;
  logic [0:0] f1414_rst;
  logic [31:0] f1414_rdata;
  sr_buffer_32_1 f1414(.wen(f1414_wen), .wdata(f1414_wdata), .clk(f1414_clk), .rst(f1414_rst), .rdata(f1414_rdata));
  assign f1414_clk = clk;
  assign f1414_rst = rst;
  // Bindings to f1414

  // f1416
  logic [0:0] f1416_wen;
  logic [31:0] f1416_wdata;
  logic [0:0] f1416_clk;
  logic [0:0] f1416_rst;
  logic [31:0] f1416_rdata;
  sr_buffer_32_1 f1416(.wen(f1416_wen), .wdata(f1416_wdata), .clk(f1416_clk), .rst(f1416_rst), .rdata(f1416_rdata));
  assign f1416_clk = clk;
  assign f1416_rst = rst;
  // Bindings to f1416

  // f1418
  logic [0:0] f1418_wen;
  logic [31:0] f1418_wdata;
  logic [0:0] f1418_clk;
  logic [0:0] f1418_rst;
  logic [31:0] f1418_rdata;
  sr_buffer_32_1 f1418(.wen(f1418_wen), .wdata(f1418_wdata), .clk(f1418_clk), .rst(f1418_rst), .rdata(f1418_rdata));
  assign f1418_clk = clk;
  assign f1418_rst = rst;
  // Bindings to f1418

  // f1420
  logic [0:0] f1420_wen;
  logic [31:0] f1420_wdata;
  logic [0:0] f1420_clk;
  logic [0:0] f1420_rst;
  logic [31:0] f1420_rdata;
  sr_buffer_32_1 f1420(.wen(f1420_wen), .wdata(f1420_wdata), .clk(f1420_clk), .rst(f1420_rst), .rdata(f1420_rdata));
  assign f1420_clk = clk;
  assign f1420_rst = rst;
  // Bindings to f1420

  // f1422
  logic [0:0] f1422_wen;
  logic [31:0] f1422_wdata;
  logic [0:0] f1422_clk;
  logic [0:0] f1422_rst;
  logic [31:0] f1422_rdata;
  sr_buffer_32_1 f1422(.wen(f1422_wen), .wdata(f1422_wdata), .clk(f1422_clk), .rst(f1422_rst), .rdata(f1422_rdata));
  assign f1422_clk = clk;
  assign f1422_rst = rst;
  // Bindings to f1422

  // f1424
  logic [0:0] f1424_wen;
  logic [31:0] f1424_wdata;
  logic [0:0] f1424_clk;
  logic [0:0] f1424_rst;
  logic [31:0] f1424_rdata;
  sr_buffer_32_1 f1424(.wen(f1424_wen), .wdata(f1424_wdata), .clk(f1424_clk), .rst(f1424_rst), .rdata(f1424_rdata));
  assign f1424_clk = clk;
  assign f1424_rst = rst;
  // Bindings to f1424

  // f1426
  logic [0:0] f1426_wen;
  logic [31:0] f1426_wdata;
  logic [0:0] f1426_clk;
  logic [0:0] f1426_rst;
  logic [31:0] f1426_rdata;
  sr_buffer_32_1 f1426(.wen(f1426_wen), .wdata(f1426_wdata), .clk(f1426_clk), .rst(f1426_rst), .rdata(f1426_rdata));
  assign f1426_clk = clk;
  assign f1426_rst = rst;
  // Bindings to f1426

  // f1428
  logic [0:0] f1428_wen;
  logic [31:0] f1428_wdata;
  logic [0:0] f1428_clk;
  logic [0:0] f1428_rst;
  logic [31:0] f1428_rdata;
  sr_buffer_32_1 f1428(.wen(f1428_wen), .wdata(f1428_wdata), .clk(f1428_clk), .rst(f1428_rst), .rdata(f1428_rdata));
  assign f1428_clk = clk;
  assign f1428_rst = rst;
  // Bindings to f1428

  // f1430
  logic [0:0] f1430_wen;
  logic [31:0] f1430_wdata;
  logic [0:0] f1430_clk;
  logic [0:0] f1430_rst;
  logic [31:0] f1430_rdata;
  sr_buffer_32_1 f1430(.wen(f1430_wen), .wdata(f1430_wdata), .clk(f1430_clk), .rst(f1430_rst), .rdata(f1430_rdata));
  assign f1430_clk = clk;
  assign f1430_rst = rst;
  // Bindings to f1430

  // f1432
  logic [0:0] f1432_wen;
  logic [31:0] f1432_wdata;
  logic [0:0] f1432_clk;
  logic [0:0] f1432_rst;
  logic [31:0] f1432_rdata;
  sr_buffer_32_1 f1432(.wen(f1432_wen), .wdata(f1432_wdata), .clk(f1432_clk), .rst(f1432_rst), .rdata(f1432_rdata));
  assign f1432_clk = clk;
  assign f1432_rst = rst;
  // Bindings to f1432

  // f1434
  logic [0:0] f1434_wen;
  logic [31:0] f1434_wdata;
  logic [0:0] f1434_clk;
  logic [0:0] f1434_rst;
  logic [31:0] f1434_rdata;
  sr_buffer_32_1 f1434(.wen(f1434_wen), .wdata(f1434_wdata), .clk(f1434_clk), .rst(f1434_rst), .rdata(f1434_rdata));
  assign f1434_clk = clk;
  assign f1434_rst = rst;
  // Bindings to f1434

  // f1436
  logic [0:0] f1436_wen;
  logic [31:0] f1436_wdata;
  logic [0:0] f1436_clk;
  logic [0:0] f1436_rst;
  logic [31:0] f1436_rdata;
  sr_buffer_32_1 f1436(.wen(f1436_wen), .wdata(f1436_wdata), .clk(f1436_clk), .rst(f1436_rst), .rdata(f1436_rdata));
  assign f1436_clk = clk;
  assign f1436_rst = rst;
  // Bindings to f1436

  // f1438
  logic [0:0] f1438_wen;
  logic [31:0] f1438_wdata;
  logic [0:0] f1438_clk;
  logic [0:0] f1438_rst;
  logic [31:0] f1438_rdata;
  sr_buffer_32_1 f1438(.wen(f1438_wen), .wdata(f1438_wdata), .clk(f1438_clk), .rst(f1438_rst), .rdata(f1438_rdata));
  assign f1438_clk = clk;
  assign f1438_rst = rst;
  // Bindings to f1438

  // f1440
  logic [0:0] f1440_wen;
  logic [31:0] f1440_wdata;
  logic [0:0] f1440_clk;
  logic [0:0] f1440_rst;
  logic [31:0] f1440_rdata;
  sr_buffer_32_1 f1440(.wen(f1440_wen), .wdata(f1440_wdata), .clk(f1440_clk), .rst(f1440_rst), .rdata(f1440_rdata));
  assign f1440_clk = clk;
  assign f1440_rst = rst;
  // Bindings to f1440

  // f1442
  logic [0:0] f1442_wen;
  logic [31:0] f1442_wdata;
  logic [0:0] f1442_clk;
  logic [0:0] f1442_rst;
  logic [31:0] f1442_rdata;
  sr_buffer_32_1 f1442(.wen(f1442_wen), .wdata(f1442_wdata), .clk(f1442_clk), .rst(f1442_rst), .rdata(f1442_rdata));
  assign f1442_clk = clk;
  assign f1442_rst = rst;
  // Bindings to f1442

  // f1444
  logic [0:0] f1444_wen;
  logic [31:0] f1444_wdata;
  logic [0:0] f1444_clk;
  logic [0:0] f1444_rst;
  logic [31:0] f1444_rdata;
  sr_buffer_32_1 f1444(.wen(f1444_wen), .wdata(f1444_wdata), .clk(f1444_clk), .rst(f1444_rst), .rdata(f1444_rdata));
  assign f1444_clk = clk;
  assign f1444_rst = rst;
  // Bindings to f1444

  // f1446
  logic [0:0] f1446_wen;
  logic [31:0] f1446_wdata;
  logic [0:0] f1446_clk;
  logic [0:0] f1446_rst;
  logic [31:0] f1446_rdata;
  sr_buffer_32_1 f1446(.wen(f1446_wen), .wdata(f1446_wdata), .clk(f1446_clk), .rst(f1446_rst), .rdata(f1446_rdata));
  assign f1446_clk = clk;
  assign f1446_rst = rst;
  // Bindings to f1446



endmodule


module dark_weights_normed_gauss_blur_1_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1265;
    end
  end

endmodule


module fused_level_0_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (-1249 + d0 == 0 && 1248 - d1 >= 0) ? (17695) : (1248 - d1 >= 0 && 1248 - d0 >= 0) ? (17696) : (-1249 + d1 == 0) ? ((17681 - d0)) : 0;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2527;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1264;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_1_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_update_0_write_wen(output [0:0] dark_weights_normed_update_0_write_wen);

endmodule


module dark_weights_normed_gauss_blur_1_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (1259 - d0 >= 0) ? (1263) : (-1260 + d0 == 0) ? (1263) : 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_update_0_write_wdata(output [31:0] dark_weights_normed_update_0_write_wdata);

endmodule


module in_wire_dark_weights_normed_gauss_blur_1_update_0_read_dummy(output [287:0] dark_weights_normed_gauss_blur_1_update_0_read_dummy);

endmodule


module out_wire_dark_weights_normed_gauss_blur_1_update_0_read_rdata(input [287:0] dark_weights_normed_gauss_blur_1_update_0_read_rdata);

endmodule


module dark_weights_normed(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] fused_level_0_update_0_read_rdata, output [287:0] dark_weights_normed_gauss_blur_1_update_0_read_rdata, input [287:0] dark_weights_normed_gauss_blur_1_update_0_read_dummy, input [31:0] dark_weights_normed_update_0_write_wdata, input [31:0] fused_level_0_update_0_read_dummy, input [0:0] dark_weights_normed_update_0_write_wen);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_4;
  logic [287:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_4_stage_1;
  reg [287:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_4_stage_1 <= rd_4;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to fused_level_0_update_0_read_rdata
    // wr_5
  assign fused_level_0_update_0_read_rdata = rd_4;

  // Bindings to dark_weights_normed_gauss_blur_1_update_0_read_rdata
    // wr_3
  assign dark_weights_normed_gauss_blur_1_update_0_read_rdata = rd_2;

  // Bindings to dark_weights_normed_gauss_blur_1_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_weights_normed_gauss_blur_1_update_0_read_dummy;

  // Bindings to dark_weights_normed_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_normed_update_0_write_wdata;

  // selector_dark_weights_normed_gauss_blur_1_rd6_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd6_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd6_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd6_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd6_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd6_select_out;
  dark_weights_normed_gauss_blur_1_rd6_select selector_dark_weights_normed_gauss_blur_1_rd6_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd6_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd6_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd6_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd6_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd6_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd6_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd6_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd6_select

  // selector_dark_weights_normed_gauss_blur_1_rd8_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd8_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd8_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd8_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd8_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd8_select_out;
  dark_weights_normed_gauss_blur_1_rd8_select selector_dark_weights_normed_gauss_blur_1_rd8_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd8_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd8_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd8_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd8_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd8_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd8_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd8_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd8_select

  // selector_dark_weights_normed_gauss_blur_1_rd7_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd7_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd7_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd7_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd7_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd7_select_out;
  dark_weights_normed_gauss_blur_1_rd7_select selector_dark_weights_normed_gauss_blur_1_rd7_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd7_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd7_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd7_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd7_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd7_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd7_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd7_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd7_select

  // selector_dark_weights_normed_gauss_blur_1_rd5_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd5_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd5_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd5_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd5_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd5_select_out;
  dark_weights_normed_gauss_blur_1_rd5_select selector_dark_weights_normed_gauss_blur_1_rd5_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd5_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd5_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd5_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd5_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd5_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd5_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd5_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd5_select

  // selector_dark_weights_normed_gauss_blur_1_rd3_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd3_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd3_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd3_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd3_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd3_select_out;
  dark_weights_normed_gauss_blur_1_rd3_select selector_dark_weights_normed_gauss_blur_1_rd3_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd3_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd3_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd3_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd3_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd3_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd3_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd3_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd3_select

  // selector_dark_weights_normed_gauss_blur_1_rd4_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd4_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd4_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd4_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd4_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd4_select_out;
  dark_weights_normed_gauss_blur_1_rd4_select selector_dark_weights_normed_gauss_blur_1_rd4_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd4_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd4_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd4_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd4_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd4_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd4_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd4_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd4_select

  // selector_dark_weights_normed_gauss_blur_1_rd2_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd2_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd2_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd2_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd2_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd2_select_out;
  dark_weights_normed_gauss_blur_1_rd2_select selector_dark_weights_normed_gauss_blur_1_rd2_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd2_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd2_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd2_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd2_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd2_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd2_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd2_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd2_select

  // Bindings to fused_level_0_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_0_update_0_read_dummy;

  // Bindings to dark_weights_normed_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_normed_update_0_write_wen;

  // selector_dark_weights_normed_gauss_blur_1_rd0_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd0_select_out;
  dark_weights_normed_gauss_blur_1_rd0_select selector_dark_weights_normed_gauss_blur_1_rd0_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd0_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd0_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd0_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd0_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd0_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd0_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd0_select

  // selector_fused_level_0_rd0_select
  logic [0:0] selector_fused_level_0_rd0_select_clk;
  logic [0:0] selector_fused_level_0_rd0_select_rst;
  logic [31:0] selector_fused_level_0_rd0_select_d0;
  logic [31:0] selector_fused_level_0_rd0_select_d1;
  logic [31:0] selector_fused_level_0_rd0_select_out;
  fused_level_0_rd0_select selector_fused_level_0_rd0_select(.clk(selector_fused_level_0_rd0_select_clk), .rst(selector_fused_level_0_rd0_select_rst), .d0(selector_fused_level_0_rd0_select_d0), .d1(selector_fused_level_0_rd0_select_d1), .out(selector_fused_level_0_rd0_select_out));
  assign selector_fused_level_0_rd0_select_clk = clk;
  assign selector_fused_level_0_rd0_select_rst = rst;
  // Bindings to selector_fused_level_0_rd0_select

  // dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_clk;
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_rst;
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_start;
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_done;
  dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0 dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0(.clk(dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_clk), .rst(dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_rst), .start(dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_start), .done(dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_done));
  assign dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_clk = clk;
  assign dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0_rst = rst;
  // Bindings to dark_weights_normed_dark_weights_normed_update_0_write0_to_fused_level_0_rd0

  // selector_dark_weights_normed_gauss_blur_1_rd1_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd1_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_1_rd1_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd1_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd1_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_1_rd1_select_out;
  dark_weights_normed_gauss_blur_1_rd1_select selector_dark_weights_normed_gauss_blur_1_rd1_select(.clk(selector_dark_weights_normed_gauss_blur_1_rd1_select_clk), .rst(selector_dark_weights_normed_gauss_blur_1_rd1_select_rst), .d0(selector_dark_weights_normed_gauss_blur_1_rd1_select_d0), .d1(selector_dark_weights_normed_gauss_blur_1_rd1_select_d1), .out(selector_dark_weights_normed_gauss_blur_1_rd1_select_out));
  assign selector_dark_weights_normed_gauss_blur_1_rd1_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_1_rd1_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_1_rd1_select

  // dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_clk;
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_rst;
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_start;
  logic [0:0] dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_done;
  dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9 dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9(.clk(dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_clk), .rst(dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_rst), .start(dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_start), .done(dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_done));
  assign dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_clk = clk;
  assign dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9_rst = rst;
  // Bindings to dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9



endmodule


module dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module dark_weights_normed_gauss_ds_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_gauss_blur_1_update_0_write_wen(output [0:0] dark_weights_normed_gauss_blur_1_update_0_write_wen);

endmodule


module in_wire_dark_weights_normed_gauss_blur_1_update_0_write_wdata(output [31:0] dark_weights_normed_gauss_blur_1_update_0_write_wdata);

endmodule


module in_wire_dark_weights_normed_gauss_ds_1_update_0_read_dummy(output [31:0] dark_weights_normed_gauss_ds_1_update_0_read_dummy);

endmodule


module out_wire_dark_weights_normed_gauss_ds_1_update_0_read_rdata(input [31:0] dark_weights_normed_gauss_ds_1_update_0_read_rdata);

endmodule


module in_wire_dark_weights_normed_gauss_ds_2_update_0_write_wen(output [0:0] dark_weights_normed_gauss_ds_2_update_0_write_wen);

endmodule


module fused_level_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 632;
    end
  end

endmodule


module in_wire_dark_weights_normed_gauss_ds_2_update_0_write_wdata(output [31:0] dark_weights_normed_gauss_ds_2_update_0_write_wdata);

endmodule


module in_wire_dark_weights_normed_gauss_blur_3_update_0_read_dummy(output [287:0] dark_weights_normed_gauss_blur_3_update_0_read_dummy);

endmodule


module out_wire_dark_weights_normed_gauss_blur_3_update_0_read_rdata(input [287:0] dark_weights_normed_gauss_blur_3_update_0_read_rdata);

endmodule


module final_merged_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] final_merged_2_update_0_write_wen, input [31:0] final_merged_2_update_0_write_wdata, input [31:0] final_merged_1_update_0_read_dummy, output [31:0] final_merged_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to final_merged_2_update_0_write_wen
    // rd_0
  assign rd_0 = final_merged_2_update_0_write_wen;

  // final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0
  logic [0:0] final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_clk;
  logic [0:0] final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_rst;
  logic [0:0] final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_start;
  logic [0:0] final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_done;
  final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0 final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0(.clk(final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_clk), .rst(final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_rst), .start(final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_start), .done(final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_done));
  assign final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_clk = clk;
  assign final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0_rst = rst;
  // Bindings to final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0

  // Bindings to final_merged_2_update_0_write_wdata
    // rd_1
  assign rd_1 = final_merged_2_update_0_write_wdata;

  // selector_final_merged_1_rd0_select
  logic [0:0] selector_final_merged_1_rd0_select_clk;
  logic [0:0] selector_final_merged_1_rd0_select_rst;
  logic [31:0] selector_final_merged_1_rd0_select_d0;
  logic [31:0] selector_final_merged_1_rd0_select_d1;
  logic [31:0] selector_final_merged_1_rd0_select_out;
  final_merged_1_rd0_select selector_final_merged_1_rd0_select(.clk(selector_final_merged_1_rd0_select_clk), .rst(selector_final_merged_1_rd0_select_rst), .d0(selector_final_merged_1_rd0_select_d0), .d1(selector_final_merged_1_rd0_select_d1), .out(selector_final_merged_1_rd0_select_out));
  assign selector_final_merged_1_rd0_select_clk = clk;
  assign selector_final_merged_1_rd0_select_rst = rst;
  // Bindings to selector_final_merged_1_rd0_select

  // Bindings to final_merged_1_update_0_read_dummy
    // rd_2
  assign rd_2 = final_merged_1_update_0_read_dummy;

  // Bindings to final_merged_1_update_0_read_rdata
    // wr_3
  assign final_merged_1_update_0_read_rdata = rd_2;



endmodule


module fused_level_0_fused_level_0_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module fused_level_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] fused_level_0_update_0_write_wen, input [31:0] fused_level_0_update_0_write_wdata, input [31:0] final_merged_0_update_0_read_dummy, output [31:0] final_merged_0_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // fused_level_0_fused_level_0_update_0_write0_merged_banks_1
  logic [0:0] fused_level_0_fused_level_0_update_0_write0_merged_banks_1_clk;
  logic [0:0] fused_level_0_fused_level_0_update_0_write0_merged_banks_1_rst;
  logic [0:0] fused_level_0_fused_level_0_update_0_write0_merged_banks_1_start;
  logic [0:0] fused_level_0_fused_level_0_update_0_write0_merged_banks_1_done;
  fused_level_0_fused_level_0_update_0_write0_merged_banks_1 fused_level_0_fused_level_0_update_0_write0_merged_banks_1(.clk(fused_level_0_fused_level_0_update_0_write0_merged_banks_1_clk), .rst(fused_level_0_fused_level_0_update_0_write0_merged_banks_1_rst), .start(fused_level_0_fused_level_0_update_0_write0_merged_banks_1_start), .done(fused_level_0_fused_level_0_update_0_write0_merged_banks_1_done));
  assign fused_level_0_fused_level_0_update_0_write0_merged_banks_1_clk = clk;
  assign fused_level_0_fused_level_0_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to fused_level_0_fused_level_0_update_0_write0_merged_banks_1

  // Bindings to fused_level_0_update_0_write_wen
    // rd_0
  assign rd_0 = fused_level_0_update_0_write_wen;

  // selector_final_merged_0_rd0_select
  logic [0:0] selector_final_merged_0_rd0_select_clk;
  logic [0:0] selector_final_merged_0_rd0_select_rst;
  logic [31:0] selector_final_merged_0_rd0_select_d0;
  logic [31:0] selector_final_merged_0_rd0_select_d1;
  logic [31:0] selector_final_merged_0_rd0_select_out;
  final_merged_0_rd0_select selector_final_merged_0_rd0_select(.clk(selector_final_merged_0_rd0_select_clk), .rst(selector_final_merged_0_rd0_select_rst), .d0(selector_final_merged_0_rd0_select_d0), .d1(selector_final_merged_0_rd0_select_d1), .out(selector_final_merged_0_rd0_select_out));
  assign selector_final_merged_0_rd0_select_clk = clk;
  assign selector_final_merged_0_rd0_select_rst = rst;
  // Bindings to selector_final_merged_0_rd0_select

  // Bindings to fused_level_0_update_0_write_wdata
    // rd_1
  assign rd_1 = fused_level_0_update_0_write_wdata;

  // Bindings to final_merged_0_update_0_read_dummy
    // rd_2
  assign rd_2 = final_merged_0_update_0_read_dummy;

  // Bindings to final_merged_0_update_0_read_rdata
    // wr_3
  assign final_merged_0_update_0_read_rdata = rd_2;



endmodule


module fused_level_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] fused_level_1_update_0_write_wen, input [31:0] fused_level_1_update_0_write_wdata, input [31:0] final_merged_1_update_0_read_dummy, output [31:0] final_merged_1_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // fused_level_1_fused_level_1_update_0_write0_merged_banks_1
  logic [0:0] fused_level_1_fused_level_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] fused_level_1_fused_level_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] fused_level_1_fused_level_1_update_0_write0_merged_banks_1_start;
  logic [0:0] fused_level_1_fused_level_1_update_0_write0_merged_banks_1_done;
  fused_level_1_fused_level_1_update_0_write0_merged_banks_1 fused_level_1_fused_level_1_update_0_write0_merged_banks_1(.clk(fused_level_1_fused_level_1_update_0_write0_merged_banks_1_clk), .rst(fused_level_1_fused_level_1_update_0_write0_merged_banks_1_rst), .start(fused_level_1_fused_level_1_update_0_write0_merged_banks_1_start), .done(fused_level_1_fused_level_1_update_0_write0_merged_banks_1_done));
  assign fused_level_1_fused_level_1_update_0_write0_merged_banks_1_clk = clk;
  assign fused_level_1_fused_level_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to fused_level_1_fused_level_1_update_0_write0_merged_banks_1

  // selector_final_merged_1_rd0_select
  logic [0:0] selector_final_merged_1_rd0_select_clk;
  logic [0:0] selector_final_merged_1_rd0_select_rst;
  logic [31:0] selector_final_merged_1_rd0_select_d0;
  logic [31:0] selector_final_merged_1_rd0_select_d1;
  logic [31:0] selector_final_merged_1_rd0_select_out;
  final_merged_1_rd0_select selector_final_merged_1_rd0_select(.clk(selector_final_merged_1_rd0_select_clk), .rst(selector_final_merged_1_rd0_select_rst), .d0(selector_final_merged_1_rd0_select_d0), .d1(selector_final_merged_1_rd0_select_d1), .out(selector_final_merged_1_rd0_select_out));
  assign selector_final_merged_1_rd0_select_clk = clk;
  assign selector_final_merged_1_rd0_select_rst = rst;
  // Bindings to selector_final_merged_1_rd0_select

  // Bindings to fused_level_1_update_0_write_wen
    // rd_0
  assign rd_0 = fused_level_1_update_0_write_wen;

  // Bindings to fused_level_1_update_0_write_wdata
    // rd_1
  assign rd_1 = fused_level_1_update_0_write_wdata;

  // Bindings to final_merged_1_update_0_read_dummy
    // rd_2
  assign rd_2 = final_merged_1_update_0_read_dummy;

  // Bindings to final_merged_1_update_0_read_rdata
    // wr_3
  assign final_merged_1_update_0_read_rdata = rd_2;



endmodule


module fused_level_2_fused_level_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module fused_level_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] fused_level_2_update_0_write_wdata, input [0:0] fused_level_2_update_0_write_wen, input [31:0] final_merged_2_update_0_read_dummy, output [31:0] final_merged_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // fused_level_2_fused_level_2_update_0_write0_merged_banks_1
  logic [0:0] fused_level_2_fused_level_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] fused_level_2_fused_level_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] fused_level_2_fused_level_2_update_0_write0_merged_banks_1_start;
  logic [0:0] fused_level_2_fused_level_2_update_0_write0_merged_banks_1_done;
  fused_level_2_fused_level_2_update_0_write0_merged_banks_1 fused_level_2_fused_level_2_update_0_write0_merged_banks_1(.clk(fused_level_2_fused_level_2_update_0_write0_merged_banks_1_clk), .rst(fused_level_2_fused_level_2_update_0_write0_merged_banks_1_rst), .start(fused_level_2_fused_level_2_update_0_write0_merged_banks_1_start), .done(fused_level_2_fused_level_2_update_0_write0_merged_banks_1_done));
  assign fused_level_2_fused_level_2_update_0_write0_merged_banks_1_clk = clk;
  assign fused_level_2_fused_level_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to fused_level_2_fused_level_2_update_0_write0_merged_banks_1

  // selector_final_merged_2_rd0_select
  logic [0:0] selector_final_merged_2_rd0_select_clk;
  logic [0:0] selector_final_merged_2_rd0_select_rst;
  logic [31:0] selector_final_merged_2_rd0_select_d0;
  logic [31:0] selector_final_merged_2_rd0_select_d1;
  logic [31:0] selector_final_merged_2_rd0_select_out;
  final_merged_2_rd0_select selector_final_merged_2_rd0_select(.clk(selector_final_merged_2_rd0_select_clk), .rst(selector_final_merged_2_rd0_select_rst), .d0(selector_final_merged_2_rd0_select_d0), .d1(selector_final_merged_2_rd0_select_d1), .out(selector_final_merged_2_rd0_select_out));
  assign selector_final_merged_2_rd0_select_clk = clk;
  assign selector_final_merged_2_rd0_select_rst = rst;
  // Bindings to selector_final_merged_2_rd0_select

  // Bindings to fused_level_2_update_0_write_wdata
    // rd_1
  assign rd_1 = fused_level_2_update_0_write_wdata;

  // Bindings to fused_level_2_update_0_write_wen
    // rd_0
  assign rd_0 = fused_level_2_update_0_write_wen;

  // Bindings to final_merged_2_update_0_read_dummy
    // rd_2
  assign rd_2 = final_merged_2_update_0_read_dummy;

  // Bindings to final_merged_2_update_0_read_rdata
    // wr_3
  assign final_merged_2_update_0_read_rdata = rd_2;



endmodule


module fused_level_1_fused_level_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module bright_gauss_ds_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module dark_laplace_us_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module dark_laplace_us_0_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_weights_normed_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_weights_normed_gauss_blur_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_gauss_blur_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_weights_normed_gauss_ds_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_weights_normed_gauss_ds_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_laplace_us_0_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_laplace_diff_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_laplace_diff_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_weights_normed_gauss_blur_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_gauss_ds_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_laplace_diff_0_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_weights_normed_gauss_blur_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_gauss_blur_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] bright_gauss_ds_2_update_0_read_rdata, input [31:0] bright_gauss_blur_2_update_0_write_wdata, input [31:0] bright_gauss_ds_2_update_0_read_dummy, input [0:0] bright_gauss_blur_2_update_0_write_wen);

  logic [31:0] rd_2;
  logic [0:0] rd_0;
  logic [31:0] rd_1;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_2_stage_1;
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_2_stage_1 <= rd_2;
      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;


    end

  end


  // Data processing units...
  // Bindings to bright_gauss_ds_2_update_0_read_rdata
    // wr_3
  assign bright_gauss_ds_2_update_0_read_rdata = rd_2;

  // Bindings to bright_gauss_blur_2_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_gauss_blur_2_update_0_write_wdata;

  // Bindings to bright_gauss_ds_2_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_gauss_ds_2_update_0_read_dummy;

  // selector_bright_gauss_ds_2_rd0_select
  logic [0:0] selector_bright_gauss_ds_2_rd0_select_clk;
  logic [0:0] selector_bright_gauss_ds_2_rd0_select_rst;
  logic [31:0] selector_bright_gauss_ds_2_rd0_select_d0;
  logic [31:0] selector_bright_gauss_ds_2_rd0_select_d1;
  logic [31:0] selector_bright_gauss_ds_2_rd0_select_out;
  bright_gauss_ds_2_rd0_select selector_bright_gauss_ds_2_rd0_select(.clk(selector_bright_gauss_ds_2_rd0_select_clk), .rst(selector_bright_gauss_ds_2_rd0_select_rst), .d0(selector_bright_gauss_ds_2_rd0_select_d0), .d1(selector_bright_gauss_ds_2_rd0_select_d1), .out(selector_bright_gauss_ds_2_rd0_select_out));
  assign selector_bright_gauss_ds_2_rd0_select_clk = clk;
  assign selector_bright_gauss_ds_2_rd0_select_rst = rst;
  // Bindings to selector_bright_gauss_ds_2_rd0_select

  // bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1
  logic [0:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_done;
  bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1 bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1(.clk(bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_clk), .rst(bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_rst), .start(bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_start), .done(bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_done));
  assign bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_clk = clk;
  assign bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1

  // Bindings to bright_gauss_blur_2_update_0_write_wen
    // rd_0
  assign rd_0 = bright_gauss_blur_2_update_0_write_wen;



endmodule


module sr_buffer_32_1(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 1;

  reg [31:0] data [0:0];

  reg [31:0] rdata_d;

  reg [0:0] waddr;

  wire [0:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module bright_bright_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_1260 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_1260 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10



endmodule


module bright_gauss_ds_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module sr_buffer_32_16431(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 16431;

  reg [31:0] data [16430:0];

  reg [31:0] rdata_d;

  reg [14:0] waddr;

  wire [14:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module sr_buffer_32_1260(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 1260;

  reg [31:0] data [1259:0];

  reg [31:0] rdata_d;

  reg [10:0] waddr;

  wire [10:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module in_wire_bright_gauss_blur_3_update_0_write_wen(output [0:0] bright_gauss_blur_3_update_0_write_wen);

endmodule


module bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_gauss_blur_3_update_0_write_wdata(output [31:0] bright_gauss_blur_3_update_0_write_wdata);

endmodule


module in_wire_bright_gauss_ds_3_update_0_read_dummy(output [31:0] bright_gauss_ds_3_update_0_read_dummy);

endmodule


module out_wire_bright_gauss_ds_3_update_0_read_rdata(input [31:0] bright_gauss_ds_3_update_0_read_rdata);

endmodule


module bright_gauss_blur_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] bright_gauss_ds_3_update_0_read_dummy, output [31:0] bright_gauss_ds_3_update_0_read_rdata, input [31:0] bright_gauss_blur_3_update_0_write_wdata, input [0:0] bright_gauss_blur_3_update_0_write_wen);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to bright_gauss_ds_3_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_gauss_ds_3_update_0_read_dummy;

  // bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1
  logic [0:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_done;
  bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1 bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1(.clk(bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_clk), .rst(bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_rst), .start(bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_start), .done(bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_done));
  assign bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_clk = clk;
  assign bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_gauss_blur_3_bright_gauss_blur_3_update_0_write0_merged_banks_1

  // Bindings to bright_gauss_ds_3_update_0_read_rdata
    // wr_3
  assign bright_gauss_ds_3_update_0_read_rdata = rd_2;

  // Bindings to bright_gauss_blur_3_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_gauss_blur_3_update_0_write_wdata;

  // selector_bright_gauss_ds_3_rd0_select
  logic [0:0] selector_bright_gauss_ds_3_rd0_select_clk;
  logic [0:0] selector_bright_gauss_ds_3_rd0_select_rst;
  logic [31:0] selector_bright_gauss_ds_3_rd0_select_d0;
  logic [31:0] selector_bright_gauss_ds_3_rd0_select_d1;
  logic [31:0] selector_bright_gauss_ds_3_rd0_select_out;
  bright_gauss_ds_3_rd0_select selector_bright_gauss_ds_3_rd0_select(.clk(selector_bright_gauss_ds_3_rd0_select_clk), .rst(selector_bright_gauss_ds_3_rd0_select_rst), .d0(selector_bright_gauss_ds_3_rd0_select_d0), .d1(selector_bright_gauss_ds_3_rd0_select_d1), .out(selector_bright_gauss_ds_3_rd0_select_out));
  assign selector_bright_gauss_ds_3_rd0_select_clk = clk;
  assign selector_bright_gauss_ds_3_rd0_select_rst = rst;
  // Bindings to selector_bright_gauss_ds_3_rd0_select

  // Bindings to bright_gauss_blur_3_update_0_write_wen
    // rd_0
  assign rd_0 = bright_gauss_blur_3_update_0_write_wen;



endmodule


module in_wire_bright_gauss_ds_3_update_0_write_wdata(output [31:0] bright_gauss_ds_3_update_0_write_wdata);

endmodule


module in_wire_bright_laplace_us_2_update_0_read_dummy(output [31:0] bright_laplace_us_2_update_0_read_dummy);

endmodule


module out_wire_bright_laplace_us_2_update_0_read_rdata(input [31:0] bright_laplace_us_2_update_0_read_rdata);

endmodule


module bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_628 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_628 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f17
  logic [0:0] f17_wen;
  logic [31:0] f17_wdata;
  logic [0:0] f17_clk;
  logic [0:0] f17_rst;
  logic [31:0] f17_rdata;
  sr_buffer_32_2527 f17(.wen(f17_wen), .wdata(f17_wdata), .clk(f17_clk), .rst(f17_rst), .rdata(f17_rdata));
  assign f17_clk = clk;
  assign f17_rst = rst;
  // Bindings to f17

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18



endmodule


module sr_buffer_32_628(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 628;

  reg [31:0] data [627:0];

  reg [31:0] rdata_d;

  reg [9:0] waddr;

  wire [9:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module sr_buffer_32_2527(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 2527;

  reg [31:0] data [2526:0];

  reg [31:0] rdata_d;

  reg [11:0] waddr;

  wire [11:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module sr_buffer_32_3790(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 3790;

  reg [31:0] data [3789:0];

  reg [31:0] rdata_d;

  reg [11:0] waddr;

  wire [11:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module in_wire_fused_level_3_update_0_read_dummy(output [31:0] fused_level_3_update_0_read_dummy);

endmodule


module out_wire_fused_level_3_update_0_read_rdata(input [31:0] fused_level_3_update_0_read_rdata);

endmodule


module bright_weights_normed_gauss_blur_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_weights_normed_gauss_blur_2_update_0_write_wen, input [31:0] bright_weights_normed_gauss_ds_2_update_0_read_dummy, input [31:0] bright_weights_normed_gauss_blur_2_update_0_write_wdata, output [31:0] bright_weights_normed_gauss_ds_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to bright_weights_normed_gauss_blur_2_update_0_write_wen
    // rd_0
  assign rd_0 = bright_weights_normed_gauss_blur_2_update_0_write_wen;

  // Bindings to bright_weights_normed_gauss_ds_2_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_gauss_ds_2_update_0_read_dummy;

  // selector_bright_weights_normed_gauss_ds_2_rd0_select
  logic [0:0] selector_bright_weights_normed_gauss_ds_2_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_gauss_ds_2_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_gauss_ds_2_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_gauss_ds_2_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_gauss_ds_2_rd0_select_out;
  bright_weights_normed_gauss_ds_2_rd0_select selector_bright_weights_normed_gauss_ds_2_rd0_select(.clk(selector_bright_weights_normed_gauss_ds_2_rd0_select_clk), .rst(selector_bright_weights_normed_gauss_ds_2_rd0_select_rst), .d0(selector_bright_weights_normed_gauss_ds_2_rd0_select_d0), .d1(selector_bright_weights_normed_gauss_ds_2_rd0_select_d1), .out(selector_bright_weights_normed_gauss_ds_2_rd0_select_out));
  assign selector_bright_weights_normed_gauss_ds_2_rd0_select_clk = clk;
  assign selector_bright_weights_normed_gauss_ds_2_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_gauss_ds_2_rd0_select

  // bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1
  logic [0:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_done;
  bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1 bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1(.clk(bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_clk), .rst(bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_rst), .start(bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_start), .done(bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_done));
  assign bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_clk = clk;
  assign bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1

  // Bindings to bright_weights_normed_gauss_blur_2_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_weights_normed_gauss_blur_2_update_0_write_wdata;

  // Bindings to bright_weights_normed_gauss_ds_2_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_gauss_ds_2_update_0_read_rdata = rd_2;



endmodule


module in_wire_bright_weights_normed_gauss_blur_3_update_0_write_wen(output [0:0] bright_weights_normed_gauss_blur_3_update_0_write_wen);

endmodule


module bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_weights_normed_gauss_blur_3_update_0_write_wdata(output [31:0] bright_weights_normed_gauss_blur_3_update_0_write_wdata);

endmodule


module bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_weights_normed_gauss_ds_3_update_0_read_dummy(output [31:0] bright_weights_normed_gauss_ds_3_update_0_read_dummy);

endmodule


module bright_weights_normed_gauss_ds_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module out_wire_bright_weights_normed_gauss_ds_3_update_0_read_rdata(input [31:0] bright_weights_normed_gauss_ds_3_update_0_read_rdata);

endmodule


module in_wire_bright_weights_normed_gauss_ds_3_update_0_write_wen(output [0:0] bright_weights_normed_gauss_ds_3_update_0_write_wen);

endmodule


module in_wire_dark_gauss_blur_2_update_0_write_wen(output [0:0] dark_gauss_blur_2_update_0_write_wen);

endmodule


module in_wire_dark_gauss_blur_2_update_0_write_wdata(output [31:0] dark_gauss_blur_2_update_0_write_wdata);

endmodule


module dark_gauss_ds_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_gauss_ds_2_update_0_read_dummy(output [31:0] dark_gauss_ds_2_update_0_read_dummy);

endmodule


module out_wire_dark_gauss_ds_2_update_0_read_rdata(input [31:0] dark_gauss_ds_2_update_0_read_rdata);

endmodule


module dark_gauss_blur_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_gauss_blur_2_update_0_write_wen, input [31:0] dark_gauss_ds_2_update_0_read_dummy, output [31:0] dark_gauss_ds_2_update_0_read_rdata, input [31:0] dark_gauss_blur_2_update_0_write_wdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_gauss_blur_2_update_0_write_wen
    // rd_0
  assign rd_0 = dark_gauss_blur_2_update_0_write_wen;

  // Bindings to dark_gauss_ds_2_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_gauss_ds_2_update_0_read_dummy;

  // selector_dark_gauss_ds_2_rd0_select
  logic [0:0] selector_dark_gauss_ds_2_rd0_select_clk;
  logic [0:0] selector_dark_gauss_ds_2_rd0_select_rst;
  logic [31:0] selector_dark_gauss_ds_2_rd0_select_d0;
  logic [31:0] selector_dark_gauss_ds_2_rd0_select_d1;
  logic [31:0] selector_dark_gauss_ds_2_rd0_select_out;
  dark_gauss_ds_2_rd0_select selector_dark_gauss_ds_2_rd0_select(.clk(selector_dark_gauss_ds_2_rd0_select_clk), .rst(selector_dark_gauss_ds_2_rd0_select_rst), .d0(selector_dark_gauss_ds_2_rd0_select_d0), .d1(selector_dark_gauss_ds_2_rd0_select_d1), .out(selector_dark_gauss_ds_2_rd0_select_out));
  assign selector_dark_gauss_ds_2_rd0_select_clk = clk;
  assign selector_dark_gauss_ds_2_rd0_select_rst = rst;
  // Bindings to selector_dark_gauss_ds_2_rd0_select

  // dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1
  logic [0:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_done;
  dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1 dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1(.clk(dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_clk), .rst(dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_rst), .start(dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_start), .done(dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_done));
  assign dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_clk = clk;
  assign dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_gauss_blur_2_dark_gauss_blur_2_update_0_write0_merged_banks_1

  // Bindings to dark_gauss_ds_2_update_0_read_rdata
    // wr_3
  assign dark_gauss_ds_2_update_0_read_rdata = rd_2;

  // Bindings to dark_gauss_blur_2_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_gauss_blur_2_update_0_write_wdata;



endmodule


module in_wire_dark_gauss_blur_3_update_0_write_wen(output [0:0] dark_gauss_blur_3_update_0_write_wen);

endmodule


module dark_gauss_ds_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_gauss_blur_3_update_0_write_wdata(output [31:0] dark_gauss_blur_3_update_0_write_wdata);

endmodule


module in_wire_dark_gauss_ds_3_update_0_read_dummy(output [31:0] dark_gauss_ds_3_update_0_read_dummy);

endmodule


module out_wire_dark_gauss_ds_3_update_0_read_rdata(input [31:0] dark_gauss_ds_3_update_0_read_rdata);

endmodule


module dark_gauss_blur_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] dark_gauss_ds_3_update_0_read_rdata, input [31:0] dark_gauss_blur_3_update_0_write_wdata, input [0:0] dark_gauss_blur_3_update_0_write_wen, input [31:0] dark_gauss_ds_3_update_0_read_dummy);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_gauss_ds_3_update_0_read_rdata
    // wr_3
  assign dark_gauss_ds_3_update_0_read_rdata = rd_2;

  // Bindings to dark_gauss_blur_3_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_gauss_blur_3_update_0_write_wdata;

  // selector_dark_gauss_ds_3_rd0_select
  logic [0:0] selector_dark_gauss_ds_3_rd0_select_clk;
  logic [0:0] selector_dark_gauss_ds_3_rd0_select_rst;
  logic [31:0] selector_dark_gauss_ds_3_rd0_select_d0;
  logic [31:0] selector_dark_gauss_ds_3_rd0_select_d1;
  logic [31:0] selector_dark_gauss_ds_3_rd0_select_out;
  dark_gauss_ds_3_rd0_select selector_dark_gauss_ds_3_rd0_select(.clk(selector_dark_gauss_ds_3_rd0_select_clk), .rst(selector_dark_gauss_ds_3_rd0_select_rst), .d0(selector_dark_gauss_ds_3_rd0_select_d0), .d1(selector_dark_gauss_ds_3_rd0_select_d1), .out(selector_dark_gauss_ds_3_rd0_select_out));
  assign selector_dark_gauss_ds_3_rd0_select_clk = clk;
  assign selector_dark_gauss_ds_3_rd0_select_rst = rst;
  // Bindings to selector_dark_gauss_ds_3_rd0_select

  // dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1
  logic [0:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_done;
  dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1 dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1(.clk(dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_clk), .rst(dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_rst), .start(dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_start), .done(dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_done));
  assign dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_clk = clk;
  assign dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_gauss_blur_3_dark_gauss_blur_3_update_0_write0_merged_banks_1

  // Bindings to dark_gauss_blur_3_update_0_write_wen
    // rd_0
  assign rd_0 = dark_gauss_blur_3_update_0_write_wen;

  // Bindings to dark_gauss_ds_3_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_gauss_ds_3_update_0_read_dummy;



endmodule


module dark_gauss_ds_1_dark_gauss_ds_1_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f17
  logic [0:0] f17_wen;
  logic [31:0] f17_wdata;
  logic [0:0] f17_clk;
  logic [0:0] f17_rst;
  logic [31:0] f17_rdata;
  sr_buffer_32_2527 f17(.wen(f17_wen), .wdata(f17_wdata), .clk(f17_clk), .rst(f17_rst), .rdata(f17_rdata));
  assign f17_clk = clk;
  assign f17_rst = rst;
  // Bindings to f17

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_628 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_628 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2



endmodule


module in_wire_dark_gauss_ds_2_update_0_write_wen(output [0:0] dark_gauss_ds_2_update_0_write_wen);

endmodule


module dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_631 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f314
  logic [0:0] f314_wen;
  logic [31:0] f314_wdata;
  logic [0:0] f314_clk;
  logic [0:0] f314_rst;
  logic [31:0] f314_rdata;
  sr_buffer_32_1 f314(.wen(f314_wen), .wdata(f314_wdata), .clk(f314_clk), .rst(f314_rst), .rdata(f314_rdata));
  assign f314_clk = clk;
  assign f314_rst = rst;
  // Bindings to f314

  // f316
  logic [0:0] f316_wen;
  logic [31:0] f316_wdata;
  logic [0:0] f316_clk;
  logic [0:0] f316_rst;
  logic [31:0] f316_rdata;
  sr_buffer_32_1 f316(.wen(f316_wen), .wdata(f316_wdata), .clk(f316_clk), .rst(f316_rst), .rdata(f316_rdata));
  assign f316_clk = clk;
  assign f316_rst = rst;
  // Bindings to f316

  // f318
  logic [0:0] f318_wen;
  logic [31:0] f318_wdata;
  logic [0:0] f318_clk;
  logic [0:0] f318_rst;
  logic [31:0] f318_rdata;
  sr_buffer_32_1 f318(.wen(f318_wen), .wdata(f318_wdata), .clk(f318_clk), .rst(f318_rst), .rdata(f318_rdata));
  assign f318_clk = clk;
  assign f318_rst = rst;
  // Bindings to f318

  // f320
  logic [0:0] f320_wen;
  logic [31:0] f320_wdata;
  logic [0:0] f320_clk;
  logic [0:0] f320_rst;
  logic [31:0] f320_rdata;
  sr_buffer_32_1 f320(.wen(f320_wen), .wdata(f320_wdata), .clk(f320_clk), .rst(f320_rst), .rdata(f320_rdata));
  assign f320_clk = clk;
  assign f320_rst = rst;
  // Bindings to f320

  // f322
  logic [0:0] f322_wen;
  logic [31:0] f322_wdata;
  logic [0:0] f322_clk;
  logic [0:0] f322_rst;
  logic [31:0] f322_rdata;
  sr_buffer_32_1 f322(.wen(f322_wen), .wdata(f322_wdata), .clk(f322_clk), .rst(f322_rst), .rdata(f322_rdata));
  assign f322_clk = clk;
  assign f322_rst = rst;
  // Bindings to f322

  // f324
  logic [0:0] f324_wen;
  logic [31:0] f324_wdata;
  logic [0:0] f324_clk;
  logic [0:0] f324_rst;
  logic [31:0] f324_rdata;
  sr_buffer_32_1 f324(.wen(f324_wen), .wdata(f324_wdata), .clk(f324_clk), .rst(f324_rst), .rdata(f324_rdata));
  assign f324_clk = clk;
  assign f324_rst = rst;
  // Bindings to f324

  // f326
  logic [0:0] f326_wen;
  logic [31:0] f326_wdata;
  logic [0:0] f326_clk;
  logic [0:0] f326_rst;
  logic [31:0] f326_rdata;
  sr_buffer_32_1 f326(.wen(f326_wen), .wdata(f326_wdata), .clk(f326_clk), .rst(f326_rst), .rdata(f326_rdata));
  assign f326_clk = clk;
  assign f326_rst = rst;
  // Bindings to f326

  // f328
  logic [0:0] f328_wen;
  logic [31:0] f328_wdata;
  logic [0:0] f328_clk;
  logic [0:0] f328_rst;
  logic [31:0] f328_rdata;
  sr_buffer_32_1 f328(.wen(f328_wen), .wdata(f328_wdata), .clk(f328_clk), .rst(f328_rst), .rdata(f328_rdata));
  assign f328_clk = clk;
  assign f328_rst = rst;
  // Bindings to f328

  // f330
  logic [0:0] f330_wen;
  logic [31:0] f330_wdata;
  logic [0:0] f330_clk;
  logic [0:0] f330_rst;
  logic [31:0] f330_rdata;
  sr_buffer_32_1 f330(.wen(f330_wen), .wdata(f330_wdata), .clk(f330_clk), .rst(f330_rst), .rdata(f330_rdata));
  assign f330_clk = clk;
  assign f330_rst = rst;
  // Bindings to f330

  // f332
  logic [0:0] f332_wen;
  logic [31:0] f332_wdata;
  logic [0:0] f332_clk;
  logic [0:0] f332_rst;
  logic [31:0] f332_rdata;
  sr_buffer_32_1 f332(.wen(f332_wen), .wdata(f332_wdata), .clk(f332_clk), .rst(f332_rst), .rdata(f332_rdata));
  assign f332_clk = clk;
  assign f332_rst = rst;
  // Bindings to f332

  // f334
  logic [0:0] f334_wen;
  logic [31:0] f334_wdata;
  logic [0:0] f334_clk;
  logic [0:0] f334_rst;
  logic [31:0] f334_rdata;
  sr_buffer_32_1 f334(.wen(f334_wen), .wdata(f334_wdata), .clk(f334_clk), .rst(f334_rst), .rdata(f334_rdata));
  assign f334_clk = clk;
  assign f334_rst = rst;
  // Bindings to f334

  // f336
  logic [0:0] f336_wen;
  logic [31:0] f336_wdata;
  logic [0:0] f336_clk;
  logic [0:0] f336_rst;
  logic [31:0] f336_rdata;
  sr_buffer_32_1 f336(.wen(f336_wen), .wdata(f336_wdata), .clk(f336_clk), .rst(f336_rst), .rdata(f336_rdata));
  assign f336_clk = clk;
  assign f336_rst = rst;
  // Bindings to f336

  // f338
  logic [0:0] f338_wen;
  logic [31:0] f338_wdata;
  logic [0:0] f338_clk;
  logic [0:0] f338_rst;
  logic [31:0] f338_rdata;
  sr_buffer_32_1 f338(.wen(f338_wen), .wdata(f338_wdata), .clk(f338_clk), .rst(f338_rst), .rdata(f338_rdata));
  assign f338_clk = clk;
  assign f338_rst = rst;
  // Bindings to f338

  // f340
  logic [0:0] f340_wen;
  logic [31:0] f340_wdata;
  logic [0:0] f340_clk;
  logic [0:0] f340_rst;
  logic [31:0] f340_rdata;
  sr_buffer_32_1 f340(.wen(f340_wen), .wdata(f340_wdata), .clk(f340_clk), .rst(f340_rst), .rdata(f340_rdata));
  assign f340_clk = clk;
  assign f340_rst = rst;
  // Bindings to f340

  // f342
  logic [0:0] f342_wen;
  logic [31:0] f342_wdata;
  logic [0:0] f342_clk;
  logic [0:0] f342_rst;
  logic [31:0] f342_rdata;
  sr_buffer_32_1 f342(.wen(f342_wen), .wdata(f342_wdata), .clk(f342_clk), .rst(f342_rst), .rdata(f342_rdata));
  assign f342_clk = clk;
  assign f342_rst = rst;
  // Bindings to f342

  // f344
  logic [0:0] f344_wen;
  logic [31:0] f344_wdata;
  logic [0:0] f344_clk;
  logic [0:0] f344_rst;
  logic [31:0] f344_rdata;
  sr_buffer_32_1 f344(.wen(f344_wen), .wdata(f344_wdata), .clk(f344_clk), .rst(f344_rst), .rdata(f344_rdata));
  assign f344_clk = clk;
  assign f344_rst = rst;
  // Bindings to f344

  // f346
  logic [0:0] f346_wen;
  logic [31:0] f346_wdata;
  logic [0:0] f346_clk;
  logic [0:0] f346_rst;
  logic [31:0] f346_rdata;
  sr_buffer_32_1 f346(.wen(f346_wen), .wdata(f346_wdata), .clk(f346_clk), .rst(f346_rst), .rdata(f346_rdata));
  assign f346_clk = clk;
  assign f346_rst = rst;
  // Bindings to f346

  // f348
  logic [0:0] f348_wen;
  logic [31:0] f348_wdata;
  logic [0:0] f348_clk;
  logic [0:0] f348_rst;
  logic [31:0] f348_rdata;
  sr_buffer_32_1 f348(.wen(f348_wen), .wdata(f348_wdata), .clk(f348_clk), .rst(f348_rst), .rdata(f348_rdata));
  assign f348_clk = clk;
  assign f348_rst = rst;
  // Bindings to f348

  // f350
  logic [0:0] f350_wen;
  logic [31:0] f350_wdata;
  logic [0:0] f350_clk;
  logic [0:0] f350_rst;
  logic [31:0] f350_rdata;
  sr_buffer_32_1 f350(.wen(f350_wen), .wdata(f350_wdata), .clk(f350_clk), .rst(f350_rst), .rdata(f350_rdata));
  assign f350_clk = clk;
  assign f350_rst = rst;
  // Bindings to f350

  // f352
  logic [0:0] f352_wen;
  logic [31:0] f352_wdata;
  logic [0:0] f352_clk;
  logic [0:0] f352_rst;
  logic [31:0] f352_rdata;
  sr_buffer_32_1 f352(.wen(f352_wen), .wdata(f352_wdata), .clk(f352_clk), .rst(f352_rst), .rdata(f352_rdata));
  assign f352_clk = clk;
  assign f352_rst = rst;
  // Bindings to f352

  // f354
  logic [0:0] f354_wen;
  logic [31:0] f354_wdata;
  logic [0:0] f354_clk;
  logic [0:0] f354_rst;
  logic [31:0] f354_rdata;
  sr_buffer_32_1 f354(.wen(f354_wen), .wdata(f354_wdata), .clk(f354_clk), .rst(f354_rst), .rdata(f354_rdata));
  assign f354_clk = clk;
  assign f354_rst = rst;
  // Bindings to f354

  // f356
  logic [0:0] f356_wen;
  logic [31:0] f356_wdata;
  logic [0:0] f356_clk;
  logic [0:0] f356_rst;
  logic [31:0] f356_rdata;
  sr_buffer_32_1 f356(.wen(f356_wen), .wdata(f356_wdata), .clk(f356_clk), .rst(f356_rst), .rdata(f356_rdata));
  assign f356_clk = clk;
  assign f356_rst = rst;
  // Bindings to f356

  // f358
  logic [0:0] f358_wen;
  logic [31:0] f358_wdata;
  logic [0:0] f358_clk;
  logic [0:0] f358_rst;
  logic [31:0] f358_rdata;
  sr_buffer_32_1 f358(.wen(f358_wen), .wdata(f358_wdata), .clk(f358_clk), .rst(f358_rst), .rdata(f358_rdata));
  assign f358_clk = clk;
  assign f358_rst = rst;
  // Bindings to f358

  // f360
  logic [0:0] f360_wen;
  logic [31:0] f360_wdata;
  logic [0:0] f360_clk;
  logic [0:0] f360_rst;
  logic [31:0] f360_rdata;
  sr_buffer_32_1 f360(.wen(f360_wen), .wdata(f360_wdata), .clk(f360_clk), .rst(f360_rst), .rdata(f360_rdata));
  assign f360_clk = clk;
  assign f360_rst = rst;
  // Bindings to f360

  // f362
  logic [0:0] f362_wen;
  logic [31:0] f362_wdata;
  logic [0:0] f362_clk;
  logic [0:0] f362_rst;
  logic [31:0] f362_rdata;
  sr_buffer_32_1 f362(.wen(f362_wen), .wdata(f362_wdata), .clk(f362_clk), .rst(f362_rst), .rdata(f362_rdata));
  assign f362_clk = clk;
  assign f362_rst = rst;
  // Bindings to f362

  // f364
  logic [0:0] f364_wen;
  logic [31:0] f364_wdata;
  logic [0:0] f364_clk;
  logic [0:0] f364_rst;
  logic [31:0] f364_rdata;
  sr_buffer_32_1 f364(.wen(f364_wen), .wdata(f364_wdata), .clk(f364_clk), .rst(f364_rst), .rdata(f364_rdata));
  assign f364_clk = clk;
  assign f364_rst = rst;
  // Bindings to f364

  // f366
  logic [0:0] f366_wen;
  logic [31:0] f366_wdata;
  logic [0:0] f366_clk;
  logic [0:0] f366_rst;
  logic [31:0] f366_rdata;
  sr_buffer_32_1 f366(.wen(f366_wen), .wdata(f366_wdata), .clk(f366_clk), .rst(f366_rst), .rdata(f366_rdata));
  assign f366_clk = clk;
  assign f366_rst = rst;
  // Bindings to f366

  // f368
  logic [0:0] f368_wen;
  logic [31:0] f368_wdata;
  logic [0:0] f368_clk;
  logic [0:0] f368_rst;
  logic [31:0] f368_rdata;
  sr_buffer_32_1 f368(.wen(f368_wen), .wdata(f368_wdata), .clk(f368_clk), .rst(f368_rst), .rdata(f368_rdata));
  assign f368_clk = clk;
  assign f368_rst = rst;
  // Bindings to f368

  // f370
  logic [0:0] f370_wen;
  logic [31:0] f370_wdata;
  logic [0:0] f370_clk;
  logic [0:0] f370_rst;
  logic [31:0] f370_rdata;
  sr_buffer_32_1 f370(.wen(f370_wen), .wdata(f370_wdata), .clk(f370_clk), .rst(f370_rst), .rdata(f370_rdata));
  assign f370_clk = clk;
  assign f370_rst = rst;
  // Bindings to f370

  // f372
  logic [0:0] f372_wen;
  logic [31:0] f372_wdata;
  logic [0:0] f372_clk;
  logic [0:0] f372_rst;
  logic [31:0] f372_rdata;
  sr_buffer_32_1 f372(.wen(f372_wen), .wdata(f372_wdata), .clk(f372_clk), .rst(f372_rst), .rdata(f372_rdata));
  assign f372_clk = clk;
  assign f372_rst = rst;
  // Bindings to f372

  // f374
  logic [0:0] f374_wen;
  logic [31:0] f374_wdata;
  logic [0:0] f374_clk;
  logic [0:0] f374_rst;
  logic [31:0] f374_rdata;
  sr_buffer_32_1 f374(.wen(f374_wen), .wdata(f374_wdata), .clk(f374_clk), .rst(f374_rst), .rdata(f374_rdata));
  assign f374_clk = clk;
  assign f374_rst = rst;
  // Bindings to f374

  // f376
  logic [0:0] f376_wen;
  logic [31:0] f376_wdata;
  logic [0:0] f376_clk;
  logic [0:0] f376_rst;
  logic [31:0] f376_rdata;
  sr_buffer_32_1 f376(.wen(f376_wen), .wdata(f376_wdata), .clk(f376_clk), .rst(f376_rst), .rdata(f376_rdata));
  assign f376_clk = clk;
  assign f376_rst = rst;
  // Bindings to f376

  // f378
  logic [0:0] f378_wen;
  logic [31:0] f378_wdata;
  logic [0:0] f378_clk;
  logic [0:0] f378_rst;
  logic [31:0] f378_rdata;
  sr_buffer_32_1 f378(.wen(f378_wen), .wdata(f378_wdata), .clk(f378_clk), .rst(f378_rst), .rdata(f378_rdata));
  assign f378_clk = clk;
  assign f378_rst = rst;
  // Bindings to f378

  // f380
  logic [0:0] f380_wen;
  logic [31:0] f380_wdata;
  logic [0:0] f380_clk;
  logic [0:0] f380_rst;
  logic [31:0] f380_rdata;
  sr_buffer_32_1 f380(.wen(f380_wen), .wdata(f380_wdata), .clk(f380_clk), .rst(f380_rst), .rdata(f380_rdata));
  assign f380_clk = clk;
  assign f380_rst = rst;
  // Bindings to f380

  // f382
  logic [0:0] f382_wen;
  logic [31:0] f382_wdata;
  logic [0:0] f382_clk;
  logic [0:0] f382_rst;
  logic [31:0] f382_rdata;
  sr_buffer_32_1 f382(.wen(f382_wen), .wdata(f382_wdata), .clk(f382_clk), .rst(f382_rst), .rdata(f382_rdata));
  assign f382_clk = clk;
  assign f382_rst = rst;
  // Bindings to f382

  // f384
  logic [0:0] f384_wen;
  logic [31:0] f384_wdata;
  logic [0:0] f384_clk;
  logic [0:0] f384_rst;
  logic [31:0] f384_rdata;
  sr_buffer_32_1 f384(.wen(f384_wen), .wdata(f384_wdata), .clk(f384_clk), .rst(f384_rst), .rdata(f384_rdata));
  assign f384_clk = clk;
  assign f384_rst = rst;
  // Bindings to f384

  // f386
  logic [0:0] f386_wen;
  logic [31:0] f386_wdata;
  logic [0:0] f386_clk;
  logic [0:0] f386_rst;
  logic [31:0] f386_rdata;
  sr_buffer_32_1 f386(.wen(f386_wen), .wdata(f386_wdata), .clk(f386_clk), .rst(f386_rst), .rdata(f386_rdata));
  assign f386_clk = clk;
  assign f386_rst = rst;
  // Bindings to f386

  // f388
  logic [0:0] f388_wen;
  logic [31:0] f388_wdata;
  logic [0:0] f388_clk;
  logic [0:0] f388_rst;
  logic [31:0] f388_rdata;
  sr_buffer_32_1 f388(.wen(f388_wen), .wdata(f388_wdata), .clk(f388_clk), .rst(f388_rst), .rdata(f388_rdata));
  assign f388_clk = clk;
  assign f388_rst = rst;
  // Bindings to f388

  // f390
  logic [0:0] f390_wen;
  logic [31:0] f390_wdata;
  logic [0:0] f390_clk;
  logic [0:0] f390_rst;
  logic [31:0] f390_rdata;
  sr_buffer_32_1 f390(.wen(f390_wen), .wdata(f390_wdata), .clk(f390_clk), .rst(f390_rst), .rdata(f390_rdata));
  assign f390_clk = clk;
  assign f390_rst = rst;
  // Bindings to f390

  // f392
  logic [0:0] f392_wen;
  logic [31:0] f392_wdata;
  logic [0:0] f392_clk;
  logic [0:0] f392_rst;
  logic [31:0] f392_rdata;
  sr_buffer_32_1 f392(.wen(f392_wen), .wdata(f392_wdata), .clk(f392_clk), .rst(f392_rst), .rdata(f392_rdata));
  assign f392_clk = clk;
  assign f392_rst = rst;
  // Bindings to f392

  // f394
  logic [0:0] f394_wen;
  logic [31:0] f394_wdata;
  logic [0:0] f394_clk;
  logic [0:0] f394_rst;
  logic [31:0] f394_rdata;
  sr_buffer_32_1 f394(.wen(f394_wen), .wdata(f394_wdata), .clk(f394_clk), .rst(f394_rst), .rdata(f394_rdata));
  assign f394_clk = clk;
  assign f394_rst = rst;
  // Bindings to f394

  // f396
  logic [0:0] f396_wen;
  logic [31:0] f396_wdata;
  logic [0:0] f396_clk;
  logic [0:0] f396_rst;
  logic [31:0] f396_rdata;
  sr_buffer_32_1 f396(.wen(f396_wen), .wdata(f396_wdata), .clk(f396_clk), .rst(f396_rst), .rdata(f396_rdata));
  assign f396_clk = clk;
  assign f396_rst = rst;
  // Bindings to f396

  // f398
  logic [0:0] f398_wen;
  logic [31:0] f398_wdata;
  logic [0:0] f398_clk;
  logic [0:0] f398_rst;
  logic [31:0] f398_rdata;
  sr_buffer_32_1 f398(.wen(f398_wen), .wdata(f398_wdata), .clk(f398_clk), .rst(f398_rst), .rdata(f398_rdata));
  assign f398_clk = clk;
  assign f398_rst = rst;
  // Bindings to f398

  // f400
  logic [0:0] f400_wen;
  logic [31:0] f400_wdata;
  logic [0:0] f400_clk;
  logic [0:0] f400_rst;
  logic [31:0] f400_rdata;
  sr_buffer_32_1 f400(.wen(f400_wen), .wdata(f400_wdata), .clk(f400_clk), .rst(f400_rst), .rdata(f400_rdata));
  assign f400_clk = clk;
  assign f400_rst = rst;
  // Bindings to f400

  // f402
  logic [0:0] f402_wen;
  logic [31:0] f402_wdata;
  logic [0:0] f402_clk;
  logic [0:0] f402_rst;
  logic [31:0] f402_rdata;
  sr_buffer_32_1 f402(.wen(f402_wen), .wdata(f402_wdata), .clk(f402_clk), .rst(f402_rst), .rdata(f402_rdata));
  assign f402_clk = clk;
  assign f402_rst = rst;
  // Bindings to f402

  // f404
  logic [0:0] f404_wen;
  logic [31:0] f404_wdata;
  logic [0:0] f404_clk;
  logic [0:0] f404_rst;
  logic [31:0] f404_rdata;
  sr_buffer_32_1 f404(.wen(f404_wen), .wdata(f404_wdata), .clk(f404_clk), .rst(f404_rst), .rdata(f404_rdata));
  assign f404_clk = clk;
  assign f404_rst = rst;
  // Bindings to f404

  // f406
  logic [0:0] f406_wen;
  logic [31:0] f406_wdata;
  logic [0:0] f406_clk;
  logic [0:0] f406_rst;
  logic [31:0] f406_rdata;
  sr_buffer_32_1 f406(.wen(f406_wen), .wdata(f406_wdata), .clk(f406_clk), .rst(f406_rst), .rdata(f406_rdata));
  assign f406_clk = clk;
  assign f406_rst = rst;
  // Bindings to f406

  // f408
  logic [0:0] f408_wen;
  logic [31:0] f408_wdata;
  logic [0:0] f408_clk;
  logic [0:0] f408_rst;
  logic [31:0] f408_rdata;
  sr_buffer_32_1 f408(.wen(f408_wen), .wdata(f408_wdata), .clk(f408_clk), .rst(f408_rst), .rdata(f408_rdata));
  assign f408_clk = clk;
  assign f408_rst = rst;
  // Bindings to f408

  // f410
  logic [0:0] f410_wen;
  logic [31:0] f410_wdata;
  logic [0:0] f410_clk;
  logic [0:0] f410_rst;
  logic [31:0] f410_rdata;
  sr_buffer_32_1 f410(.wen(f410_wen), .wdata(f410_wdata), .clk(f410_clk), .rst(f410_rst), .rdata(f410_rdata));
  assign f410_clk = clk;
  assign f410_rst = rst;
  // Bindings to f410

  // f412
  logic [0:0] f412_wen;
  logic [31:0] f412_wdata;
  logic [0:0] f412_clk;
  logic [0:0] f412_rst;
  logic [31:0] f412_rdata;
  sr_buffer_32_1 f412(.wen(f412_wen), .wdata(f412_wdata), .clk(f412_clk), .rst(f412_rst), .rdata(f412_rdata));
  assign f412_clk = clk;
  assign f412_rst = rst;
  // Bindings to f412

  // f414
  logic [0:0] f414_wen;
  logic [31:0] f414_wdata;
  logic [0:0] f414_clk;
  logic [0:0] f414_rst;
  logic [31:0] f414_rdata;
  sr_buffer_32_1 f414(.wen(f414_wen), .wdata(f414_wdata), .clk(f414_clk), .rst(f414_rst), .rdata(f414_rdata));
  assign f414_clk = clk;
  assign f414_rst = rst;
  // Bindings to f414

  // f416
  logic [0:0] f416_wen;
  logic [31:0] f416_wdata;
  logic [0:0] f416_clk;
  logic [0:0] f416_rst;
  logic [31:0] f416_rdata;
  sr_buffer_32_1 f416(.wen(f416_wen), .wdata(f416_wdata), .clk(f416_clk), .rst(f416_rst), .rdata(f416_rdata));
  assign f416_clk = clk;
  assign f416_rst = rst;
  // Bindings to f416

  // f418
  logic [0:0] f418_wen;
  logic [31:0] f418_wdata;
  logic [0:0] f418_clk;
  logic [0:0] f418_rst;
  logic [31:0] f418_rdata;
  sr_buffer_32_1 f418(.wen(f418_wen), .wdata(f418_wdata), .clk(f418_clk), .rst(f418_rst), .rdata(f418_rdata));
  assign f418_clk = clk;
  assign f418_rst = rst;
  // Bindings to f418

  // f420
  logic [0:0] f420_wen;
  logic [31:0] f420_wdata;
  logic [0:0] f420_clk;
  logic [0:0] f420_rst;
  logic [31:0] f420_rdata;
  sr_buffer_32_1 f420(.wen(f420_wen), .wdata(f420_wdata), .clk(f420_clk), .rst(f420_rst), .rdata(f420_rdata));
  assign f420_clk = clk;
  assign f420_rst = rst;
  // Bindings to f420

  // f422
  logic [0:0] f422_wen;
  logic [31:0] f422_wdata;
  logic [0:0] f422_clk;
  logic [0:0] f422_rst;
  logic [31:0] f422_rdata;
  sr_buffer_32_1 f422(.wen(f422_wen), .wdata(f422_wdata), .clk(f422_clk), .rst(f422_rst), .rdata(f422_rdata));
  assign f422_clk = clk;
  assign f422_rst = rst;
  // Bindings to f422

  // f424
  logic [0:0] f424_wen;
  logic [31:0] f424_wdata;
  logic [0:0] f424_clk;
  logic [0:0] f424_rst;
  logic [31:0] f424_rdata;
  sr_buffer_32_1 f424(.wen(f424_wen), .wdata(f424_wdata), .clk(f424_clk), .rst(f424_rst), .rdata(f424_rdata));
  assign f424_clk = clk;
  assign f424_rst = rst;
  // Bindings to f424

  // f426
  logic [0:0] f426_wen;
  logic [31:0] f426_wdata;
  logic [0:0] f426_clk;
  logic [0:0] f426_rst;
  logic [31:0] f426_rdata;
  sr_buffer_32_1 f426(.wen(f426_wen), .wdata(f426_wdata), .clk(f426_clk), .rst(f426_rst), .rdata(f426_rdata));
  assign f426_clk = clk;
  assign f426_rst = rst;
  // Bindings to f426

  // f428
  logic [0:0] f428_wen;
  logic [31:0] f428_wdata;
  logic [0:0] f428_clk;
  logic [0:0] f428_rst;
  logic [31:0] f428_rdata;
  sr_buffer_32_1 f428(.wen(f428_wen), .wdata(f428_wdata), .clk(f428_clk), .rst(f428_rst), .rdata(f428_rdata));
  assign f428_clk = clk;
  assign f428_rst = rst;
  // Bindings to f428

  // f430
  logic [0:0] f430_wen;
  logic [31:0] f430_wdata;
  logic [0:0] f430_clk;
  logic [0:0] f430_rst;
  logic [31:0] f430_rdata;
  sr_buffer_32_1 f430(.wen(f430_wen), .wdata(f430_wdata), .clk(f430_clk), .rst(f430_rst), .rdata(f430_rdata));
  assign f430_clk = clk;
  assign f430_rst = rst;
  // Bindings to f430

  // f432
  logic [0:0] f432_wen;
  logic [31:0] f432_wdata;
  logic [0:0] f432_clk;
  logic [0:0] f432_rst;
  logic [31:0] f432_rdata;
  sr_buffer_32_1 f432(.wen(f432_wen), .wdata(f432_wdata), .clk(f432_clk), .rst(f432_rst), .rdata(f432_rdata));
  assign f432_clk = clk;
  assign f432_rst = rst;
  // Bindings to f432

  // f434
  logic [0:0] f434_wen;
  logic [31:0] f434_wdata;
  logic [0:0] f434_clk;
  logic [0:0] f434_rst;
  logic [31:0] f434_rdata;
  sr_buffer_32_1 f434(.wen(f434_wen), .wdata(f434_wdata), .clk(f434_clk), .rst(f434_rst), .rdata(f434_rdata));
  assign f434_clk = clk;
  assign f434_rst = rst;
  // Bindings to f434

  // f436
  logic [0:0] f436_wen;
  logic [31:0] f436_wdata;
  logic [0:0] f436_clk;
  logic [0:0] f436_rst;
  logic [31:0] f436_rdata;
  sr_buffer_32_1 f436(.wen(f436_wen), .wdata(f436_wdata), .clk(f436_clk), .rst(f436_rst), .rdata(f436_rdata));
  assign f436_clk = clk;
  assign f436_rst = rst;
  // Bindings to f436

  // f438
  logic [0:0] f438_wen;
  logic [31:0] f438_wdata;
  logic [0:0] f438_clk;
  logic [0:0] f438_rst;
  logic [31:0] f438_rdata;
  sr_buffer_32_1 f438(.wen(f438_wen), .wdata(f438_wdata), .clk(f438_clk), .rst(f438_rst), .rdata(f438_rdata));
  assign f438_clk = clk;
  assign f438_rst = rst;
  // Bindings to f438

  // f440
  logic [0:0] f440_wen;
  logic [31:0] f440_wdata;
  logic [0:0] f440_clk;
  logic [0:0] f440_rst;
  logic [31:0] f440_rdata;
  sr_buffer_32_1 f440(.wen(f440_wen), .wdata(f440_wdata), .clk(f440_clk), .rst(f440_rst), .rdata(f440_rdata));
  assign f440_clk = clk;
  assign f440_rst = rst;
  // Bindings to f440

  // f442
  logic [0:0] f442_wen;
  logic [31:0] f442_wdata;
  logic [0:0] f442_clk;
  logic [0:0] f442_rst;
  logic [31:0] f442_rdata;
  sr_buffer_32_1 f442(.wen(f442_wen), .wdata(f442_wdata), .clk(f442_clk), .rst(f442_rst), .rdata(f442_rdata));
  assign f442_clk = clk;
  assign f442_rst = rst;
  // Bindings to f442

  // f444
  logic [0:0] f444_wen;
  logic [31:0] f444_wdata;
  logic [0:0] f444_clk;
  logic [0:0] f444_rst;
  logic [31:0] f444_rdata;
  sr_buffer_32_1 f444(.wen(f444_wen), .wdata(f444_wdata), .clk(f444_clk), .rst(f444_rst), .rdata(f444_rdata));
  assign f444_clk = clk;
  assign f444_rst = rst;
  // Bindings to f444

  // f446
  logic [0:0] f446_wen;
  logic [31:0] f446_wdata;
  logic [0:0] f446_clk;
  logic [0:0] f446_rst;
  logic [31:0] f446_rdata;
  sr_buffer_32_1 f446(.wen(f446_wen), .wdata(f446_wdata), .clk(f446_clk), .rst(f446_rst), .rdata(f446_rdata));
  assign f446_clk = clk;
  assign f446_rst = rst;
  // Bindings to f446

  // f448
  logic [0:0] f448_wen;
  logic [31:0] f448_wdata;
  logic [0:0] f448_clk;
  logic [0:0] f448_rst;
  logic [31:0] f448_rdata;
  sr_buffer_32_1 f448(.wen(f448_wen), .wdata(f448_wdata), .clk(f448_clk), .rst(f448_rst), .rdata(f448_rdata));
  assign f448_clk = clk;
  assign f448_rst = rst;
  // Bindings to f448

  // f450
  logic [0:0] f450_wen;
  logic [31:0] f450_wdata;
  logic [0:0] f450_clk;
  logic [0:0] f450_rst;
  logic [31:0] f450_rdata;
  sr_buffer_32_1 f450(.wen(f450_wen), .wdata(f450_wdata), .clk(f450_clk), .rst(f450_rst), .rdata(f450_rdata));
  assign f450_clk = clk;
  assign f450_rst = rst;
  // Bindings to f450

  // f452
  logic [0:0] f452_wen;
  logic [31:0] f452_wdata;
  logic [0:0] f452_clk;
  logic [0:0] f452_rst;
  logic [31:0] f452_rdata;
  sr_buffer_32_1 f452(.wen(f452_wen), .wdata(f452_wdata), .clk(f452_clk), .rst(f452_rst), .rdata(f452_rdata));
  assign f452_clk = clk;
  assign f452_rst = rst;
  // Bindings to f452

  // f454
  logic [0:0] f454_wen;
  logic [31:0] f454_wdata;
  logic [0:0] f454_clk;
  logic [0:0] f454_rst;
  logic [31:0] f454_rdata;
  sr_buffer_32_1 f454(.wen(f454_wen), .wdata(f454_wdata), .clk(f454_clk), .rst(f454_rst), .rdata(f454_rdata));
  assign f454_clk = clk;
  assign f454_rst = rst;
  // Bindings to f454

  // f456
  logic [0:0] f456_wen;
  logic [31:0] f456_wdata;
  logic [0:0] f456_clk;
  logic [0:0] f456_rst;
  logic [31:0] f456_rdata;
  sr_buffer_32_1 f456(.wen(f456_wen), .wdata(f456_wdata), .clk(f456_clk), .rst(f456_rst), .rdata(f456_rdata));
  assign f456_clk = clk;
  assign f456_rst = rst;
  // Bindings to f456

  // f458
  logic [0:0] f458_wen;
  logic [31:0] f458_wdata;
  logic [0:0] f458_clk;
  logic [0:0] f458_rst;
  logic [31:0] f458_rdata;
  sr_buffer_32_1 f458(.wen(f458_wen), .wdata(f458_wdata), .clk(f458_clk), .rst(f458_rst), .rdata(f458_rdata));
  assign f458_clk = clk;
  assign f458_rst = rst;
  // Bindings to f458

  // f460
  logic [0:0] f460_wen;
  logic [31:0] f460_wdata;
  logic [0:0] f460_clk;
  logic [0:0] f460_rst;
  logic [31:0] f460_rdata;
  sr_buffer_32_1 f460(.wen(f460_wen), .wdata(f460_wdata), .clk(f460_clk), .rst(f460_rst), .rdata(f460_rdata));
  assign f460_clk = clk;
  assign f460_rst = rst;
  // Bindings to f460

  // f462
  logic [0:0] f462_wen;
  logic [31:0] f462_wdata;
  logic [0:0] f462_clk;
  logic [0:0] f462_rst;
  logic [31:0] f462_rdata;
  sr_buffer_32_1 f462(.wen(f462_wen), .wdata(f462_wdata), .clk(f462_clk), .rst(f462_rst), .rdata(f462_rdata));
  assign f462_clk = clk;
  assign f462_rst = rst;
  // Bindings to f462

  // f464
  logic [0:0] f464_wen;
  logic [31:0] f464_wdata;
  logic [0:0] f464_clk;
  logic [0:0] f464_rst;
  logic [31:0] f464_rdata;
  sr_buffer_32_1 f464(.wen(f464_wen), .wdata(f464_wdata), .clk(f464_clk), .rst(f464_rst), .rdata(f464_rdata));
  assign f464_clk = clk;
  assign f464_rst = rst;
  // Bindings to f464

  // f466
  logic [0:0] f466_wen;
  logic [31:0] f466_wdata;
  logic [0:0] f466_clk;
  logic [0:0] f466_rst;
  logic [31:0] f466_rdata;
  sr_buffer_32_1 f466(.wen(f466_wen), .wdata(f466_wdata), .clk(f466_clk), .rst(f466_rst), .rdata(f466_rdata));
  assign f466_clk = clk;
  assign f466_rst = rst;
  // Bindings to f466

  // f468
  logic [0:0] f468_wen;
  logic [31:0] f468_wdata;
  logic [0:0] f468_clk;
  logic [0:0] f468_rst;
  logic [31:0] f468_rdata;
  sr_buffer_32_1 f468(.wen(f468_wen), .wdata(f468_wdata), .clk(f468_clk), .rst(f468_rst), .rdata(f468_rdata));
  assign f468_clk = clk;
  assign f468_rst = rst;
  // Bindings to f468

  // f470
  logic [0:0] f470_wen;
  logic [31:0] f470_wdata;
  logic [0:0] f470_clk;
  logic [0:0] f470_rst;
  logic [31:0] f470_rdata;
  sr_buffer_32_1 f470(.wen(f470_wen), .wdata(f470_wdata), .clk(f470_clk), .rst(f470_rst), .rdata(f470_rdata));
  assign f470_clk = clk;
  assign f470_rst = rst;
  // Bindings to f470

  // f472
  logic [0:0] f472_wen;
  logic [31:0] f472_wdata;
  logic [0:0] f472_clk;
  logic [0:0] f472_rst;
  logic [31:0] f472_rdata;
  sr_buffer_32_1 f472(.wen(f472_wen), .wdata(f472_wdata), .clk(f472_clk), .rst(f472_rst), .rdata(f472_rdata));
  assign f472_clk = clk;
  assign f472_rst = rst;
  // Bindings to f472

  // f474
  logic [0:0] f474_wen;
  logic [31:0] f474_wdata;
  logic [0:0] f474_clk;
  logic [0:0] f474_rst;
  logic [31:0] f474_rdata;
  sr_buffer_32_1 f474(.wen(f474_wen), .wdata(f474_wdata), .clk(f474_clk), .rst(f474_rst), .rdata(f474_rdata));
  assign f474_clk = clk;
  assign f474_rst = rst;
  // Bindings to f474

  // f476
  logic [0:0] f476_wen;
  logic [31:0] f476_wdata;
  logic [0:0] f476_clk;
  logic [0:0] f476_rst;
  logic [31:0] f476_rdata;
  sr_buffer_32_1 f476(.wen(f476_wen), .wdata(f476_wdata), .clk(f476_clk), .rst(f476_rst), .rdata(f476_rdata));
  assign f476_clk = clk;
  assign f476_rst = rst;
  // Bindings to f476

  // f478
  logic [0:0] f478_wen;
  logic [31:0] f478_wdata;
  logic [0:0] f478_clk;
  logic [0:0] f478_rst;
  logic [31:0] f478_rdata;
  sr_buffer_32_1 f478(.wen(f478_wen), .wdata(f478_wdata), .clk(f478_clk), .rst(f478_rst), .rdata(f478_rdata));
  assign f478_clk = clk;
  assign f478_rst = rst;
  // Bindings to f478

  // f480
  logic [0:0] f480_wen;
  logic [31:0] f480_wdata;
  logic [0:0] f480_clk;
  logic [0:0] f480_rst;
  logic [31:0] f480_rdata;
  sr_buffer_32_1 f480(.wen(f480_wen), .wdata(f480_wdata), .clk(f480_clk), .rst(f480_rst), .rdata(f480_rdata));
  assign f480_clk = clk;
  assign f480_rst = rst;
  // Bindings to f480

  // f482
  logic [0:0] f482_wen;
  logic [31:0] f482_wdata;
  logic [0:0] f482_clk;
  logic [0:0] f482_rst;
  logic [31:0] f482_rdata;
  sr_buffer_32_1 f482(.wen(f482_wen), .wdata(f482_wdata), .clk(f482_clk), .rst(f482_rst), .rdata(f482_rdata));
  assign f482_clk = clk;
  assign f482_rst = rst;
  // Bindings to f482

  // f484
  logic [0:0] f484_wen;
  logic [31:0] f484_wdata;
  logic [0:0] f484_clk;
  logic [0:0] f484_rst;
  logic [31:0] f484_rdata;
  sr_buffer_32_1 f484(.wen(f484_wen), .wdata(f484_wdata), .clk(f484_clk), .rst(f484_rst), .rdata(f484_rdata));
  assign f484_clk = clk;
  assign f484_rst = rst;
  // Bindings to f484

  // f486
  logic [0:0] f486_wen;
  logic [31:0] f486_wdata;
  logic [0:0] f486_clk;
  logic [0:0] f486_rst;
  logic [31:0] f486_rdata;
  sr_buffer_32_1 f486(.wen(f486_wen), .wdata(f486_wdata), .clk(f486_clk), .rst(f486_rst), .rdata(f486_rdata));
  assign f486_clk = clk;
  assign f486_rst = rst;
  // Bindings to f486

  // f488
  logic [0:0] f488_wen;
  logic [31:0] f488_wdata;
  logic [0:0] f488_clk;
  logic [0:0] f488_rst;
  logic [31:0] f488_rdata;
  sr_buffer_32_1 f488(.wen(f488_wen), .wdata(f488_wdata), .clk(f488_clk), .rst(f488_rst), .rdata(f488_rdata));
  assign f488_clk = clk;
  assign f488_rst = rst;
  // Bindings to f488

  // f490
  logic [0:0] f490_wen;
  logic [31:0] f490_wdata;
  logic [0:0] f490_clk;
  logic [0:0] f490_rst;
  logic [31:0] f490_rdata;
  sr_buffer_32_1 f490(.wen(f490_wen), .wdata(f490_wdata), .clk(f490_clk), .rst(f490_rst), .rdata(f490_rdata));
  assign f490_clk = clk;
  assign f490_rst = rst;
  // Bindings to f490

  // f492
  logic [0:0] f492_wen;
  logic [31:0] f492_wdata;
  logic [0:0] f492_clk;
  logic [0:0] f492_rst;
  logic [31:0] f492_rdata;
  sr_buffer_32_1 f492(.wen(f492_wen), .wdata(f492_wdata), .clk(f492_clk), .rst(f492_rst), .rdata(f492_rdata));
  assign f492_clk = clk;
  assign f492_rst = rst;
  // Bindings to f492

  // f494
  logic [0:0] f494_wen;
  logic [31:0] f494_wdata;
  logic [0:0] f494_clk;
  logic [0:0] f494_rst;
  logic [31:0] f494_rdata;
  sr_buffer_32_1 f494(.wen(f494_wen), .wdata(f494_wdata), .clk(f494_clk), .rst(f494_rst), .rdata(f494_rdata));
  assign f494_clk = clk;
  assign f494_rst = rst;
  // Bindings to f494

  // f496
  logic [0:0] f496_wen;
  logic [31:0] f496_wdata;
  logic [0:0] f496_clk;
  logic [0:0] f496_rst;
  logic [31:0] f496_rdata;
  sr_buffer_32_1 f496(.wen(f496_wen), .wdata(f496_wdata), .clk(f496_clk), .rst(f496_rst), .rdata(f496_rdata));
  assign f496_clk = clk;
  assign f496_rst = rst;
  // Bindings to f496

  // f498
  logic [0:0] f498_wen;
  logic [31:0] f498_wdata;
  logic [0:0] f498_clk;
  logic [0:0] f498_rst;
  logic [31:0] f498_rdata;
  sr_buffer_32_1 f498(.wen(f498_wen), .wdata(f498_wdata), .clk(f498_clk), .rst(f498_rst), .rdata(f498_rdata));
  assign f498_clk = clk;
  assign f498_rst = rst;
  // Bindings to f498

  // f500
  logic [0:0] f500_wen;
  logic [31:0] f500_wdata;
  logic [0:0] f500_clk;
  logic [0:0] f500_rst;
  logic [31:0] f500_rdata;
  sr_buffer_32_1 f500(.wen(f500_wen), .wdata(f500_wdata), .clk(f500_clk), .rst(f500_rst), .rdata(f500_rdata));
  assign f500_clk = clk;
  assign f500_rst = rst;
  // Bindings to f500

  // f502
  logic [0:0] f502_wen;
  logic [31:0] f502_wdata;
  logic [0:0] f502_clk;
  logic [0:0] f502_rst;
  logic [31:0] f502_rdata;
  sr_buffer_32_1 f502(.wen(f502_wen), .wdata(f502_wdata), .clk(f502_clk), .rst(f502_rst), .rdata(f502_rdata));
  assign f502_clk = clk;
  assign f502_rst = rst;
  // Bindings to f502

  // f504
  logic [0:0] f504_wen;
  logic [31:0] f504_wdata;
  logic [0:0] f504_clk;
  logic [0:0] f504_rst;
  logic [31:0] f504_rdata;
  sr_buffer_32_1 f504(.wen(f504_wen), .wdata(f504_wdata), .clk(f504_clk), .rst(f504_rst), .rdata(f504_rdata));
  assign f504_clk = clk;
  assign f504_rst = rst;
  // Bindings to f504

  // f506
  logic [0:0] f506_wen;
  logic [31:0] f506_wdata;
  logic [0:0] f506_clk;
  logic [0:0] f506_rst;
  logic [31:0] f506_rdata;
  sr_buffer_32_1 f506(.wen(f506_wen), .wdata(f506_wdata), .clk(f506_clk), .rst(f506_rst), .rdata(f506_rdata));
  assign f506_clk = clk;
  assign f506_rst = rst;
  // Bindings to f506

  // f508
  logic [0:0] f508_wen;
  logic [31:0] f508_wdata;
  logic [0:0] f508_clk;
  logic [0:0] f508_rst;
  logic [31:0] f508_rdata;
  sr_buffer_32_1 f508(.wen(f508_wen), .wdata(f508_wdata), .clk(f508_clk), .rst(f508_rst), .rdata(f508_rdata));
  assign f508_clk = clk;
  assign f508_rst = rst;
  // Bindings to f508

  // f510
  logic [0:0] f510_wen;
  logic [31:0] f510_wdata;
  logic [0:0] f510_clk;
  logic [0:0] f510_rst;
  logic [31:0] f510_rdata;
  sr_buffer_32_1 f510(.wen(f510_wen), .wdata(f510_wdata), .clk(f510_clk), .rst(f510_rst), .rdata(f510_rdata));
  assign f510_clk = clk;
  assign f510_rst = rst;
  // Bindings to f510

  // f512
  logic [0:0] f512_wen;
  logic [31:0] f512_wdata;
  logic [0:0] f512_clk;
  logic [0:0] f512_rst;
  logic [31:0] f512_rdata;
  sr_buffer_32_1 f512(.wen(f512_wen), .wdata(f512_wdata), .clk(f512_clk), .rst(f512_rst), .rdata(f512_rdata));
  assign f512_clk = clk;
  assign f512_rst = rst;
  // Bindings to f512

  // f514
  logic [0:0] f514_wen;
  logic [31:0] f514_wdata;
  logic [0:0] f514_clk;
  logic [0:0] f514_rst;
  logic [31:0] f514_rdata;
  sr_buffer_32_1 f514(.wen(f514_wen), .wdata(f514_wdata), .clk(f514_clk), .rst(f514_rst), .rdata(f514_rdata));
  assign f514_clk = clk;
  assign f514_rst = rst;
  // Bindings to f514

  // f516
  logic [0:0] f516_wen;
  logic [31:0] f516_wdata;
  logic [0:0] f516_clk;
  logic [0:0] f516_rst;
  logic [31:0] f516_rdata;
  sr_buffer_32_1 f516(.wen(f516_wen), .wdata(f516_wdata), .clk(f516_clk), .rst(f516_rst), .rdata(f516_rdata));
  assign f516_clk = clk;
  assign f516_rst = rst;
  // Bindings to f516

  // f518
  logic [0:0] f518_wen;
  logic [31:0] f518_wdata;
  logic [0:0] f518_clk;
  logic [0:0] f518_rst;
  logic [31:0] f518_rdata;
  sr_buffer_32_1 f518(.wen(f518_wen), .wdata(f518_wdata), .clk(f518_clk), .rst(f518_rst), .rdata(f518_rdata));
  assign f518_clk = clk;
  assign f518_rst = rst;
  // Bindings to f518

  // f520
  logic [0:0] f520_wen;
  logic [31:0] f520_wdata;
  logic [0:0] f520_clk;
  logic [0:0] f520_rst;
  logic [31:0] f520_rdata;
  sr_buffer_32_1 f520(.wen(f520_wen), .wdata(f520_wdata), .clk(f520_clk), .rst(f520_rst), .rdata(f520_rdata));
  assign f520_clk = clk;
  assign f520_rst = rst;
  // Bindings to f520

  // f522
  logic [0:0] f522_wen;
  logic [31:0] f522_wdata;
  logic [0:0] f522_clk;
  logic [0:0] f522_rst;
  logic [31:0] f522_rdata;
  sr_buffer_32_1 f522(.wen(f522_wen), .wdata(f522_wdata), .clk(f522_clk), .rst(f522_rst), .rdata(f522_rdata));
  assign f522_clk = clk;
  assign f522_rst = rst;
  // Bindings to f522

  // f524
  logic [0:0] f524_wen;
  logic [31:0] f524_wdata;
  logic [0:0] f524_clk;
  logic [0:0] f524_rst;
  logic [31:0] f524_rdata;
  sr_buffer_32_1 f524(.wen(f524_wen), .wdata(f524_wdata), .clk(f524_clk), .rst(f524_rst), .rdata(f524_rdata));
  assign f524_clk = clk;
  assign f524_rst = rst;
  // Bindings to f524

  // f526
  logic [0:0] f526_wen;
  logic [31:0] f526_wdata;
  logic [0:0] f526_clk;
  logic [0:0] f526_rst;
  logic [31:0] f526_rdata;
  sr_buffer_32_1 f526(.wen(f526_wen), .wdata(f526_wdata), .clk(f526_clk), .rst(f526_rst), .rdata(f526_rdata));
  assign f526_clk = clk;
  assign f526_rst = rst;
  // Bindings to f526

  // f528
  logic [0:0] f528_wen;
  logic [31:0] f528_wdata;
  logic [0:0] f528_clk;
  logic [0:0] f528_rst;
  logic [31:0] f528_rdata;
  sr_buffer_32_1 f528(.wen(f528_wen), .wdata(f528_wdata), .clk(f528_clk), .rst(f528_rst), .rdata(f528_rdata));
  assign f528_clk = clk;
  assign f528_rst = rst;
  // Bindings to f528

  // f530
  logic [0:0] f530_wen;
  logic [31:0] f530_wdata;
  logic [0:0] f530_clk;
  logic [0:0] f530_rst;
  logic [31:0] f530_rdata;
  sr_buffer_32_1 f530(.wen(f530_wen), .wdata(f530_wdata), .clk(f530_clk), .rst(f530_rst), .rdata(f530_rdata));
  assign f530_clk = clk;
  assign f530_rst = rst;
  // Bindings to f530

  // f532
  logic [0:0] f532_wen;
  logic [31:0] f532_wdata;
  logic [0:0] f532_clk;
  logic [0:0] f532_rst;
  logic [31:0] f532_rdata;
  sr_buffer_32_1 f532(.wen(f532_wen), .wdata(f532_wdata), .clk(f532_clk), .rst(f532_rst), .rdata(f532_rdata));
  assign f532_clk = clk;
  assign f532_rst = rst;
  // Bindings to f532

  // f534
  logic [0:0] f534_wen;
  logic [31:0] f534_wdata;
  logic [0:0] f534_clk;
  logic [0:0] f534_rst;
  logic [31:0] f534_rdata;
  sr_buffer_32_1 f534(.wen(f534_wen), .wdata(f534_wdata), .clk(f534_clk), .rst(f534_rst), .rdata(f534_rdata));
  assign f534_clk = clk;
  assign f534_rst = rst;
  // Bindings to f534

  // f536
  logic [0:0] f536_wen;
  logic [31:0] f536_wdata;
  logic [0:0] f536_clk;
  logic [0:0] f536_rst;
  logic [31:0] f536_rdata;
  sr_buffer_32_1 f536(.wen(f536_wen), .wdata(f536_wdata), .clk(f536_clk), .rst(f536_rst), .rdata(f536_rdata));
  assign f536_clk = clk;
  assign f536_rst = rst;
  // Bindings to f536

  // f538
  logic [0:0] f538_wen;
  logic [31:0] f538_wdata;
  logic [0:0] f538_clk;
  logic [0:0] f538_rst;
  logic [31:0] f538_rdata;
  sr_buffer_32_1 f538(.wen(f538_wen), .wdata(f538_wdata), .clk(f538_clk), .rst(f538_rst), .rdata(f538_rdata));
  assign f538_clk = clk;
  assign f538_rst = rst;
  // Bindings to f538

  // f540
  logic [0:0] f540_wen;
  logic [31:0] f540_wdata;
  logic [0:0] f540_clk;
  logic [0:0] f540_rst;
  logic [31:0] f540_rdata;
  sr_buffer_32_1 f540(.wen(f540_wen), .wdata(f540_wdata), .clk(f540_clk), .rst(f540_rst), .rdata(f540_rdata));
  assign f540_clk = clk;
  assign f540_rst = rst;
  // Bindings to f540

  // f542
  logic [0:0] f542_wen;
  logic [31:0] f542_wdata;
  logic [0:0] f542_clk;
  logic [0:0] f542_rst;
  logic [31:0] f542_rdata;
  sr_buffer_32_1 f542(.wen(f542_wen), .wdata(f542_wdata), .clk(f542_clk), .rst(f542_rst), .rdata(f542_rdata));
  assign f542_clk = clk;
  assign f542_rst = rst;
  // Bindings to f542

  // f544
  logic [0:0] f544_wen;
  logic [31:0] f544_wdata;
  logic [0:0] f544_clk;
  logic [0:0] f544_rst;
  logic [31:0] f544_rdata;
  sr_buffer_32_1 f544(.wen(f544_wen), .wdata(f544_wdata), .clk(f544_clk), .rst(f544_rst), .rdata(f544_rdata));
  assign f544_clk = clk;
  assign f544_rst = rst;
  // Bindings to f544

  // f546
  logic [0:0] f546_wen;
  logic [31:0] f546_wdata;
  logic [0:0] f546_clk;
  logic [0:0] f546_rst;
  logic [31:0] f546_rdata;
  sr_buffer_32_1 f546(.wen(f546_wen), .wdata(f546_wdata), .clk(f546_clk), .rst(f546_rst), .rdata(f546_rdata));
  assign f546_clk = clk;
  assign f546_rst = rst;
  // Bindings to f546

  // f548
  logic [0:0] f548_wen;
  logic [31:0] f548_wdata;
  logic [0:0] f548_clk;
  logic [0:0] f548_rst;
  logic [31:0] f548_rdata;
  sr_buffer_32_1 f548(.wen(f548_wen), .wdata(f548_wdata), .clk(f548_clk), .rst(f548_rst), .rdata(f548_rdata));
  assign f548_clk = clk;
  assign f548_rst = rst;
  // Bindings to f548

  // f550
  logic [0:0] f550_wen;
  logic [31:0] f550_wdata;
  logic [0:0] f550_clk;
  logic [0:0] f550_rst;
  logic [31:0] f550_rdata;
  sr_buffer_32_1 f550(.wen(f550_wen), .wdata(f550_wdata), .clk(f550_clk), .rst(f550_rst), .rdata(f550_rdata));
  assign f550_clk = clk;
  assign f550_rst = rst;
  // Bindings to f550

  // f552
  logic [0:0] f552_wen;
  logic [31:0] f552_wdata;
  logic [0:0] f552_clk;
  logic [0:0] f552_rst;
  logic [31:0] f552_rdata;
  sr_buffer_32_1 f552(.wen(f552_wen), .wdata(f552_wdata), .clk(f552_clk), .rst(f552_rst), .rdata(f552_rdata));
  assign f552_clk = clk;
  assign f552_rst = rst;
  // Bindings to f552

  // f554
  logic [0:0] f554_wen;
  logic [31:0] f554_wdata;
  logic [0:0] f554_clk;
  logic [0:0] f554_rst;
  logic [31:0] f554_rdata;
  sr_buffer_32_1 f554(.wen(f554_wen), .wdata(f554_wdata), .clk(f554_clk), .rst(f554_rst), .rdata(f554_rdata));
  assign f554_clk = clk;
  assign f554_rst = rst;
  // Bindings to f554

  // f556
  logic [0:0] f556_wen;
  logic [31:0] f556_wdata;
  logic [0:0] f556_clk;
  logic [0:0] f556_rst;
  logic [31:0] f556_rdata;
  sr_buffer_32_1 f556(.wen(f556_wen), .wdata(f556_wdata), .clk(f556_clk), .rst(f556_rst), .rdata(f556_rdata));
  assign f556_clk = clk;
  assign f556_rst = rst;
  // Bindings to f556

  // f558
  logic [0:0] f558_wen;
  logic [31:0] f558_wdata;
  logic [0:0] f558_clk;
  logic [0:0] f558_rst;
  logic [31:0] f558_rdata;
  sr_buffer_32_1 f558(.wen(f558_wen), .wdata(f558_wdata), .clk(f558_clk), .rst(f558_rst), .rdata(f558_rdata));
  assign f558_clk = clk;
  assign f558_rst = rst;
  // Bindings to f558

  // f560
  logic [0:0] f560_wen;
  logic [31:0] f560_wdata;
  logic [0:0] f560_clk;
  logic [0:0] f560_rst;
  logic [31:0] f560_rdata;
  sr_buffer_32_1 f560(.wen(f560_wen), .wdata(f560_wdata), .clk(f560_clk), .rst(f560_rst), .rdata(f560_rdata));
  assign f560_clk = clk;
  assign f560_rst = rst;
  // Bindings to f560

  // f562
  logic [0:0] f562_wen;
  logic [31:0] f562_wdata;
  logic [0:0] f562_clk;
  logic [0:0] f562_rst;
  logic [31:0] f562_rdata;
  sr_buffer_32_1 f562(.wen(f562_wen), .wdata(f562_wdata), .clk(f562_clk), .rst(f562_rst), .rdata(f562_rdata));
  assign f562_clk = clk;
  assign f562_rst = rst;
  // Bindings to f562

  // f564
  logic [0:0] f564_wen;
  logic [31:0] f564_wdata;
  logic [0:0] f564_clk;
  logic [0:0] f564_rst;
  logic [31:0] f564_rdata;
  sr_buffer_32_1 f564(.wen(f564_wen), .wdata(f564_wdata), .clk(f564_clk), .rst(f564_rst), .rdata(f564_rdata));
  assign f564_clk = clk;
  assign f564_rst = rst;
  // Bindings to f564

  // f566
  logic [0:0] f566_wen;
  logic [31:0] f566_wdata;
  logic [0:0] f566_clk;
  logic [0:0] f566_rst;
  logic [31:0] f566_rdata;
  sr_buffer_32_1 f566(.wen(f566_wen), .wdata(f566_wdata), .clk(f566_clk), .rst(f566_rst), .rdata(f566_rdata));
  assign f566_clk = clk;
  assign f566_rst = rst;
  // Bindings to f566

  // f568
  logic [0:0] f568_wen;
  logic [31:0] f568_wdata;
  logic [0:0] f568_clk;
  logic [0:0] f568_rst;
  logic [31:0] f568_rdata;
  sr_buffer_32_1 f568(.wen(f568_wen), .wdata(f568_wdata), .clk(f568_clk), .rst(f568_rst), .rdata(f568_rdata));
  assign f568_clk = clk;
  assign f568_rst = rst;
  // Bindings to f568

  // f570
  logic [0:0] f570_wen;
  logic [31:0] f570_wdata;
  logic [0:0] f570_clk;
  logic [0:0] f570_rst;
  logic [31:0] f570_rdata;
  sr_buffer_32_1 f570(.wen(f570_wen), .wdata(f570_wdata), .clk(f570_clk), .rst(f570_rst), .rdata(f570_rdata));
  assign f570_clk = clk;
  assign f570_rst = rst;
  // Bindings to f570

  // f572
  logic [0:0] f572_wen;
  logic [31:0] f572_wdata;
  logic [0:0] f572_clk;
  logic [0:0] f572_rst;
  logic [31:0] f572_rdata;
  sr_buffer_32_1 f572(.wen(f572_wen), .wdata(f572_wdata), .clk(f572_clk), .rst(f572_rst), .rdata(f572_rdata));
  assign f572_clk = clk;
  assign f572_rst = rst;
  // Bindings to f572

  // f574
  logic [0:0] f574_wen;
  logic [31:0] f574_wdata;
  logic [0:0] f574_clk;
  logic [0:0] f574_rst;
  logic [31:0] f574_rdata;
  sr_buffer_32_1 f574(.wen(f574_wen), .wdata(f574_wdata), .clk(f574_clk), .rst(f574_rst), .rdata(f574_rdata));
  assign f574_clk = clk;
  assign f574_rst = rst;
  // Bindings to f574

  // f576
  logic [0:0] f576_wen;
  logic [31:0] f576_wdata;
  logic [0:0] f576_clk;
  logic [0:0] f576_rst;
  logic [31:0] f576_rdata;
  sr_buffer_32_1 f576(.wen(f576_wen), .wdata(f576_wdata), .clk(f576_clk), .rst(f576_rst), .rdata(f576_rdata));
  assign f576_clk = clk;
  assign f576_rst = rst;
  // Bindings to f576

  // f578
  logic [0:0] f578_wen;
  logic [31:0] f578_wdata;
  logic [0:0] f578_clk;
  logic [0:0] f578_rst;
  logic [31:0] f578_rdata;
  sr_buffer_32_1 f578(.wen(f578_wen), .wdata(f578_wdata), .clk(f578_clk), .rst(f578_rst), .rdata(f578_rdata));
  assign f578_clk = clk;
  assign f578_rst = rst;
  // Bindings to f578

  // f580
  logic [0:0] f580_wen;
  logic [31:0] f580_wdata;
  logic [0:0] f580_clk;
  logic [0:0] f580_rst;
  logic [31:0] f580_rdata;
  sr_buffer_32_1 f580(.wen(f580_wen), .wdata(f580_wdata), .clk(f580_clk), .rst(f580_rst), .rdata(f580_rdata));
  assign f580_clk = clk;
  assign f580_rst = rst;
  // Bindings to f580

  // f582
  logic [0:0] f582_wen;
  logic [31:0] f582_wdata;
  logic [0:0] f582_clk;
  logic [0:0] f582_rst;
  logic [31:0] f582_rdata;
  sr_buffer_32_1 f582(.wen(f582_wen), .wdata(f582_wdata), .clk(f582_clk), .rst(f582_rst), .rdata(f582_rdata));
  assign f582_clk = clk;
  assign f582_rst = rst;
  // Bindings to f582

  // f584
  logic [0:0] f584_wen;
  logic [31:0] f584_wdata;
  logic [0:0] f584_clk;
  logic [0:0] f584_rst;
  logic [31:0] f584_rdata;
  sr_buffer_32_1 f584(.wen(f584_wen), .wdata(f584_wdata), .clk(f584_clk), .rst(f584_rst), .rdata(f584_rdata));
  assign f584_clk = clk;
  assign f584_rst = rst;
  // Bindings to f584

  // f586
  logic [0:0] f586_wen;
  logic [31:0] f586_wdata;
  logic [0:0] f586_clk;
  logic [0:0] f586_rst;
  logic [31:0] f586_rdata;
  sr_buffer_32_1 f586(.wen(f586_wen), .wdata(f586_wdata), .clk(f586_clk), .rst(f586_rst), .rdata(f586_rdata));
  assign f586_clk = clk;
  assign f586_rst = rst;
  // Bindings to f586

  // f588
  logic [0:0] f588_wen;
  logic [31:0] f588_wdata;
  logic [0:0] f588_clk;
  logic [0:0] f588_rst;
  logic [31:0] f588_rdata;
  sr_buffer_32_1 f588(.wen(f588_wen), .wdata(f588_wdata), .clk(f588_clk), .rst(f588_rst), .rdata(f588_rdata));
  assign f588_clk = clk;
  assign f588_rst = rst;
  // Bindings to f588

  // f590
  logic [0:0] f590_wen;
  logic [31:0] f590_wdata;
  logic [0:0] f590_clk;
  logic [0:0] f590_rst;
  logic [31:0] f590_rdata;
  sr_buffer_32_1 f590(.wen(f590_wen), .wdata(f590_wdata), .clk(f590_clk), .rst(f590_rst), .rdata(f590_rdata));
  assign f590_clk = clk;
  assign f590_rst = rst;
  // Bindings to f590

  // f592
  logic [0:0] f592_wen;
  logic [31:0] f592_wdata;
  logic [0:0] f592_clk;
  logic [0:0] f592_rst;
  logic [31:0] f592_rdata;
  sr_buffer_32_1 f592(.wen(f592_wen), .wdata(f592_wdata), .clk(f592_clk), .rst(f592_rst), .rdata(f592_rdata));
  assign f592_clk = clk;
  assign f592_rst = rst;
  // Bindings to f592

  // f594
  logic [0:0] f594_wen;
  logic [31:0] f594_wdata;
  logic [0:0] f594_clk;
  logic [0:0] f594_rst;
  logic [31:0] f594_rdata;
  sr_buffer_32_1 f594(.wen(f594_wen), .wdata(f594_wdata), .clk(f594_clk), .rst(f594_rst), .rdata(f594_rdata));
  assign f594_clk = clk;
  assign f594_rst = rst;
  // Bindings to f594

  // f596
  logic [0:0] f596_wen;
  logic [31:0] f596_wdata;
  logic [0:0] f596_clk;
  logic [0:0] f596_rst;
  logic [31:0] f596_rdata;
  sr_buffer_32_1 f596(.wen(f596_wen), .wdata(f596_wdata), .clk(f596_clk), .rst(f596_rst), .rdata(f596_rdata));
  assign f596_clk = clk;
  assign f596_rst = rst;
  // Bindings to f596

  // f598
  logic [0:0] f598_wen;
  logic [31:0] f598_wdata;
  logic [0:0] f598_clk;
  logic [0:0] f598_rst;
  logic [31:0] f598_rdata;
  sr_buffer_32_1 f598(.wen(f598_wen), .wdata(f598_wdata), .clk(f598_clk), .rst(f598_rst), .rdata(f598_rdata));
  assign f598_clk = clk;
  assign f598_rst = rst;
  // Bindings to f598

  // f600
  logic [0:0] f600_wen;
  logic [31:0] f600_wdata;
  logic [0:0] f600_clk;
  logic [0:0] f600_rst;
  logic [31:0] f600_rdata;
  sr_buffer_32_1 f600(.wen(f600_wen), .wdata(f600_wdata), .clk(f600_clk), .rst(f600_rst), .rdata(f600_rdata));
  assign f600_clk = clk;
  assign f600_rst = rst;
  // Bindings to f600

  // f602
  logic [0:0] f602_wen;
  logic [31:0] f602_wdata;
  logic [0:0] f602_clk;
  logic [0:0] f602_rst;
  logic [31:0] f602_rdata;
  sr_buffer_32_1 f602(.wen(f602_wen), .wdata(f602_wdata), .clk(f602_clk), .rst(f602_rst), .rdata(f602_rdata));
  assign f602_clk = clk;
  assign f602_rst = rst;
  // Bindings to f602

  // f604
  logic [0:0] f604_wen;
  logic [31:0] f604_wdata;
  logic [0:0] f604_clk;
  logic [0:0] f604_rst;
  logic [31:0] f604_rdata;
  sr_buffer_32_1 f604(.wen(f604_wen), .wdata(f604_wdata), .clk(f604_clk), .rst(f604_rst), .rdata(f604_rdata));
  assign f604_clk = clk;
  assign f604_rst = rst;
  // Bindings to f604

  // f606
  logic [0:0] f606_wen;
  logic [31:0] f606_wdata;
  logic [0:0] f606_clk;
  logic [0:0] f606_rst;
  logic [31:0] f606_rdata;
  sr_buffer_32_1 f606(.wen(f606_wen), .wdata(f606_wdata), .clk(f606_clk), .rst(f606_rst), .rdata(f606_rdata));
  assign f606_clk = clk;
  assign f606_rst = rst;
  // Bindings to f606

  // f608
  logic [0:0] f608_wen;
  logic [31:0] f608_wdata;
  logic [0:0] f608_clk;
  logic [0:0] f608_rst;
  logic [31:0] f608_rdata;
  sr_buffer_32_1 f608(.wen(f608_wen), .wdata(f608_wdata), .clk(f608_clk), .rst(f608_rst), .rdata(f608_rdata));
  assign f608_clk = clk;
  assign f608_rst = rst;
  // Bindings to f608

  // f610
  logic [0:0] f610_wen;
  logic [31:0] f610_wdata;
  logic [0:0] f610_clk;
  logic [0:0] f610_rst;
  logic [31:0] f610_rdata;
  sr_buffer_32_1 f610(.wen(f610_wen), .wdata(f610_wdata), .clk(f610_clk), .rst(f610_rst), .rdata(f610_rdata));
  assign f610_clk = clk;
  assign f610_rst = rst;
  // Bindings to f610

  // f612
  logic [0:0] f612_wen;
  logic [31:0] f612_wdata;
  logic [0:0] f612_clk;
  logic [0:0] f612_rst;
  logic [31:0] f612_rdata;
  sr_buffer_32_1 f612(.wen(f612_wen), .wdata(f612_wdata), .clk(f612_clk), .rst(f612_rst), .rdata(f612_rdata));
  assign f612_clk = clk;
  assign f612_rst = rst;
  // Bindings to f612

  // f614
  logic [0:0] f614_wen;
  logic [31:0] f614_wdata;
  logic [0:0] f614_clk;
  logic [0:0] f614_rst;
  logic [31:0] f614_rdata;
  sr_buffer_32_1 f614(.wen(f614_wen), .wdata(f614_wdata), .clk(f614_clk), .rst(f614_rst), .rdata(f614_rdata));
  assign f614_clk = clk;
  assign f614_rst = rst;
  // Bindings to f614

  // f616
  logic [0:0] f616_wen;
  logic [31:0] f616_wdata;
  logic [0:0] f616_clk;
  logic [0:0] f616_rst;
  logic [31:0] f616_rdata;
  sr_buffer_32_1 f616(.wen(f616_wen), .wdata(f616_wdata), .clk(f616_clk), .rst(f616_rst), .rdata(f616_rdata));
  assign f616_clk = clk;
  assign f616_rst = rst;
  // Bindings to f616

  // f618
  logic [0:0] f618_wen;
  logic [31:0] f618_wdata;
  logic [0:0] f618_clk;
  logic [0:0] f618_rst;
  logic [31:0] f618_rdata;
  sr_buffer_32_1 f618(.wen(f618_wen), .wdata(f618_wdata), .clk(f618_clk), .rst(f618_rst), .rdata(f618_rdata));
  assign f618_clk = clk;
  assign f618_rst = rst;
  // Bindings to f618

  // f620
  logic [0:0] f620_wen;
  logic [31:0] f620_wdata;
  logic [0:0] f620_clk;
  logic [0:0] f620_rst;
  logic [31:0] f620_rdata;
  sr_buffer_32_1 f620(.wen(f620_wen), .wdata(f620_wdata), .clk(f620_clk), .rst(f620_rst), .rdata(f620_rdata));
  assign f620_clk = clk;
  assign f620_rst = rst;
  // Bindings to f620

  // f622
  logic [0:0] f622_wen;
  logic [31:0] f622_wdata;
  logic [0:0] f622_clk;
  logic [0:0] f622_rst;
  logic [31:0] f622_rdata;
  sr_buffer_32_1 f622(.wen(f622_wen), .wdata(f622_wdata), .clk(f622_clk), .rst(f622_rst), .rdata(f622_rdata));
  assign f622_clk = clk;
  assign f622_rst = rst;
  // Bindings to f622

  // f624
  logic [0:0] f624_wen;
  logic [31:0] f624_wdata;
  logic [0:0] f624_clk;
  logic [0:0] f624_rst;
  logic [31:0] f624_rdata;
  sr_buffer_32_1 f624(.wen(f624_wen), .wdata(f624_wdata), .clk(f624_clk), .rst(f624_rst), .rdata(f624_rdata));
  assign f624_clk = clk;
  assign f624_rst = rst;
  // Bindings to f624

  // f626
  logic [0:0] f626_wen;
  logic [31:0] f626_wdata;
  logic [0:0] f626_clk;
  logic [0:0] f626_rst;
  logic [31:0] f626_rdata;
  sr_buffer_32_1 f626(.wen(f626_wen), .wdata(f626_wdata), .clk(f626_clk), .rst(f626_rst), .rdata(f626_rdata));
  assign f626_clk = clk;
  assign f626_rst = rst;
  // Bindings to f626



endmodule


module bright_gauss_blur_1_bright_gauss_blur_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_gauss_blur_1_update_0_write_wen(output [0:0] bright_gauss_blur_1_update_0_write_wen);

endmodule


module in_wire_bright_gauss_blur_1_update_0_write_wdata(output [31:0] bright_gauss_blur_1_update_0_write_wdata);

endmodule


module bright_gauss_ds_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_gauss_ds_1_update_0_read_dummy(output [31:0] bright_gauss_ds_1_update_0_read_dummy);

endmodule


module out_wire_bright_gauss_ds_1_update_0_read_rdata(input [31:0] bright_gauss_ds_1_update_0_read_rdata);

endmodule


module bright_gauss_blur_2_bright_gauss_blur_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_gauss_ds_2_update_0_read_dummy(output [31:0] bright_gauss_ds_2_update_0_read_dummy);

endmodule


module out_wire_bright_gauss_ds_2_update_0_read_rdata(input [31:0] bright_gauss_ds_2_update_0_read_rdata);

endmodule


module bright_gauss_ds_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_bright_gauss_blur_2_update_0_write_wen(output [0:0] bright_gauss_blur_2_update_0_write_wen);

endmodule


module in_wire_bright_gauss_blur_2_update_0_write_wdata(output [31:0] bright_gauss_blur_2_update_0_write_wdata);

endmodule


module bright_gauss_ds_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_gauss_ds_1_update_0_write_wen, input [31:0] bright_gauss_ds_1_update_0_write_wdata, input [287:0] bright_gauss_blur_2_update_0_read_dummy, output [287:0] bright_gauss_blur_2_update_0_read_rdata, input [31:0] bright_laplace_diff_1_update_0_read_dummy, output [31:0] bright_laplace_diff_1_update_0_read_rdata, input [31:0] bright_laplace_us_0_update_0_read_dummy, output [31:0] bright_laplace_us_0_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;
  logic [31:0] rd_6;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;
  reg [31:0] rd_6_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;
      rd_6_stage_1 <= rd_6;


    end

  end


  // Data processing units...
  // bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_clk;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_rst;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_start;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_done;
  bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0 bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0(.clk(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_clk), .rst(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_rst), .start(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_start), .done(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_done));
  assign bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_clk = clk;
  assign bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0_rst = rst;
  // Bindings to bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_to_bright_laplace_us_0_rd0

  // selector_bright_gauss_blur_2_rd0_select
  logic [0:0] selector_bright_gauss_blur_2_rd0_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd0_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd0_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd0_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd0_select_out;
  bright_gauss_blur_2_rd0_select selector_bright_gauss_blur_2_rd0_select(.clk(selector_bright_gauss_blur_2_rd0_select_clk), .rst(selector_bright_gauss_blur_2_rd0_select_rst), .d0(selector_bright_gauss_blur_2_rd0_select_d0), .d1(selector_bright_gauss_blur_2_rd0_select_d1), .out(selector_bright_gauss_blur_2_rd0_select_out));
  assign selector_bright_gauss_blur_2_rd0_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd0_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd0_select

  // selector_bright_gauss_blur_2_rd1_select
  logic [0:0] selector_bright_gauss_blur_2_rd1_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd1_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd1_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd1_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd1_select_out;
  bright_gauss_blur_2_rd1_select selector_bright_gauss_blur_2_rd1_select(.clk(selector_bright_gauss_blur_2_rd1_select_clk), .rst(selector_bright_gauss_blur_2_rd1_select_rst), .d0(selector_bright_gauss_blur_2_rd1_select_d0), .d1(selector_bright_gauss_blur_2_rd1_select_d1), .out(selector_bright_gauss_blur_2_rd1_select_out));
  assign selector_bright_gauss_blur_2_rd1_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd1_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd1_select

  // Bindings to bright_gauss_ds_1_update_0_write_wen
    // rd_0
  assign rd_0 = bright_gauss_ds_1_update_0_write_wen;

  // selector_bright_gauss_blur_2_rd2_select
  logic [0:0] selector_bright_gauss_blur_2_rd2_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd2_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd2_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd2_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd2_select_out;
  bright_gauss_blur_2_rd2_select selector_bright_gauss_blur_2_rd2_select(.clk(selector_bright_gauss_blur_2_rd2_select_clk), .rst(selector_bright_gauss_blur_2_rd2_select_rst), .d0(selector_bright_gauss_blur_2_rd2_select_d0), .d1(selector_bright_gauss_blur_2_rd2_select_d1), .out(selector_bright_gauss_blur_2_rd2_select_out));
  assign selector_bright_gauss_blur_2_rd2_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd2_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd2_select

  // selector_bright_gauss_blur_2_rd3_select
  logic [0:0] selector_bright_gauss_blur_2_rd3_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd3_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd3_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd3_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd3_select_out;
  bright_gauss_blur_2_rd3_select selector_bright_gauss_blur_2_rd3_select(.clk(selector_bright_gauss_blur_2_rd3_select_clk), .rst(selector_bright_gauss_blur_2_rd3_select_rst), .d0(selector_bright_gauss_blur_2_rd3_select_d0), .d1(selector_bright_gauss_blur_2_rd3_select_d1), .out(selector_bright_gauss_blur_2_rd3_select_out));
  assign selector_bright_gauss_blur_2_rd3_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd3_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd3_select

  // selector_bright_gauss_blur_2_rd4_select
  logic [0:0] selector_bright_gauss_blur_2_rd4_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd4_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd4_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd4_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd4_select_out;
  bright_gauss_blur_2_rd4_select selector_bright_gauss_blur_2_rd4_select(.clk(selector_bright_gauss_blur_2_rd4_select_clk), .rst(selector_bright_gauss_blur_2_rd4_select_rst), .d0(selector_bright_gauss_blur_2_rd4_select_d0), .d1(selector_bright_gauss_blur_2_rd4_select_d1), .out(selector_bright_gauss_blur_2_rd4_select_out));
  assign selector_bright_gauss_blur_2_rd4_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd4_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd4_select

  // selector_bright_gauss_blur_2_rd5_select
  logic [0:0] selector_bright_gauss_blur_2_rd5_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd5_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd5_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd5_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd5_select_out;
  bright_gauss_blur_2_rd5_select selector_bright_gauss_blur_2_rd5_select(.clk(selector_bright_gauss_blur_2_rd5_select_clk), .rst(selector_bright_gauss_blur_2_rd5_select_rst), .d0(selector_bright_gauss_blur_2_rd5_select_d0), .d1(selector_bright_gauss_blur_2_rd5_select_d1), .out(selector_bright_gauss_blur_2_rd5_select_out));
  assign selector_bright_gauss_blur_2_rd5_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd5_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd5_select

  // selector_bright_gauss_blur_2_rd6_select
  logic [0:0] selector_bright_gauss_blur_2_rd6_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd6_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd6_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd6_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd6_select_out;
  bright_gauss_blur_2_rd6_select selector_bright_gauss_blur_2_rd6_select(.clk(selector_bright_gauss_blur_2_rd6_select_clk), .rst(selector_bright_gauss_blur_2_rd6_select_rst), .d0(selector_bright_gauss_blur_2_rd6_select_d0), .d1(selector_bright_gauss_blur_2_rd6_select_d1), .out(selector_bright_gauss_blur_2_rd6_select_out));
  assign selector_bright_gauss_blur_2_rd6_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd6_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd6_select

  // selector_bright_gauss_blur_2_rd7_select
  logic [0:0] selector_bright_gauss_blur_2_rd7_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd7_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd7_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd7_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd7_select_out;
  bright_gauss_blur_2_rd7_select selector_bright_gauss_blur_2_rd7_select(.clk(selector_bright_gauss_blur_2_rd7_select_clk), .rst(selector_bright_gauss_blur_2_rd7_select_rst), .d0(selector_bright_gauss_blur_2_rd7_select_d0), .d1(selector_bright_gauss_blur_2_rd7_select_d1), .out(selector_bright_gauss_blur_2_rd7_select_out));
  assign selector_bright_gauss_blur_2_rd7_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd7_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd7_select

  // selector_bright_gauss_blur_2_rd8_select
  logic [0:0] selector_bright_gauss_blur_2_rd8_select_clk;
  logic [0:0] selector_bright_gauss_blur_2_rd8_select_rst;
  logic [31:0] selector_bright_gauss_blur_2_rd8_select_d0;
  logic [31:0] selector_bright_gauss_blur_2_rd8_select_d1;
  logic [31:0] selector_bright_gauss_blur_2_rd8_select_out;
  bright_gauss_blur_2_rd8_select selector_bright_gauss_blur_2_rd8_select(.clk(selector_bright_gauss_blur_2_rd8_select_clk), .rst(selector_bright_gauss_blur_2_rd8_select_rst), .d0(selector_bright_gauss_blur_2_rd8_select_d0), .d1(selector_bright_gauss_blur_2_rd8_select_d1), .out(selector_bright_gauss_blur_2_rd8_select_out));
  assign selector_bright_gauss_blur_2_rd8_select_clk = clk;
  assign selector_bright_gauss_blur_2_rd8_select_rst = rst;
  // Bindings to selector_bright_gauss_blur_2_rd8_select

  // selector_bright_laplace_us_0_rd0_select
  logic [0:0] selector_bright_laplace_us_0_rd0_select_clk;
  logic [0:0] selector_bright_laplace_us_0_rd0_select_rst;
  logic [31:0] selector_bright_laplace_us_0_rd0_select_d0;
  logic [31:0] selector_bright_laplace_us_0_rd0_select_d1;
  logic [31:0] selector_bright_laplace_us_0_rd0_select_out;
  bright_laplace_us_0_rd0_select selector_bright_laplace_us_0_rd0_select(.clk(selector_bright_laplace_us_0_rd0_select_clk), .rst(selector_bright_laplace_us_0_rd0_select_rst), .d0(selector_bright_laplace_us_0_rd0_select_d0), .d1(selector_bright_laplace_us_0_rd0_select_d1), .out(selector_bright_laplace_us_0_rd0_select_out));
  assign selector_bright_laplace_us_0_rd0_select_clk = clk;
  assign selector_bright_laplace_us_0_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_us_0_rd0_select

  // selector_bright_laplace_diff_1_rd0_select
  logic [0:0] selector_bright_laplace_diff_1_rd0_select_clk;
  logic [0:0] selector_bright_laplace_diff_1_rd0_select_rst;
  logic [31:0] selector_bright_laplace_diff_1_rd0_select_d0;
  logic [31:0] selector_bright_laplace_diff_1_rd0_select_d1;
  logic [31:0] selector_bright_laplace_diff_1_rd0_select_out;
  bright_laplace_diff_1_rd0_select selector_bright_laplace_diff_1_rd0_select(.clk(selector_bright_laplace_diff_1_rd0_select_clk), .rst(selector_bright_laplace_diff_1_rd0_select_rst), .d0(selector_bright_laplace_diff_1_rd0_select_d0), .d1(selector_bright_laplace_diff_1_rd0_select_d1), .out(selector_bright_laplace_diff_1_rd0_select_out));
  assign selector_bright_laplace_diff_1_rd0_select_clk = clk;
  assign selector_bright_laplace_diff_1_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_diff_1_rd0_select

  // Bindings to bright_gauss_ds_1_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_gauss_ds_1_update_0_write_wdata;

  // Bindings to bright_gauss_blur_2_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_gauss_blur_2_update_0_read_dummy;

  // Bindings to bright_gauss_blur_2_update_0_read_rdata
    // wr_3
  assign bright_gauss_blur_2_update_0_read_rdata = rd_2;

  // Bindings to bright_laplace_diff_1_update_0_read_dummy
    // rd_4
  assign rd_4 = bright_laplace_diff_1_update_0_read_dummy;

  // Bindings to bright_laplace_diff_1_update_0_read_rdata
    // wr_5
  assign bright_laplace_diff_1_update_0_read_rdata = rd_4;

  // Bindings to bright_laplace_us_0_update_0_read_dummy
    // rd_6
  assign rd_6 = bright_laplace_us_0_update_0_read_dummy;

  // Bindings to bright_laplace_us_0_update_0_read_rdata
    // wr_7
  assign bright_laplace_us_0_update_0_read_rdata = rd_6;

  // bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10_clk;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10_rst;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10_start;
  logic [0:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10_done;
  bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10 bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10(.clk(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10_clk), .rst(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10_rst), .start(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10_start), .done(bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10_done));
  assign bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10_clk = clk;
  assign bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to bright_gauss_ds_1_bright_gauss_ds_1_update_0_write0_merged_banks_10



endmodule


module bright_gauss_ds_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] bright_gauss_ds_3_update_0_write_wen, input [31:0] fused_level_3_update_0_read_dummy, output [31:0] fused_level_3_update_0_read_rdata, output [31:0] bright_laplace_us_2_update_0_read_rdata, input [31:0] bright_gauss_ds_3_update_0_write_wdata, input [31:0] bright_laplace_us_2_update_0_read_dummy);

  logic [0:0] rd_0;
  logic [31:0] rd_2;
  logic [31:0] rd_1;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_2_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_2_stage_1 <= rd_2;
      rd_1_stage_1 <= rd_1;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_clk;
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_rst;
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_start;
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_done;
  bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0 bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0(.clk(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_clk), .rst(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_rst), .start(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_start), .done(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_done));
  assign bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_clk = clk;
  assign bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0_rst = rst;
  // Bindings to bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_to_bright_laplace_us_2_rd0

  // bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_start;
  logic [0:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_done;
  bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1 bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1(.clk(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_clk), .rst(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_rst), .start(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_start), .done(bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_done));
  assign bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_clk = clk;
  assign bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to bright_gauss_ds_3_bright_gauss_ds_3_update_0_write0_merged_banks_1

  // selector_bright_laplace_us_2_rd0_select
  logic [0:0] selector_bright_laplace_us_2_rd0_select_clk;
  logic [0:0] selector_bright_laplace_us_2_rd0_select_rst;
  logic [31:0] selector_bright_laplace_us_2_rd0_select_d0;
  logic [31:0] selector_bright_laplace_us_2_rd0_select_d1;
  logic [31:0] selector_bright_laplace_us_2_rd0_select_out;
  bright_laplace_us_2_rd0_select selector_bright_laplace_us_2_rd0_select(.clk(selector_bright_laplace_us_2_rd0_select_clk), .rst(selector_bright_laplace_us_2_rd0_select_rst), .d0(selector_bright_laplace_us_2_rd0_select_d0), .d1(selector_bright_laplace_us_2_rd0_select_d1), .out(selector_bright_laplace_us_2_rd0_select_out));
  assign selector_bright_laplace_us_2_rd0_select_clk = clk;
  assign selector_bright_laplace_us_2_rd0_select_rst = rst;
  // Bindings to selector_bright_laplace_us_2_rd0_select

  // Bindings to bright_gauss_ds_3_update_0_write_wen
    // rd_0
  assign rd_0 = bright_gauss_ds_3_update_0_write_wen;

  // selector_fused_level_3_rd0_select
  logic [0:0] selector_fused_level_3_rd0_select_clk;
  logic [0:0] selector_fused_level_3_rd0_select_rst;
  logic [31:0] selector_fused_level_3_rd0_select_d0;
  logic [31:0] selector_fused_level_3_rd0_select_d1;
  logic [31:0] selector_fused_level_3_rd0_select_out;
  fused_level_3_rd0_select selector_fused_level_3_rd0_select(.clk(selector_fused_level_3_rd0_select_clk), .rst(selector_fused_level_3_rd0_select_rst), .d0(selector_fused_level_3_rd0_select_d0), .d1(selector_fused_level_3_rd0_select_d1), .out(selector_fused_level_3_rd0_select_out));
  assign selector_fused_level_3_rd0_select_clk = clk;
  assign selector_fused_level_3_rd0_select_rst = rst;
  // Bindings to selector_fused_level_3_rd0_select

  // Bindings to fused_level_3_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_3_update_0_read_dummy;

  // Bindings to fused_level_3_update_0_read_rdata
    // wr_5
  assign fused_level_3_update_0_read_rdata = rd_4;

  // Bindings to bright_laplace_us_2_update_0_read_rdata
    // wr_3
  assign bright_laplace_us_2_update_0_read_rdata = rd_2;

  // Bindings to bright_gauss_ds_3_update_0_write_wdata
    // rd_1
  assign rd_1 = bright_gauss_ds_3_update_0_write_wdata;

  // Bindings to bright_laplace_us_2_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_laplace_us_2_update_0_read_dummy;



endmodule


module sr_buffer_32_312(input [0:0] wen, input [31:0] wdata, input [0:0] clk, input [0:0] rst, output [31:0] rdata);
  localparam DEPTH = 312;

  reg [31:0] data [311:0];

  reg [31:0] rdata_d;

  reg [8:0] waddr;

  wire [8:0] raddr;

  assign raddr = DEPTH - 1;

  assign rdata = rdata_d;

  always @(posedge clk) begin
    if (rst) begin
      waddr <= 0;
    end else begin
      if (wen) begin
        data[waddr] <= wdata;
        waddr <= (waddr + 1) % DEPTH;
      end

      rdata_d <= data[(waddr + raddr) % DEPTH];
    end
  end

endmodule


module in_wire_bright_laplace_diff_0_update_0_write_wen(output [0:0] bright_laplace_diff_0_update_0_write_wen);

endmodule


module bright_laplace_diff_0_bright_laplace_diff_0_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_bright_laplace_diff_0_update_0_write_wdata(output [31:0] bright_laplace_diff_0_update_0_write_wdata);

endmodule


module in_wire_fused_level_0_update_0_read_dummy(output [31:0] fused_level_0_update_0_read_dummy);

endmodule


module out_wire_fused_level_0_update_0_read_rdata(input [31:0] fused_level_0_update_0_read_rdata);

endmodule


module in_wire_bright_weights_normed_gauss_ds_3_update_0_write_wdata(output [31:0] bright_weights_normed_gauss_ds_3_update_0_write_wdata);

endmodule


module in_wire_dark_laplace_diff_1_update_0_write_wen(output [0:0] dark_laplace_diff_1_update_0_write_wen);

endmodule


module in_wire_dark_laplace_diff_1_update_0_write_wdata(output [31:0] dark_laplace_diff_1_update_0_write_wdata);

endmodule


module in_wire_dark_laplace_diff_2_update_0_write_wen(output [0:0] dark_laplace_diff_2_update_0_write_wen);

endmodule


module in_wire_dark_laplace_diff_2_update_0_write_wdata(output [31:0] dark_laplace_diff_2_update_0_write_wdata);

endmodule


module in_wire_dark_laplace_us_0_update_0_write_wen(output [0:0] dark_laplace_us_0_update_0_write_wen);

endmodule


module in_wire_dark_laplace_us_0_update_0_write_wdata(output [31:0] dark_laplace_us_0_update_0_write_wdata);

endmodule


module dark_laplace_diff_0_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_gauss_ds_3_update_0_write_wen(output [0:0] dark_weights_normed_gauss_ds_3_update_0_write_wen);

endmodule


module fused_level_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_gauss_ds_3_update_0_write_wdata(output [31:0] dark_weights_normed_gauss_ds_3_update_0_write_wdata);

endmodule


module final_merged_0_final_merged_0_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_final_merged_0_update_0_write_wen(output [0:0] final_merged_0_update_0_write_wen);

endmodule


module in_wire_final_merged_0_update_0_write_wdata(output [31:0] final_merged_0_update_0_write_wdata);

endmodule


module pyramid_synthetic_exposure_fusion_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_pyramid_synthetic_exposure_fusion_update_0_read_dummy(output [31:0] pyramid_synthetic_exposure_fusion_update_0_read_dummy);

endmodule


module out_wire_pyramid_synthetic_exposure_fusion_update_0_read_rdata(input [31:0] pyramid_synthetic_exposure_fusion_update_0_read_rdata);

endmodule


module final_merged_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] pyramid_synthetic_exposure_fusion_update_0_read_dummy, input [0:0] final_merged_0_update_0_write_wen, input [31:0] final_merged_0_update_0_write_wdata, output [31:0] pyramid_synthetic_exposure_fusion_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to pyramid_synthetic_exposure_fusion_update_0_read_dummy
    // rd_2
  assign rd_2 = pyramid_synthetic_exposure_fusion_update_0_read_dummy;

  // Bindings to final_merged_0_update_0_write_wen
    // rd_0
  assign rd_0 = final_merged_0_update_0_write_wen;

  // final_merged_0_final_merged_0_update_0_write0_merged_banks_1
  logic [0:0] final_merged_0_final_merged_0_update_0_write0_merged_banks_1_clk;
  logic [0:0] final_merged_0_final_merged_0_update_0_write0_merged_banks_1_rst;
  logic [0:0] final_merged_0_final_merged_0_update_0_write0_merged_banks_1_start;
  logic [0:0] final_merged_0_final_merged_0_update_0_write0_merged_banks_1_done;
  final_merged_0_final_merged_0_update_0_write0_merged_banks_1 final_merged_0_final_merged_0_update_0_write0_merged_banks_1(.clk(final_merged_0_final_merged_0_update_0_write0_merged_banks_1_clk), .rst(final_merged_0_final_merged_0_update_0_write0_merged_banks_1_rst), .start(final_merged_0_final_merged_0_update_0_write0_merged_banks_1_start), .done(final_merged_0_final_merged_0_update_0_write0_merged_banks_1_done));
  assign final_merged_0_final_merged_0_update_0_write0_merged_banks_1_clk = clk;
  assign final_merged_0_final_merged_0_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to final_merged_0_final_merged_0_update_0_write0_merged_banks_1

  // selector_pyramid_synthetic_exposure_fusion_rd0_select
  logic [0:0] selector_pyramid_synthetic_exposure_fusion_rd0_select_clk;
  logic [0:0] selector_pyramid_synthetic_exposure_fusion_rd0_select_rst;
  logic [31:0] selector_pyramid_synthetic_exposure_fusion_rd0_select_d0;
  logic [31:0] selector_pyramid_synthetic_exposure_fusion_rd0_select_d1;
  logic [31:0] selector_pyramid_synthetic_exposure_fusion_rd0_select_out;
  pyramid_synthetic_exposure_fusion_rd0_select selector_pyramid_synthetic_exposure_fusion_rd0_select(.clk(selector_pyramid_synthetic_exposure_fusion_rd0_select_clk), .rst(selector_pyramid_synthetic_exposure_fusion_rd0_select_rst), .d0(selector_pyramid_synthetic_exposure_fusion_rd0_select_d0), .d1(selector_pyramid_synthetic_exposure_fusion_rd0_select_d1), .out(selector_pyramid_synthetic_exposure_fusion_rd0_select_out));
  assign selector_pyramid_synthetic_exposure_fusion_rd0_select_clk = clk;
  assign selector_pyramid_synthetic_exposure_fusion_rd0_select_rst = rst;
  // Bindings to selector_pyramid_synthetic_exposure_fusion_rd0_select

  // Bindings to final_merged_0_update_0_write_wdata
    // rd_1
  assign rd_1 = final_merged_0_update_0_write_wdata;

  // Bindings to pyramid_synthetic_exposure_fusion_update_0_read_rdata
    // wr_3
  assign pyramid_synthetic_exposure_fusion_update_0_read_rdata = rd_2;



endmodule


module in_wire_final_merged_1_update_0_write_wen(output [0:0] final_merged_1_update_0_write_wen);

endmodule


module final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f422
  logic [0:0] f422_wen;
  logic [31:0] f422_wdata;
  logic [0:0] f422_clk;
  logic [0:0] f422_rst;
  logic [31:0] f422_rdata;
  sr_buffer_32_1 f422(.wen(f422_wen), .wdata(f422_wdata), .clk(f422_clk), .rst(f422_rst), .rdata(f422_rdata));
  assign f422_clk = clk;
  assign f422_rst = rst;
  // Bindings to f422

  // f420
  logic [0:0] f420_wen;
  logic [31:0] f420_wdata;
  logic [0:0] f420_clk;
  logic [0:0] f420_rst;
  logic [31:0] f420_rdata;
  sr_buffer_32_1 f420(.wen(f420_wen), .wdata(f420_wdata), .clk(f420_clk), .rst(f420_rst), .rdata(f420_rdata));
  assign f420_clk = clk;
  assign f420_rst = rst;
  // Bindings to f420

  // f416
  logic [0:0] f416_wen;
  logic [31:0] f416_wdata;
  logic [0:0] f416_clk;
  logic [0:0] f416_rst;
  logic [31:0] f416_rdata;
  sr_buffer_32_1 f416(.wen(f416_wen), .wdata(f416_wdata), .clk(f416_clk), .rst(f416_rst), .rdata(f416_rdata));
  assign f416_clk = clk;
  assign f416_rst = rst;
  // Bindings to f416

  // f418
  logic [0:0] f418_wen;
  logic [31:0] f418_wdata;
  logic [0:0] f418_clk;
  logic [0:0] f418_rst;
  logic [31:0] f418_rdata;
  sr_buffer_32_1 f418(.wen(f418_wen), .wdata(f418_wdata), .clk(f418_clk), .rst(f418_rst), .rdata(f418_rdata));
  assign f418_clk = clk;
  assign f418_rst = rst;
  // Bindings to f418

  // f414
  logic [0:0] f414_wen;
  logic [31:0] f414_wdata;
  logic [0:0] f414_clk;
  logic [0:0] f414_rst;
  logic [31:0] f414_rdata;
  sr_buffer_32_1 f414(.wen(f414_wen), .wdata(f414_wdata), .clk(f414_clk), .rst(f414_rst), .rdata(f414_rdata));
  assign f414_clk = clk;
  assign f414_rst = rst;
  // Bindings to f414

  // f410
  logic [0:0] f410_wen;
  logic [31:0] f410_wdata;
  logic [0:0] f410_clk;
  logic [0:0] f410_rst;
  logic [31:0] f410_rdata;
  sr_buffer_32_1 f410(.wen(f410_wen), .wdata(f410_wdata), .clk(f410_clk), .rst(f410_rst), .rdata(f410_rdata));
  assign f410_clk = clk;
  assign f410_rst = rst;
  // Bindings to f410

  // f412
  logic [0:0] f412_wen;
  logic [31:0] f412_wdata;
  logic [0:0] f412_clk;
  logic [0:0] f412_rst;
  logic [31:0] f412_rdata;
  sr_buffer_32_1 f412(.wen(f412_wen), .wdata(f412_wdata), .clk(f412_clk), .rst(f412_rst), .rdata(f412_rdata));
  assign f412_clk = clk;
  assign f412_rst = rst;
  // Bindings to f412

  // f406
  logic [0:0] f406_wen;
  logic [31:0] f406_wdata;
  logic [0:0] f406_clk;
  logic [0:0] f406_rst;
  logic [31:0] f406_rdata;
  sr_buffer_32_1 f406(.wen(f406_wen), .wdata(f406_wdata), .clk(f406_clk), .rst(f406_rst), .rdata(f406_rdata));
  assign f406_clk = clk;
  assign f406_rst = rst;
  // Bindings to f406

  // f408
  logic [0:0] f408_wen;
  logic [31:0] f408_wdata;
  logic [0:0] f408_clk;
  logic [0:0] f408_rst;
  logic [31:0] f408_rdata;
  sr_buffer_32_1 f408(.wen(f408_wen), .wdata(f408_wdata), .clk(f408_clk), .rst(f408_rst), .rdata(f408_rdata));
  assign f408_clk = clk;
  assign f408_rst = rst;
  // Bindings to f408

  // f400
  logic [0:0] f400_wen;
  logic [31:0] f400_wdata;
  logic [0:0] f400_clk;
  logic [0:0] f400_rst;
  logic [31:0] f400_rdata;
  sr_buffer_32_1 f400(.wen(f400_wen), .wdata(f400_wdata), .clk(f400_clk), .rst(f400_rst), .rdata(f400_rdata));
  assign f400_clk = clk;
  assign f400_rst = rst;
  // Bindings to f400

  // f404
  logic [0:0] f404_wen;
  logic [31:0] f404_wdata;
  logic [0:0] f404_clk;
  logic [0:0] f404_rst;
  logic [31:0] f404_rdata;
  sr_buffer_32_1 f404(.wen(f404_wen), .wdata(f404_wdata), .clk(f404_clk), .rst(f404_rst), .rdata(f404_rdata));
  assign f404_clk = clk;
  assign f404_rst = rst;
  // Bindings to f404

  // f402
  logic [0:0] f402_wen;
  logic [31:0] f402_wdata;
  logic [0:0] f402_clk;
  logic [0:0] f402_rst;
  logic [31:0] f402_rdata;
  sr_buffer_32_1 f402(.wen(f402_wen), .wdata(f402_wdata), .clk(f402_clk), .rst(f402_rst), .rdata(f402_rdata));
  assign f402_clk = clk;
  assign f402_rst = rst;
  // Bindings to f402

  // f398
  logic [0:0] f398_wen;
  logic [31:0] f398_wdata;
  logic [0:0] f398_clk;
  logic [0:0] f398_rst;
  logic [31:0] f398_rdata;
  sr_buffer_32_1 f398(.wen(f398_wen), .wdata(f398_wdata), .clk(f398_clk), .rst(f398_rst), .rdata(f398_rdata));
  assign f398_clk = clk;
  assign f398_rst = rst;
  // Bindings to f398

  // f396
  logic [0:0] f396_wen;
  logic [31:0] f396_wdata;
  logic [0:0] f396_clk;
  logic [0:0] f396_rst;
  logic [31:0] f396_rdata;
  sr_buffer_32_1 f396(.wen(f396_wen), .wdata(f396_wdata), .clk(f396_clk), .rst(f396_rst), .rdata(f396_rdata));
  assign f396_clk = clk;
  assign f396_rst = rst;
  // Bindings to f396

  // f394
  logic [0:0] f394_wen;
  logic [31:0] f394_wdata;
  logic [0:0] f394_clk;
  logic [0:0] f394_rst;
  logic [31:0] f394_rdata;
  sr_buffer_32_1 f394(.wen(f394_wen), .wdata(f394_wdata), .clk(f394_clk), .rst(f394_rst), .rdata(f394_rdata));
  assign f394_clk = clk;
  assign f394_rst = rst;
  // Bindings to f394

  // f390
  logic [0:0] f390_wen;
  logic [31:0] f390_wdata;
  logic [0:0] f390_clk;
  logic [0:0] f390_rst;
  logic [31:0] f390_rdata;
  sr_buffer_32_1 f390(.wen(f390_wen), .wdata(f390_wdata), .clk(f390_clk), .rst(f390_rst), .rdata(f390_rdata));
  assign f390_clk = clk;
  assign f390_rst = rst;
  // Bindings to f390

  // f392
  logic [0:0] f392_wen;
  logic [31:0] f392_wdata;
  logic [0:0] f392_clk;
  logic [0:0] f392_rst;
  logic [31:0] f392_rdata;
  sr_buffer_32_1 f392(.wen(f392_wen), .wdata(f392_wdata), .clk(f392_clk), .rst(f392_rst), .rdata(f392_rdata));
  assign f392_clk = clk;
  assign f392_rst = rst;
  // Bindings to f392

  // f388
  logic [0:0] f388_wen;
  logic [31:0] f388_wdata;
  logic [0:0] f388_clk;
  logic [0:0] f388_rst;
  logic [31:0] f388_rdata;
  sr_buffer_32_1 f388(.wen(f388_wen), .wdata(f388_wdata), .clk(f388_clk), .rst(f388_rst), .rdata(f388_rdata));
  assign f388_clk = clk;
  assign f388_rst = rst;
  // Bindings to f388

  // f384
  logic [0:0] f384_wen;
  logic [31:0] f384_wdata;
  logic [0:0] f384_clk;
  logic [0:0] f384_rst;
  logic [31:0] f384_rdata;
  sr_buffer_32_1 f384(.wen(f384_wen), .wdata(f384_wdata), .clk(f384_clk), .rst(f384_rst), .rdata(f384_rdata));
  assign f384_clk = clk;
  assign f384_rst = rst;
  // Bindings to f384

  // f386
  logic [0:0] f386_wen;
  logic [31:0] f386_wdata;
  logic [0:0] f386_clk;
  logic [0:0] f386_rst;
  logic [31:0] f386_rdata;
  sr_buffer_32_1 f386(.wen(f386_wen), .wdata(f386_wdata), .clk(f386_clk), .rst(f386_rst), .rdata(f386_rdata));
  assign f386_clk = clk;
  assign f386_rst = rst;
  // Bindings to f386

  // f376
  logic [0:0] f376_wen;
  logic [31:0] f376_wdata;
  logic [0:0] f376_clk;
  logic [0:0] f376_rst;
  logic [31:0] f376_rdata;
  sr_buffer_32_1 f376(.wen(f376_wen), .wdata(f376_wdata), .clk(f376_clk), .rst(f376_rst), .rdata(f376_rdata));
  assign f376_clk = clk;
  assign f376_rst = rst;
  // Bindings to f376

  // f382
  logic [0:0] f382_wen;
  logic [31:0] f382_wdata;
  logic [0:0] f382_clk;
  logic [0:0] f382_rst;
  logic [31:0] f382_rdata;
  sr_buffer_32_1 f382(.wen(f382_wen), .wdata(f382_wdata), .clk(f382_clk), .rst(f382_rst), .rdata(f382_rdata));
  assign f382_clk = clk;
  assign f382_rst = rst;
  // Bindings to f382

  // f380
  logic [0:0] f380_wen;
  logic [31:0] f380_wdata;
  logic [0:0] f380_clk;
  logic [0:0] f380_rst;
  logic [31:0] f380_rdata;
  sr_buffer_32_1 f380(.wen(f380_wen), .wdata(f380_wdata), .clk(f380_clk), .rst(f380_rst), .rdata(f380_rdata));
  assign f380_clk = clk;
  assign f380_rst = rst;
  // Bindings to f380

  // f378
  logic [0:0] f378_wen;
  logic [31:0] f378_wdata;
  logic [0:0] f378_clk;
  logic [0:0] f378_rst;
  logic [31:0] f378_rdata;
  sr_buffer_32_1 f378(.wen(f378_wen), .wdata(f378_wdata), .clk(f378_clk), .rst(f378_rst), .rdata(f378_rdata));
  assign f378_clk = clk;
  assign f378_rst = rst;
  // Bindings to f378

  // f374
  logic [0:0] f374_wen;
  logic [31:0] f374_wdata;
  logic [0:0] f374_clk;
  logic [0:0] f374_rst;
  logic [31:0] f374_rdata;
  sr_buffer_32_1 f374(.wen(f374_wen), .wdata(f374_wdata), .clk(f374_clk), .rst(f374_rst), .rdata(f374_rdata));
  assign f374_clk = clk;
  assign f374_rst = rst;
  // Bindings to f374

  // f372
  logic [0:0] f372_wen;
  logic [31:0] f372_wdata;
  logic [0:0] f372_clk;
  logic [0:0] f372_rst;
  logic [31:0] f372_rdata;
  sr_buffer_32_1 f372(.wen(f372_wen), .wdata(f372_wdata), .clk(f372_clk), .rst(f372_rst), .rdata(f372_rdata));
  assign f372_clk = clk;
  assign f372_rst = rst;
  // Bindings to f372

  // f370
  logic [0:0] f370_wen;
  logic [31:0] f370_wdata;
  logic [0:0] f370_clk;
  logic [0:0] f370_rst;
  logic [31:0] f370_rdata;
  sr_buffer_32_1 f370(.wen(f370_wen), .wdata(f370_wdata), .clk(f370_clk), .rst(f370_rst), .rdata(f370_rdata));
  assign f370_clk = clk;
  assign f370_rst = rst;
  // Bindings to f370

  // f366
  logic [0:0] f366_wen;
  logic [31:0] f366_wdata;
  logic [0:0] f366_clk;
  logic [0:0] f366_rst;
  logic [31:0] f366_rdata;
  sr_buffer_32_1 f366(.wen(f366_wen), .wdata(f366_wdata), .clk(f366_clk), .rst(f366_rst), .rdata(f366_rdata));
  assign f366_clk = clk;
  assign f366_rst = rst;
  // Bindings to f366

  // f368
  logic [0:0] f368_wen;
  logic [31:0] f368_wdata;
  logic [0:0] f368_clk;
  logic [0:0] f368_rst;
  logic [31:0] f368_rdata;
  sr_buffer_32_1 f368(.wen(f368_wen), .wdata(f368_wdata), .clk(f368_clk), .rst(f368_rst), .rdata(f368_rdata));
  assign f368_clk = clk;
  assign f368_rst = rst;
  // Bindings to f368

  // f356
  logic [0:0] f356_wen;
  logic [31:0] f356_wdata;
  logic [0:0] f356_clk;
  logic [0:0] f356_rst;
  logic [31:0] f356_rdata;
  sr_buffer_32_1 f356(.wen(f356_wen), .wdata(f356_wdata), .clk(f356_clk), .rst(f356_rst), .rdata(f356_rdata));
  assign f356_clk = clk;
  assign f356_rst = rst;
  // Bindings to f356

  // f364
  logic [0:0] f364_wen;
  logic [31:0] f364_wdata;
  logic [0:0] f364_clk;
  logic [0:0] f364_rst;
  logic [31:0] f364_rdata;
  sr_buffer_32_1 f364(.wen(f364_wen), .wdata(f364_wdata), .clk(f364_clk), .rst(f364_rst), .rdata(f364_rdata));
  assign f364_clk = clk;
  assign f364_rst = rst;
  // Bindings to f364

  // f362
  logic [0:0] f362_wen;
  logic [31:0] f362_wdata;
  logic [0:0] f362_clk;
  logic [0:0] f362_rst;
  logic [31:0] f362_rdata;
  sr_buffer_32_1 f362(.wen(f362_wen), .wdata(f362_wdata), .clk(f362_clk), .rst(f362_rst), .rdata(f362_rdata));
  assign f362_clk = clk;
  assign f362_rst = rst;
  // Bindings to f362

  // f358
  logic [0:0] f358_wen;
  logic [31:0] f358_wdata;
  logic [0:0] f358_clk;
  logic [0:0] f358_rst;
  logic [31:0] f358_rdata;
  sr_buffer_32_1 f358(.wen(f358_wen), .wdata(f358_wdata), .clk(f358_clk), .rst(f358_rst), .rdata(f358_rdata));
  assign f358_clk = clk;
  assign f358_rst = rst;
  // Bindings to f358

  // f360
  logic [0:0] f360_wen;
  logic [31:0] f360_wdata;
  logic [0:0] f360_clk;
  logic [0:0] f360_rst;
  logic [31:0] f360_rdata;
  sr_buffer_32_1 f360(.wen(f360_wen), .wdata(f360_wdata), .clk(f360_clk), .rst(f360_rst), .rdata(f360_rdata));
  assign f360_clk = clk;
  assign f360_rst = rst;
  // Bindings to f360

  // f354
  logic [0:0] f354_wen;
  logic [31:0] f354_wdata;
  logic [0:0] f354_clk;
  logic [0:0] f354_rst;
  logic [31:0] f354_rdata;
  sr_buffer_32_1 f354(.wen(f354_wen), .wdata(f354_wdata), .clk(f354_clk), .rst(f354_rst), .rdata(f354_rdata));
  assign f354_clk = clk;
  assign f354_rst = rst;
  // Bindings to f354

  // f352
  logic [0:0] f352_wen;
  logic [31:0] f352_wdata;
  logic [0:0] f352_clk;
  logic [0:0] f352_rst;
  logic [31:0] f352_rdata;
  sr_buffer_32_1 f352(.wen(f352_wen), .wdata(f352_wdata), .clk(f352_clk), .rst(f352_rst), .rdata(f352_rdata));
  assign f352_clk = clk;
  assign f352_rst = rst;
  // Bindings to f352

  // f346
  logic [0:0] f346_wen;
  logic [31:0] f346_wdata;
  logic [0:0] f346_clk;
  logic [0:0] f346_rst;
  logic [31:0] f346_rdata;
  sr_buffer_32_1 f346(.wen(f346_wen), .wdata(f346_wdata), .clk(f346_clk), .rst(f346_rst), .rdata(f346_rdata));
  assign f346_clk = clk;
  assign f346_rst = rst;
  // Bindings to f346

  // f350
  logic [0:0] f350_wen;
  logic [31:0] f350_wdata;
  logic [0:0] f350_clk;
  logic [0:0] f350_rst;
  logic [31:0] f350_rdata;
  sr_buffer_32_1 f350(.wen(f350_wen), .wdata(f350_wdata), .clk(f350_clk), .rst(f350_rst), .rdata(f350_rdata));
  assign f350_clk = clk;
  assign f350_rst = rst;
  // Bindings to f350

  // f348
  logic [0:0] f348_wen;
  logic [31:0] f348_wdata;
  logic [0:0] f348_clk;
  logic [0:0] f348_rst;
  logic [31:0] f348_rdata;
  sr_buffer_32_1 f348(.wen(f348_wen), .wdata(f348_wdata), .clk(f348_clk), .rst(f348_rst), .rdata(f348_rdata));
  assign f348_clk = clk;
  assign f348_rst = rst;
  // Bindings to f348

  // f344
  logic [0:0] f344_wen;
  logic [31:0] f344_wdata;
  logic [0:0] f344_clk;
  logic [0:0] f344_rst;
  logic [31:0] f344_rdata;
  sr_buffer_32_1 f344(.wen(f344_wen), .wdata(f344_wdata), .clk(f344_clk), .rst(f344_rst), .rdata(f344_rdata));
  assign f344_clk = clk;
  assign f344_rst = rst;
  // Bindings to f344

  // f342
  logic [0:0] f342_wen;
  logic [31:0] f342_wdata;
  logic [0:0] f342_clk;
  logic [0:0] f342_rst;
  logic [31:0] f342_rdata;
  sr_buffer_32_1 f342(.wen(f342_wen), .wdata(f342_wdata), .clk(f342_clk), .rst(f342_rst), .rdata(f342_rdata));
  assign f342_clk = clk;
  assign f342_rst = rst;
  // Bindings to f342

  // f340
  logic [0:0] f340_wen;
  logic [31:0] f340_wdata;
  logic [0:0] f340_clk;
  logic [0:0] f340_rst;
  logic [31:0] f340_rdata;
  sr_buffer_32_1 f340(.wen(f340_wen), .wdata(f340_wdata), .clk(f340_clk), .rst(f340_rst), .rdata(f340_rdata));
  assign f340_clk = clk;
  assign f340_rst = rst;
  // Bindings to f340

  // f330
  logic [0:0] f330_wen;
  logic [31:0] f330_wdata;
  logic [0:0] f330_clk;
  logic [0:0] f330_rst;
  logic [31:0] f330_rdata;
  sr_buffer_32_1 f330(.wen(f330_wen), .wdata(f330_wdata), .clk(f330_clk), .rst(f330_rst), .rdata(f330_rdata));
  assign f330_clk = clk;
  assign f330_rst = rst;
  // Bindings to f330

  // f338
  logic [0:0] f338_wen;
  logic [31:0] f338_wdata;
  logic [0:0] f338_clk;
  logic [0:0] f338_rst;
  logic [31:0] f338_rdata;
  sr_buffer_32_1 f338(.wen(f338_wen), .wdata(f338_wdata), .clk(f338_clk), .rst(f338_rst), .rdata(f338_rdata));
  assign f338_clk = clk;
  assign f338_rst = rst;
  // Bindings to f338

  // f336
  logic [0:0] f336_wen;
  logic [31:0] f336_wdata;
  logic [0:0] f336_clk;
  logic [0:0] f336_rst;
  logic [31:0] f336_rdata;
  sr_buffer_32_1 f336(.wen(f336_wen), .wdata(f336_wdata), .clk(f336_clk), .rst(f336_rst), .rdata(f336_rdata));
  assign f336_clk = clk;
  assign f336_rst = rst;
  // Bindings to f336

  // f332
  logic [0:0] f332_wen;
  logic [31:0] f332_wdata;
  logic [0:0] f332_clk;
  logic [0:0] f332_rst;
  logic [31:0] f332_rdata;
  sr_buffer_32_1 f332(.wen(f332_wen), .wdata(f332_wdata), .clk(f332_clk), .rst(f332_rst), .rdata(f332_rdata));
  assign f332_clk = clk;
  assign f332_rst = rst;
  // Bindings to f332

  // f334
  logic [0:0] f334_wen;
  logic [31:0] f334_wdata;
  logic [0:0] f334_clk;
  logic [0:0] f334_rst;
  logic [31:0] f334_rdata;
  sr_buffer_32_1 f334(.wen(f334_wen), .wdata(f334_wdata), .clk(f334_clk), .rst(f334_rst), .rdata(f334_rdata));
  assign f334_clk = clk;
  assign f334_rst = rst;
  // Bindings to f334

  // f328
  logic [0:0] f328_wen;
  logic [31:0] f328_wdata;
  logic [0:0] f328_clk;
  logic [0:0] f328_rst;
  logic [31:0] f328_rdata;
  sr_buffer_32_1 f328(.wen(f328_wen), .wdata(f328_wdata), .clk(f328_clk), .rst(f328_rst), .rdata(f328_rdata));
  assign f328_clk = clk;
  assign f328_rst = rst;
  // Bindings to f328

  // f324
  logic [0:0] f324_wen;
  logic [31:0] f324_wdata;
  logic [0:0] f324_clk;
  logic [0:0] f324_rst;
  logic [31:0] f324_rdata;
  sr_buffer_32_1 f324(.wen(f324_wen), .wdata(f324_wdata), .clk(f324_clk), .rst(f324_rst), .rdata(f324_rdata));
  assign f324_clk = clk;
  assign f324_rst = rst;
  // Bindings to f324

  // f326
  logic [0:0] f326_wen;
  logic [31:0] f326_wdata;
  logic [0:0] f326_clk;
  logic [0:0] f326_rst;
  logic [31:0] f326_rdata;
  sr_buffer_32_1 f326(.wen(f326_wen), .wdata(f326_wdata), .clk(f326_clk), .rst(f326_rst), .rdata(f326_rdata));
  assign f326_clk = clk;
  assign f326_rst = rst;
  // Bindings to f326

  // f320
  logic [0:0] f320_wen;
  logic [31:0] f320_wdata;
  logic [0:0] f320_clk;
  logic [0:0] f320_rst;
  logic [31:0] f320_rdata;
  sr_buffer_32_1 f320(.wen(f320_wen), .wdata(f320_wdata), .clk(f320_clk), .rst(f320_rst), .rdata(f320_rdata));
  assign f320_clk = clk;
  assign f320_rst = rst;
  // Bindings to f320

  // f322
  logic [0:0] f322_wen;
  logic [31:0] f322_wdata;
  logic [0:0] f322_clk;
  logic [0:0] f322_rst;
  logic [31:0] f322_rdata;
  sr_buffer_32_1 f322(.wen(f322_wen), .wdata(f322_wdata), .clk(f322_clk), .rst(f322_rst), .rdata(f322_rdata));
  assign f322_clk = clk;
  assign f322_rst = rst;
  // Bindings to f322

  // f318
  logic [0:0] f318_wen;
  logic [31:0] f318_wdata;
  logic [0:0] f318_clk;
  logic [0:0] f318_rst;
  logic [31:0] f318_rdata;
  sr_buffer_32_1 f318(.wen(f318_wen), .wdata(f318_wdata), .clk(f318_clk), .rst(f318_rst), .rdata(f318_rdata));
  assign f318_clk = clk;
  assign f318_rst = rst;
  // Bindings to f318

  // f316
  logic [0:0] f316_wen;
  logic [31:0] f316_wdata;
  logic [0:0] f316_clk;
  logic [0:0] f316_rst;
  logic [31:0] f316_rdata;
  sr_buffer_32_1 f316(.wen(f316_wen), .wdata(f316_wdata), .clk(f316_clk), .rst(f316_rst), .rdata(f316_rdata));
  assign f316_clk = clk;
  assign f316_rst = rst;
  // Bindings to f316

  // f314
  logic [0:0] f314_wen;
  logic [31:0] f314_wdata;
  logic [0:0] f314_clk;
  logic [0:0] f314_rst;
  logic [31:0] f314_rdata;
  sr_buffer_32_1 f314(.wen(f314_wen), .wdata(f314_wdata), .clk(f314_clk), .rst(f314_rst), .rdata(f314_rdata));
  assign f314_clk = clk;
  assign f314_rst = rst;
  // Bindings to f314

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f424
  logic [0:0] f424_wen;
  logic [31:0] f424_wdata;
  logic [0:0] f424_clk;
  logic [0:0] f424_rst;
  logic [31:0] f424_rdata;
  sr_buffer_32_1 f424(.wen(f424_wen), .wdata(f424_wdata), .clk(f424_clk), .rst(f424_rst), .rdata(f424_rdata));
  assign f424_clk = clk;
  assign f424_rst = rst;
  // Bindings to f424

  // f426
  logic [0:0] f426_wen;
  logic [31:0] f426_wdata;
  logic [0:0] f426_clk;
  logic [0:0] f426_rst;
  logic [31:0] f426_rdata;
  sr_buffer_32_1 f426(.wen(f426_wen), .wdata(f426_wdata), .clk(f426_clk), .rst(f426_rst), .rdata(f426_rdata));
  assign f426_clk = clk;
  assign f426_rst = rst;
  // Bindings to f426

  // f428
  logic [0:0] f428_wen;
  logic [31:0] f428_wdata;
  logic [0:0] f428_clk;
  logic [0:0] f428_rst;
  logic [31:0] f428_rdata;
  sr_buffer_32_1 f428(.wen(f428_wen), .wdata(f428_wdata), .clk(f428_clk), .rst(f428_rst), .rdata(f428_rdata));
  assign f428_clk = clk;
  assign f428_rst = rst;
  // Bindings to f428

  // f430
  logic [0:0] f430_wen;
  logic [31:0] f430_wdata;
  logic [0:0] f430_clk;
  logic [0:0] f430_rst;
  logic [31:0] f430_rdata;
  sr_buffer_32_1 f430(.wen(f430_wen), .wdata(f430_wdata), .clk(f430_clk), .rst(f430_rst), .rdata(f430_rdata));
  assign f430_clk = clk;
  assign f430_rst = rst;
  // Bindings to f430

  // f432
  logic [0:0] f432_wen;
  logic [31:0] f432_wdata;
  logic [0:0] f432_clk;
  logic [0:0] f432_rst;
  logic [31:0] f432_rdata;
  sr_buffer_32_1 f432(.wen(f432_wen), .wdata(f432_wdata), .clk(f432_clk), .rst(f432_rst), .rdata(f432_rdata));
  assign f432_clk = clk;
  assign f432_rst = rst;
  // Bindings to f432

  // f434
  logic [0:0] f434_wen;
  logic [31:0] f434_wdata;
  logic [0:0] f434_clk;
  logic [0:0] f434_rst;
  logic [31:0] f434_rdata;
  sr_buffer_32_1 f434(.wen(f434_wen), .wdata(f434_wdata), .clk(f434_clk), .rst(f434_rst), .rdata(f434_rdata));
  assign f434_clk = clk;
  assign f434_rst = rst;
  // Bindings to f434

  // f436
  logic [0:0] f436_wen;
  logic [31:0] f436_wdata;
  logic [0:0] f436_clk;
  logic [0:0] f436_rst;
  logic [31:0] f436_rdata;
  sr_buffer_32_1 f436(.wen(f436_wen), .wdata(f436_wdata), .clk(f436_clk), .rst(f436_rst), .rdata(f436_rdata));
  assign f436_clk = clk;
  assign f436_rst = rst;
  // Bindings to f436

  // f438
  logic [0:0] f438_wen;
  logic [31:0] f438_wdata;
  logic [0:0] f438_clk;
  logic [0:0] f438_rst;
  logic [31:0] f438_rdata;
  sr_buffer_32_1 f438(.wen(f438_wen), .wdata(f438_wdata), .clk(f438_clk), .rst(f438_rst), .rdata(f438_rdata));
  assign f438_clk = clk;
  assign f438_rst = rst;
  // Bindings to f438

  // f440
  logic [0:0] f440_wen;
  logic [31:0] f440_wdata;
  logic [0:0] f440_clk;
  logic [0:0] f440_rst;
  logic [31:0] f440_rdata;
  sr_buffer_32_1 f440(.wen(f440_wen), .wdata(f440_wdata), .clk(f440_clk), .rst(f440_rst), .rdata(f440_rdata));
  assign f440_clk = clk;
  assign f440_rst = rst;
  // Bindings to f440

  // f442
  logic [0:0] f442_wen;
  logic [31:0] f442_wdata;
  logic [0:0] f442_clk;
  logic [0:0] f442_rst;
  logic [31:0] f442_rdata;
  sr_buffer_32_1 f442(.wen(f442_wen), .wdata(f442_wdata), .clk(f442_clk), .rst(f442_rst), .rdata(f442_rdata));
  assign f442_clk = clk;
  assign f442_rst = rst;
  // Bindings to f442

  // f444
  logic [0:0] f444_wen;
  logic [31:0] f444_wdata;
  logic [0:0] f444_clk;
  logic [0:0] f444_rst;
  logic [31:0] f444_rdata;
  sr_buffer_32_1 f444(.wen(f444_wen), .wdata(f444_wdata), .clk(f444_clk), .rst(f444_rst), .rdata(f444_rdata));
  assign f444_clk = clk;
  assign f444_rst = rst;
  // Bindings to f444

  // f446
  logic [0:0] f446_wen;
  logic [31:0] f446_wdata;
  logic [0:0] f446_clk;
  logic [0:0] f446_rst;
  logic [31:0] f446_rdata;
  sr_buffer_32_1 f446(.wen(f446_wen), .wdata(f446_wdata), .clk(f446_clk), .rst(f446_rst), .rdata(f446_rdata));
  assign f446_clk = clk;
  assign f446_rst = rst;
  // Bindings to f446

  // f448
  logic [0:0] f448_wen;
  logic [31:0] f448_wdata;
  logic [0:0] f448_clk;
  logic [0:0] f448_rst;
  logic [31:0] f448_rdata;
  sr_buffer_32_1 f448(.wen(f448_wen), .wdata(f448_wdata), .clk(f448_clk), .rst(f448_rst), .rdata(f448_rdata));
  assign f448_clk = clk;
  assign f448_rst = rst;
  // Bindings to f448

  // f450
  logic [0:0] f450_wen;
  logic [31:0] f450_wdata;
  logic [0:0] f450_clk;
  logic [0:0] f450_rst;
  logic [31:0] f450_rdata;
  sr_buffer_32_1 f450(.wen(f450_wen), .wdata(f450_wdata), .clk(f450_clk), .rst(f450_rst), .rdata(f450_rdata));
  assign f450_clk = clk;
  assign f450_rst = rst;
  // Bindings to f450

  // f452
  logic [0:0] f452_wen;
  logic [31:0] f452_wdata;
  logic [0:0] f452_clk;
  logic [0:0] f452_rst;
  logic [31:0] f452_rdata;
  sr_buffer_32_1 f452(.wen(f452_wen), .wdata(f452_wdata), .clk(f452_clk), .rst(f452_rst), .rdata(f452_rdata));
  assign f452_clk = clk;
  assign f452_rst = rst;
  // Bindings to f452

  // f454
  logic [0:0] f454_wen;
  logic [31:0] f454_wdata;
  logic [0:0] f454_clk;
  logic [0:0] f454_rst;
  logic [31:0] f454_rdata;
  sr_buffer_32_1 f454(.wen(f454_wen), .wdata(f454_wdata), .clk(f454_clk), .rst(f454_rst), .rdata(f454_rdata));
  assign f454_clk = clk;
  assign f454_rst = rst;
  // Bindings to f454

  // f456
  logic [0:0] f456_wen;
  logic [31:0] f456_wdata;
  logic [0:0] f456_clk;
  logic [0:0] f456_rst;
  logic [31:0] f456_rdata;
  sr_buffer_32_1 f456(.wen(f456_wen), .wdata(f456_wdata), .clk(f456_clk), .rst(f456_rst), .rdata(f456_rdata));
  assign f456_clk = clk;
  assign f456_rst = rst;
  // Bindings to f456

  // f458
  logic [0:0] f458_wen;
  logic [31:0] f458_wdata;
  logic [0:0] f458_clk;
  logic [0:0] f458_rst;
  logic [31:0] f458_rdata;
  sr_buffer_32_1 f458(.wen(f458_wen), .wdata(f458_wdata), .clk(f458_clk), .rst(f458_rst), .rdata(f458_rdata));
  assign f458_clk = clk;
  assign f458_rst = rst;
  // Bindings to f458

  // f460
  logic [0:0] f460_wen;
  logic [31:0] f460_wdata;
  logic [0:0] f460_clk;
  logic [0:0] f460_rst;
  logic [31:0] f460_rdata;
  sr_buffer_32_1 f460(.wen(f460_wen), .wdata(f460_wdata), .clk(f460_clk), .rst(f460_rst), .rdata(f460_rdata));
  assign f460_clk = clk;
  assign f460_rst = rst;
  // Bindings to f460

  // f462
  logic [0:0] f462_wen;
  logic [31:0] f462_wdata;
  logic [0:0] f462_clk;
  logic [0:0] f462_rst;
  logic [31:0] f462_rdata;
  sr_buffer_32_1 f462(.wen(f462_wen), .wdata(f462_wdata), .clk(f462_clk), .rst(f462_rst), .rdata(f462_rdata));
  assign f462_clk = clk;
  assign f462_rst = rst;
  // Bindings to f462

  // f464
  logic [0:0] f464_wen;
  logic [31:0] f464_wdata;
  logic [0:0] f464_clk;
  logic [0:0] f464_rst;
  logic [31:0] f464_rdata;
  sr_buffer_32_1 f464(.wen(f464_wen), .wdata(f464_wdata), .clk(f464_clk), .rst(f464_rst), .rdata(f464_rdata));
  assign f464_clk = clk;
  assign f464_rst = rst;
  // Bindings to f464

  // f466
  logic [0:0] f466_wen;
  logic [31:0] f466_wdata;
  logic [0:0] f466_clk;
  logic [0:0] f466_rst;
  logic [31:0] f466_rdata;
  sr_buffer_32_1 f466(.wen(f466_wen), .wdata(f466_wdata), .clk(f466_clk), .rst(f466_rst), .rdata(f466_rdata));
  assign f466_clk = clk;
  assign f466_rst = rst;
  // Bindings to f466

  // f468
  logic [0:0] f468_wen;
  logic [31:0] f468_wdata;
  logic [0:0] f468_clk;
  logic [0:0] f468_rst;
  logic [31:0] f468_rdata;
  sr_buffer_32_1 f468(.wen(f468_wen), .wdata(f468_wdata), .clk(f468_clk), .rst(f468_rst), .rdata(f468_rdata));
  assign f468_clk = clk;
  assign f468_rst = rst;
  // Bindings to f468

  // f470
  logic [0:0] f470_wen;
  logic [31:0] f470_wdata;
  logic [0:0] f470_clk;
  logic [0:0] f470_rst;
  logic [31:0] f470_rdata;
  sr_buffer_32_1 f470(.wen(f470_wen), .wdata(f470_wdata), .clk(f470_clk), .rst(f470_rst), .rdata(f470_rdata));
  assign f470_clk = clk;
  assign f470_rst = rst;
  // Bindings to f470

  // f472
  logic [0:0] f472_wen;
  logic [31:0] f472_wdata;
  logic [0:0] f472_clk;
  logic [0:0] f472_rst;
  logic [31:0] f472_rdata;
  sr_buffer_32_1 f472(.wen(f472_wen), .wdata(f472_wdata), .clk(f472_clk), .rst(f472_rst), .rdata(f472_rdata));
  assign f472_clk = clk;
  assign f472_rst = rst;
  // Bindings to f472

  // f474
  logic [0:0] f474_wen;
  logic [31:0] f474_wdata;
  logic [0:0] f474_clk;
  logic [0:0] f474_rst;
  logic [31:0] f474_rdata;
  sr_buffer_32_1 f474(.wen(f474_wen), .wdata(f474_wdata), .clk(f474_clk), .rst(f474_rst), .rdata(f474_rdata));
  assign f474_clk = clk;
  assign f474_rst = rst;
  // Bindings to f474

  // f476
  logic [0:0] f476_wen;
  logic [31:0] f476_wdata;
  logic [0:0] f476_clk;
  logic [0:0] f476_rst;
  logic [31:0] f476_rdata;
  sr_buffer_32_1 f476(.wen(f476_wen), .wdata(f476_wdata), .clk(f476_clk), .rst(f476_rst), .rdata(f476_rdata));
  assign f476_clk = clk;
  assign f476_rst = rst;
  // Bindings to f476

  // f478
  logic [0:0] f478_wen;
  logic [31:0] f478_wdata;
  logic [0:0] f478_clk;
  logic [0:0] f478_rst;
  logic [31:0] f478_rdata;
  sr_buffer_32_1 f478(.wen(f478_wen), .wdata(f478_wdata), .clk(f478_clk), .rst(f478_rst), .rdata(f478_rdata));
  assign f478_clk = clk;
  assign f478_rst = rst;
  // Bindings to f478

  // f480
  logic [0:0] f480_wen;
  logic [31:0] f480_wdata;
  logic [0:0] f480_clk;
  logic [0:0] f480_rst;
  logic [31:0] f480_rdata;
  sr_buffer_32_1 f480(.wen(f480_wen), .wdata(f480_wdata), .clk(f480_clk), .rst(f480_rst), .rdata(f480_rdata));
  assign f480_clk = clk;
  assign f480_rst = rst;
  // Bindings to f480

  // f482
  logic [0:0] f482_wen;
  logic [31:0] f482_wdata;
  logic [0:0] f482_clk;
  logic [0:0] f482_rst;
  logic [31:0] f482_rdata;
  sr_buffer_32_1 f482(.wen(f482_wen), .wdata(f482_wdata), .clk(f482_clk), .rst(f482_rst), .rdata(f482_rdata));
  assign f482_clk = clk;
  assign f482_rst = rst;
  // Bindings to f482

  // f484
  logic [0:0] f484_wen;
  logic [31:0] f484_wdata;
  logic [0:0] f484_clk;
  logic [0:0] f484_rst;
  logic [31:0] f484_rdata;
  sr_buffer_32_1 f484(.wen(f484_wen), .wdata(f484_wdata), .clk(f484_clk), .rst(f484_rst), .rdata(f484_rdata));
  assign f484_clk = clk;
  assign f484_rst = rst;
  // Bindings to f484

  // f486
  logic [0:0] f486_wen;
  logic [31:0] f486_wdata;
  logic [0:0] f486_clk;
  logic [0:0] f486_rst;
  logic [31:0] f486_rdata;
  sr_buffer_32_1 f486(.wen(f486_wen), .wdata(f486_wdata), .clk(f486_clk), .rst(f486_rst), .rdata(f486_rdata));
  assign f486_clk = clk;
  assign f486_rst = rst;
  // Bindings to f486

  // f488
  logic [0:0] f488_wen;
  logic [31:0] f488_wdata;
  logic [0:0] f488_clk;
  logic [0:0] f488_rst;
  logic [31:0] f488_rdata;
  sr_buffer_32_1 f488(.wen(f488_wen), .wdata(f488_wdata), .clk(f488_clk), .rst(f488_rst), .rdata(f488_rdata));
  assign f488_clk = clk;
  assign f488_rst = rst;
  // Bindings to f488

  // f490
  logic [0:0] f490_wen;
  logic [31:0] f490_wdata;
  logic [0:0] f490_clk;
  logic [0:0] f490_rst;
  logic [31:0] f490_rdata;
  sr_buffer_32_1 f490(.wen(f490_wen), .wdata(f490_wdata), .clk(f490_clk), .rst(f490_rst), .rdata(f490_rdata));
  assign f490_clk = clk;
  assign f490_rst = rst;
  // Bindings to f490

  // f492
  logic [0:0] f492_wen;
  logic [31:0] f492_wdata;
  logic [0:0] f492_clk;
  logic [0:0] f492_rst;
  logic [31:0] f492_rdata;
  sr_buffer_32_1 f492(.wen(f492_wen), .wdata(f492_wdata), .clk(f492_clk), .rst(f492_rst), .rdata(f492_rdata));
  assign f492_clk = clk;
  assign f492_rst = rst;
  // Bindings to f492

  // f494
  logic [0:0] f494_wen;
  logic [31:0] f494_wdata;
  logic [0:0] f494_clk;
  logic [0:0] f494_rst;
  logic [31:0] f494_rdata;
  sr_buffer_32_1 f494(.wen(f494_wen), .wdata(f494_wdata), .clk(f494_clk), .rst(f494_rst), .rdata(f494_rdata));
  assign f494_clk = clk;
  assign f494_rst = rst;
  // Bindings to f494

  // f496
  logic [0:0] f496_wen;
  logic [31:0] f496_wdata;
  logic [0:0] f496_clk;
  logic [0:0] f496_rst;
  logic [31:0] f496_rdata;
  sr_buffer_32_1 f496(.wen(f496_wen), .wdata(f496_wdata), .clk(f496_clk), .rst(f496_rst), .rdata(f496_rdata));
  assign f496_clk = clk;
  assign f496_rst = rst;
  // Bindings to f496

  // f498
  logic [0:0] f498_wen;
  logic [31:0] f498_wdata;
  logic [0:0] f498_clk;
  logic [0:0] f498_rst;
  logic [31:0] f498_rdata;
  sr_buffer_32_1 f498(.wen(f498_wen), .wdata(f498_wdata), .clk(f498_clk), .rst(f498_rst), .rdata(f498_rdata));
  assign f498_clk = clk;
  assign f498_rst = rst;
  // Bindings to f498

  // f500
  logic [0:0] f500_wen;
  logic [31:0] f500_wdata;
  logic [0:0] f500_clk;
  logic [0:0] f500_rst;
  logic [31:0] f500_rdata;
  sr_buffer_32_1 f500(.wen(f500_wen), .wdata(f500_wdata), .clk(f500_clk), .rst(f500_rst), .rdata(f500_rdata));
  assign f500_clk = clk;
  assign f500_rst = rst;
  // Bindings to f500

  // f502
  logic [0:0] f502_wen;
  logic [31:0] f502_wdata;
  logic [0:0] f502_clk;
  logic [0:0] f502_rst;
  logic [31:0] f502_rdata;
  sr_buffer_32_1 f502(.wen(f502_wen), .wdata(f502_wdata), .clk(f502_clk), .rst(f502_rst), .rdata(f502_rdata));
  assign f502_clk = clk;
  assign f502_rst = rst;
  // Bindings to f502

  // f504
  logic [0:0] f504_wen;
  logic [31:0] f504_wdata;
  logic [0:0] f504_clk;
  logic [0:0] f504_rst;
  logic [31:0] f504_rdata;
  sr_buffer_32_1 f504(.wen(f504_wen), .wdata(f504_wdata), .clk(f504_clk), .rst(f504_rst), .rdata(f504_rdata));
  assign f504_clk = clk;
  assign f504_rst = rst;
  // Bindings to f504

  // f506
  logic [0:0] f506_wen;
  logic [31:0] f506_wdata;
  logic [0:0] f506_clk;
  logic [0:0] f506_rst;
  logic [31:0] f506_rdata;
  sr_buffer_32_1 f506(.wen(f506_wen), .wdata(f506_wdata), .clk(f506_clk), .rst(f506_rst), .rdata(f506_rdata));
  assign f506_clk = clk;
  assign f506_rst = rst;
  // Bindings to f506

  // f508
  logic [0:0] f508_wen;
  logic [31:0] f508_wdata;
  logic [0:0] f508_clk;
  logic [0:0] f508_rst;
  logic [31:0] f508_rdata;
  sr_buffer_32_1 f508(.wen(f508_wen), .wdata(f508_wdata), .clk(f508_clk), .rst(f508_rst), .rdata(f508_rdata));
  assign f508_clk = clk;
  assign f508_rst = rst;
  // Bindings to f508

  // f510
  logic [0:0] f510_wen;
  logic [31:0] f510_wdata;
  logic [0:0] f510_clk;
  logic [0:0] f510_rst;
  logic [31:0] f510_rdata;
  sr_buffer_32_1 f510(.wen(f510_wen), .wdata(f510_wdata), .clk(f510_clk), .rst(f510_rst), .rdata(f510_rdata));
  assign f510_clk = clk;
  assign f510_rst = rst;
  // Bindings to f510

  // f512
  logic [0:0] f512_wen;
  logic [31:0] f512_wdata;
  logic [0:0] f512_clk;
  logic [0:0] f512_rst;
  logic [31:0] f512_rdata;
  sr_buffer_32_1 f512(.wen(f512_wen), .wdata(f512_wdata), .clk(f512_clk), .rst(f512_rst), .rdata(f512_rdata));
  assign f512_clk = clk;
  assign f512_rst = rst;
  // Bindings to f512

  // f514
  logic [0:0] f514_wen;
  logic [31:0] f514_wdata;
  logic [0:0] f514_clk;
  logic [0:0] f514_rst;
  logic [31:0] f514_rdata;
  sr_buffer_32_1 f514(.wen(f514_wen), .wdata(f514_wdata), .clk(f514_clk), .rst(f514_rst), .rdata(f514_rdata));
  assign f514_clk = clk;
  assign f514_rst = rst;
  // Bindings to f514

  // f516
  logic [0:0] f516_wen;
  logic [31:0] f516_wdata;
  logic [0:0] f516_clk;
  logic [0:0] f516_rst;
  logic [31:0] f516_rdata;
  sr_buffer_32_1 f516(.wen(f516_wen), .wdata(f516_wdata), .clk(f516_clk), .rst(f516_rst), .rdata(f516_rdata));
  assign f516_clk = clk;
  assign f516_rst = rst;
  // Bindings to f516

  // f518
  logic [0:0] f518_wen;
  logic [31:0] f518_wdata;
  logic [0:0] f518_clk;
  logic [0:0] f518_rst;
  logic [31:0] f518_rdata;
  sr_buffer_32_1 f518(.wen(f518_wen), .wdata(f518_wdata), .clk(f518_clk), .rst(f518_rst), .rdata(f518_rdata));
  assign f518_clk = clk;
  assign f518_rst = rst;
  // Bindings to f518

  // f520
  logic [0:0] f520_wen;
  logic [31:0] f520_wdata;
  logic [0:0] f520_clk;
  logic [0:0] f520_rst;
  logic [31:0] f520_rdata;
  sr_buffer_32_1 f520(.wen(f520_wen), .wdata(f520_wdata), .clk(f520_clk), .rst(f520_rst), .rdata(f520_rdata));
  assign f520_clk = clk;
  assign f520_rst = rst;
  // Bindings to f520

  // f522
  logic [0:0] f522_wen;
  logic [31:0] f522_wdata;
  logic [0:0] f522_clk;
  logic [0:0] f522_rst;
  logic [31:0] f522_rdata;
  sr_buffer_32_1 f522(.wen(f522_wen), .wdata(f522_wdata), .clk(f522_clk), .rst(f522_rst), .rdata(f522_rdata));
  assign f522_clk = clk;
  assign f522_rst = rst;
  // Bindings to f522

  // f524
  logic [0:0] f524_wen;
  logic [31:0] f524_wdata;
  logic [0:0] f524_clk;
  logic [0:0] f524_rst;
  logic [31:0] f524_rdata;
  sr_buffer_32_1 f524(.wen(f524_wen), .wdata(f524_wdata), .clk(f524_clk), .rst(f524_rst), .rdata(f524_rdata));
  assign f524_clk = clk;
  assign f524_rst = rst;
  // Bindings to f524

  // f526
  logic [0:0] f526_wen;
  logic [31:0] f526_wdata;
  logic [0:0] f526_clk;
  logic [0:0] f526_rst;
  logic [31:0] f526_rdata;
  sr_buffer_32_1 f526(.wen(f526_wen), .wdata(f526_wdata), .clk(f526_clk), .rst(f526_rst), .rdata(f526_rdata));
  assign f526_clk = clk;
  assign f526_rst = rst;
  // Bindings to f526

  // f528
  logic [0:0] f528_wen;
  logic [31:0] f528_wdata;
  logic [0:0] f528_clk;
  logic [0:0] f528_rst;
  logic [31:0] f528_rdata;
  sr_buffer_32_1 f528(.wen(f528_wen), .wdata(f528_wdata), .clk(f528_clk), .rst(f528_rst), .rdata(f528_rdata));
  assign f528_clk = clk;
  assign f528_rst = rst;
  // Bindings to f528

  // f530
  logic [0:0] f530_wen;
  logic [31:0] f530_wdata;
  logic [0:0] f530_clk;
  logic [0:0] f530_rst;
  logic [31:0] f530_rdata;
  sr_buffer_32_1 f530(.wen(f530_wen), .wdata(f530_wdata), .clk(f530_clk), .rst(f530_rst), .rdata(f530_rdata));
  assign f530_clk = clk;
  assign f530_rst = rst;
  // Bindings to f530

  // f532
  logic [0:0] f532_wen;
  logic [31:0] f532_wdata;
  logic [0:0] f532_clk;
  logic [0:0] f532_rst;
  logic [31:0] f532_rdata;
  sr_buffer_32_1 f532(.wen(f532_wen), .wdata(f532_wdata), .clk(f532_clk), .rst(f532_rst), .rdata(f532_rdata));
  assign f532_clk = clk;
  assign f532_rst = rst;
  // Bindings to f532

  // f534
  logic [0:0] f534_wen;
  logic [31:0] f534_wdata;
  logic [0:0] f534_clk;
  logic [0:0] f534_rst;
  logic [31:0] f534_rdata;
  sr_buffer_32_1 f534(.wen(f534_wen), .wdata(f534_wdata), .clk(f534_clk), .rst(f534_rst), .rdata(f534_rdata));
  assign f534_clk = clk;
  assign f534_rst = rst;
  // Bindings to f534

  // f536
  logic [0:0] f536_wen;
  logic [31:0] f536_wdata;
  logic [0:0] f536_clk;
  logic [0:0] f536_rst;
  logic [31:0] f536_rdata;
  sr_buffer_32_1 f536(.wen(f536_wen), .wdata(f536_wdata), .clk(f536_clk), .rst(f536_rst), .rdata(f536_rdata));
  assign f536_clk = clk;
  assign f536_rst = rst;
  // Bindings to f536

  // f538
  logic [0:0] f538_wen;
  logic [31:0] f538_wdata;
  logic [0:0] f538_clk;
  logic [0:0] f538_rst;
  logic [31:0] f538_rdata;
  sr_buffer_32_1 f538(.wen(f538_wen), .wdata(f538_wdata), .clk(f538_clk), .rst(f538_rst), .rdata(f538_rdata));
  assign f538_clk = clk;
  assign f538_rst = rst;
  // Bindings to f538

  // f540
  logic [0:0] f540_wen;
  logic [31:0] f540_wdata;
  logic [0:0] f540_clk;
  logic [0:0] f540_rst;
  logic [31:0] f540_rdata;
  sr_buffer_32_1 f540(.wen(f540_wen), .wdata(f540_wdata), .clk(f540_clk), .rst(f540_rst), .rdata(f540_rdata));
  assign f540_clk = clk;
  assign f540_rst = rst;
  // Bindings to f540

  // f542
  logic [0:0] f542_wen;
  logic [31:0] f542_wdata;
  logic [0:0] f542_clk;
  logic [0:0] f542_rst;
  logic [31:0] f542_rdata;
  sr_buffer_32_1 f542(.wen(f542_wen), .wdata(f542_wdata), .clk(f542_clk), .rst(f542_rst), .rdata(f542_rdata));
  assign f542_clk = clk;
  assign f542_rst = rst;
  // Bindings to f542

  // f544
  logic [0:0] f544_wen;
  logic [31:0] f544_wdata;
  logic [0:0] f544_clk;
  logic [0:0] f544_rst;
  logic [31:0] f544_rdata;
  sr_buffer_32_1 f544(.wen(f544_wen), .wdata(f544_wdata), .clk(f544_clk), .rst(f544_rst), .rdata(f544_rdata));
  assign f544_clk = clk;
  assign f544_rst = rst;
  // Bindings to f544

  // f546
  logic [0:0] f546_wen;
  logic [31:0] f546_wdata;
  logic [0:0] f546_clk;
  logic [0:0] f546_rst;
  logic [31:0] f546_rdata;
  sr_buffer_32_1 f546(.wen(f546_wen), .wdata(f546_wdata), .clk(f546_clk), .rst(f546_rst), .rdata(f546_rdata));
  assign f546_clk = clk;
  assign f546_rst = rst;
  // Bindings to f546

  // f548
  logic [0:0] f548_wen;
  logic [31:0] f548_wdata;
  logic [0:0] f548_clk;
  logic [0:0] f548_rst;
  logic [31:0] f548_rdata;
  sr_buffer_32_1 f548(.wen(f548_wen), .wdata(f548_wdata), .clk(f548_clk), .rst(f548_rst), .rdata(f548_rdata));
  assign f548_clk = clk;
  assign f548_rst = rst;
  // Bindings to f548

  // f550
  logic [0:0] f550_wen;
  logic [31:0] f550_wdata;
  logic [0:0] f550_clk;
  logic [0:0] f550_rst;
  logic [31:0] f550_rdata;
  sr_buffer_32_1 f550(.wen(f550_wen), .wdata(f550_wdata), .clk(f550_clk), .rst(f550_rst), .rdata(f550_rdata));
  assign f550_clk = clk;
  assign f550_rst = rst;
  // Bindings to f550

  // f552
  logic [0:0] f552_wen;
  logic [31:0] f552_wdata;
  logic [0:0] f552_clk;
  logic [0:0] f552_rst;
  logic [31:0] f552_rdata;
  sr_buffer_32_1 f552(.wen(f552_wen), .wdata(f552_wdata), .clk(f552_clk), .rst(f552_rst), .rdata(f552_rdata));
  assign f552_clk = clk;
  assign f552_rst = rst;
  // Bindings to f552

  // f554
  logic [0:0] f554_wen;
  logic [31:0] f554_wdata;
  logic [0:0] f554_clk;
  logic [0:0] f554_rst;
  logic [31:0] f554_rdata;
  sr_buffer_32_1 f554(.wen(f554_wen), .wdata(f554_wdata), .clk(f554_clk), .rst(f554_rst), .rdata(f554_rdata));
  assign f554_clk = clk;
  assign f554_rst = rst;
  // Bindings to f554

  // f556
  logic [0:0] f556_wen;
  logic [31:0] f556_wdata;
  logic [0:0] f556_clk;
  logic [0:0] f556_rst;
  logic [31:0] f556_rdata;
  sr_buffer_32_1 f556(.wen(f556_wen), .wdata(f556_wdata), .clk(f556_clk), .rst(f556_rst), .rdata(f556_rdata));
  assign f556_clk = clk;
  assign f556_rst = rst;
  // Bindings to f556

  // f558
  logic [0:0] f558_wen;
  logic [31:0] f558_wdata;
  logic [0:0] f558_clk;
  logic [0:0] f558_rst;
  logic [31:0] f558_rdata;
  sr_buffer_32_1 f558(.wen(f558_wen), .wdata(f558_wdata), .clk(f558_clk), .rst(f558_rst), .rdata(f558_rdata));
  assign f558_clk = clk;
  assign f558_rst = rst;
  // Bindings to f558

  // f560
  logic [0:0] f560_wen;
  logic [31:0] f560_wdata;
  logic [0:0] f560_clk;
  logic [0:0] f560_rst;
  logic [31:0] f560_rdata;
  sr_buffer_32_1 f560(.wen(f560_wen), .wdata(f560_wdata), .clk(f560_clk), .rst(f560_rst), .rdata(f560_rdata));
  assign f560_clk = clk;
  assign f560_rst = rst;
  // Bindings to f560

  // f562
  logic [0:0] f562_wen;
  logic [31:0] f562_wdata;
  logic [0:0] f562_clk;
  logic [0:0] f562_rst;
  logic [31:0] f562_rdata;
  sr_buffer_32_1 f562(.wen(f562_wen), .wdata(f562_wdata), .clk(f562_clk), .rst(f562_rst), .rdata(f562_rdata));
  assign f562_clk = clk;
  assign f562_rst = rst;
  // Bindings to f562

  // f564
  logic [0:0] f564_wen;
  logic [31:0] f564_wdata;
  logic [0:0] f564_clk;
  logic [0:0] f564_rst;
  logic [31:0] f564_rdata;
  sr_buffer_32_1 f564(.wen(f564_wen), .wdata(f564_wdata), .clk(f564_clk), .rst(f564_rst), .rdata(f564_rdata));
  assign f564_clk = clk;
  assign f564_rst = rst;
  // Bindings to f564

  // f566
  logic [0:0] f566_wen;
  logic [31:0] f566_wdata;
  logic [0:0] f566_clk;
  logic [0:0] f566_rst;
  logic [31:0] f566_rdata;
  sr_buffer_32_1 f566(.wen(f566_wen), .wdata(f566_wdata), .clk(f566_clk), .rst(f566_rst), .rdata(f566_rdata));
  assign f566_clk = clk;
  assign f566_rst = rst;
  // Bindings to f566

  // f568
  logic [0:0] f568_wen;
  logic [31:0] f568_wdata;
  logic [0:0] f568_clk;
  logic [0:0] f568_rst;
  logic [31:0] f568_rdata;
  sr_buffer_32_1 f568(.wen(f568_wen), .wdata(f568_wdata), .clk(f568_clk), .rst(f568_rst), .rdata(f568_rdata));
  assign f568_clk = clk;
  assign f568_rst = rst;
  // Bindings to f568

  // f570
  logic [0:0] f570_wen;
  logic [31:0] f570_wdata;
  logic [0:0] f570_clk;
  logic [0:0] f570_rst;
  logic [31:0] f570_rdata;
  sr_buffer_32_1 f570(.wen(f570_wen), .wdata(f570_wdata), .clk(f570_clk), .rst(f570_rst), .rdata(f570_rdata));
  assign f570_clk = clk;
  assign f570_rst = rst;
  // Bindings to f570

  // f572
  logic [0:0] f572_wen;
  logic [31:0] f572_wdata;
  logic [0:0] f572_clk;
  logic [0:0] f572_rst;
  logic [31:0] f572_rdata;
  sr_buffer_32_1 f572(.wen(f572_wen), .wdata(f572_wdata), .clk(f572_clk), .rst(f572_rst), .rdata(f572_rdata));
  assign f572_clk = clk;
  assign f572_rst = rst;
  // Bindings to f572

  // f574
  logic [0:0] f574_wen;
  logic [31:0] f574_wdata;
  logic [0:0] f574_clk;
  logic [0:0] f574_rst;
  logic [31:0] f574_rdata;
  sr_buffer_32_1 f574(.wen(f574_wen), .wdata(f574_wdata), .clk(f574_clk), .rst(f574_rst), .rdata(f574_rdata));
  assign f574_clk = clk;
  assign f574_rst = rst;
  // Bindings to f574

  // f576
  logic [0:0] f576_wen;
  logic [31:0] f576_wdata;
  logic [0:0] f576_clk;
  logic [0:0] f576_rst;
  logic [31:0] f576_rdata;
  sr_buffer_32_1 f576(.wen(f576_wen), .wdata(f576_wdata), .clk(f576_clk), .rst(f576_rst), .rdata(f576_rdata));
  assign f576_clk = clk;
  assign f576_rst = rst;
  // Bindings to f576

  // f578
  logic [0:0] f578_wen;
  logic [31:0] f578_wdata;
  logic [0:0] f578_clk;
  logic [0:0] f578_rst;
  logic [31:0] f578_rdata;
  sr_buffer_32_1 f578(.wen(f578_wen), .wdata(f578_wdata), .clk(f578_clk), .rst(f578_rst), .rdata(f578_rdata));
  assign f578_clk = clk;
  assign f578_rst = rst;
  // Bindings to f578

  // f580
  logic [0:0] f580_wen;
  logic [31:0] f580_wdata;
  logic [0:0] f580_clk;
  logic [0:0] f580_rst;
  logic [31:0] f580_rdata;
  sr_buffer_32_1 f580(.wen(f580_wen), .wdata(f580_wdata), .clk(f580_clk), .rst(f580_rst), .rdata(f580_rdata));
  assign f580_clk = clk;
  assign f580_rst = rst;
  // Bindings to f580

  // f582
  logic [0:0] f582_wen;
  logic [31:0] f582_wdata;
  logic [0:0] f582_clk;
  logic [0:0] f582_rst;
  logic [31:0] f582_rdata;
  sr_buffer_32_1 f582(.wen(f582_wen), .wdata(f582_wdata), .clk(f582_clk), .rst(f582_rst), .rdata(f582_rdata));
  assign f582_clk = clk;
  assign f582_rst = rst;
  // Bindings to f582

  // f584
  logic [0:0] f584_wen;
  logic [31:0] f584_wdata;
  logic [0:0] f584_clk;
  logic [0:0] f584_rst;
  logic [31:0] f584_rdata;
  sr_buffer_32_1 f584(.wen(f584_wen), .wdata(f584_wdata), .clk(f584_clk), .rst(f584_rst), .rdata(f584_rdata));
  assign f584_clk = clk;
  assign f584_rst = rst;
  // Bindings to f584

  // f586
  logic [0:0] f586_wen;
  logic [31:0] f586_wdata;
  logic [0:0] f586_clk;
  logic [0:0] f586_rst;
  logic [31:0] f586_rdata;
  sr_buffer_32_1 f586(.wen(f586_wen), .wdata(f586_wdata), .clk(f586_clk), .rst(f586_rst), .rdata(f586_rdata));
  assign f586_clk = clk;
  assign f586_rst = rst;
  // Bindings to f586

  // f588
  logic [0:0] f588_wen;
  logic [31:0] f588_wdata;
  logic [0:0] f588_clk;
  logic [0:0] f588_rst;
  logic [31:0] f588_rdata;
  sr_buffer_32_1 f588(.wen(f588_wen), .wdata(f588_wdata), .clk(f588_clk), .rst(f588_rst), .rdata(f588_rdata));
  assign f588_clk = clk;
  assign f588_rst = rst;
  // Bindings to f588

  // f590
  logic [0:0] f590_wen;
  logic [31:0] f590_wdata;
  logic [0:0] f590_clk;
  logic [0:0] f590_rst;
  logic [31:0] f590_rdata;
  sr_buffer_32_1 f590(.wen(f590_wen), .wdata(f590_wdata), .clk(f590_clk), .rst(f590_rst), .rdata(f590_rdata));
  assign f590_clk = clk;
  assign f590_rst = rst;
  // Bindings to f590

  // f592
  logic [0:0] f592_wen;
  logic [31:0] f592_wdata;
  logic [0:0] f592_clk;
  logic [0:0] f592_rst;
  logic [31:0] f592_rdata;
  sr_buffer_32_1 f592(.wen(f592_wen), .wdata(f592_wdata), .clk(f592_clk), .rst(f592_rst), .rdata(f592_rdata));
  assign f592_clk = clk;
  assign f592_rst = rst;
  // Bindings to f592

  // f594
  logic [0:0] f594_wen;
  logic [31:0] f594_wdata;
  logic [0:0] f594_clk;
  logic [0:0] f594_rst;
  logic [31:0] f594_rdata;
  sr_buffer_32_1 f594(.wen(f594_wen), .wdata(f594_wdata), .clk(f594_clk), .rst(f594_rst), .rdata(f594_rdata));
  assign f594_clk = clk;
  assign f594_rst = rst;
  // Bindings to f594

  // f596
  logic [0:0] f596_wen;
  logic [31:0] f596_wdata;
  logic [0:0] f596_clk;
  logic [0:0] f596_rst;
  logic [31:0] f596_rdata;
  sr_buffer_32_1 f596(.wen(f596_wen), .wdata(f596_wdata), .clk(f596_clk), .rst(f596_rst), .rdata(f596_rdata));
  assign f596_clk = clk;
  assign f596_rst = rst;
  // Bindings to f596

  // f598
  logic [0:0] f598_wen;
  logic [31:0] f598_wdata;
  logic [0:0] f598_clk;
  logic [0:0] f598_rst;
  logic [31:0] f598_rdata;
  sr_buffer_32_1 f598(.wen(f598_wen), .wdata(f598_wdata), .clk(f598_clk), .rst(f598_rst), .rdata(f598_rdata));
  assign f598_clk = clk;
  assign f598_rst = rst;
  // Bindings to f598

  // f600
  logic [0:0] f600_wen;
  logic [31:0] f600_wdata;
  logic [0:0] f600_clk;
  logic [0:0] f600_rst;
  logic [31:0] f600_rdata;
  sr_buffer_32_1 f600(.wen(f600_wen), .wdata(f600_wdata), .clk(f600_clk), .rst(f600_rst), .rdata(f600_rdata));
  assign f600_clk = clk;
  assign f600_rst = rst;
  // Bindings to f600

  // f602
  logic [0:0] f602_wen;
  logic [31:0] f602_wdata;
  logic [0:0] f602_clk;
  logic [0:0] f602_rst;
  logic [31:0] f602_rdata;
  sr_buffer_32_1 f602(.wen(f602_wen), .wdata(f602_wdata), .clk(f602_clk), .rst(f602_rst), .rdata(f602_rdata));
  assign f602_clk = clk;
  assign f602_rst = rst;
  // Bindings to f602

  // f604
  logic [0:0] f604_wen;
  logic [31:0] f604_wdata;
  logic [0:0] f604_clk;
  logic [0:0] f604_rst;
  logic [31:0] f604_rdata;
  sr_buffer_32_1 f604(.wen(f604_wen), .wdata(f604_wdata), .clk(f604_clk), .rst(f604_rst), .rdata(f604_rdata));
  assign f604_clk = clk;
  assign f604_rst = rst;
  // Bindings to f604

  // f606
  logic [0:0] f606_wen;
  logic [31:0] f606_wdata;
  logic [0:0] f606_clk;
  logic [0:0] f606_rst;
  logic [31:0] f606_rdata;
  sr_buffer_32_1 f606(.wen(f606_wen), .wdata(f606_wdata), .clk(f606_clk), .rst(f606_rst), .rdata(f606_rdata));
  assign f606_clk = clk;
  assign f606_rst = rst;
  // Bindings to f606

  // f608
  logic [0:0] f608_wen;
  logic [31:0] f608_wdata;
  logic [0:0] f608_clk;
  logic [0:0] f608_rst;
  logic [31:0] f608_rdata;
  sr_buffer_32_1 f608(.wen(f608_wen), .wdata(f608_wdata), .clk(f608_clk), .rst(f608_rst), .rdata(f608_rdata));
  assign f608_clk = clk;
  assign f608_rst = rst;
  // Bindings to f608

  // f610
  logic [0:0] f610_wen;
  logic [31:0] f610_wdata;
  logic [0:0] f610_clk;
  logic [0:0] f610_rst;
  logic [31:0] f610_rdata;
  sr_buffer_32_1 f610(.wen(f610_wen), .wdata(f610_wdata), .clk(f610_clk), .rst(f610_rst), .rdata(f610_rdata));
  assign f610_clk = clk;
  assign f610_rst = rst;
  // Bindings to f610

  // f612
  logic [0:0] f612_wen;
  logic [31:0] f612_wdata;
  logic [0:0] f612_clk;
  logic [0:0] f612_rst;
  logic [31:0] f612_rdata;
  sr_buffer_32_1 f612(.wen(f612_wen), .wdata(f612_wdata), .clk(f612_clk), .rst(f612_rst), .rdata(f612_rdata));
  assign f612_clk = clk;
  assign f612_rst = rst;
  // Bindings to f612

  // f614
  logic [0:0] f614_wen;
  logic [31:0] f614_wdata;
  logic [0:0] f614_clk;
  logic [0:0] f614_rst;
  logic [31:0] f614_rdata;
  sr_buffer_32_1 f614(.wen(f614_wen), .wdata(f614_wdata), .clk(f614_clk), .rst(f614_rst), .rdata(f614_rdata));
  assign f614_clk = clk;
  assign f614_rst = rst;
  // Bindings to f614

  // f616
  logic [0:0] f616_wen;
  logic [31:0] f616_wdata;
  logic [0:0] f616_clk;
  logic [0:0] f616_rst;
  logic [31:0] f616_rdata;
  sr_buffer_32_1 f616(.wen(f616_wen), .wdata(f616_wdata), .clk(f616_clk), .rst(f616_rst), .rdata(f616_rdata));
  assign f616_clk = clk;
  assign f616_rst = rst;
  // Bindings to f616

  // f618
  logic [0:0] f618_wen;
  logic [31:0] f618_wdata;
  logic [0:0] f618_clk;
  logic [0:0] f618_rst;
  logic [31:0] f618_rdata;
  sr_buffer_32_1 f618(.wen(f618_wen), .wdata(f618_wdata), .clk(f618_clk), .rst(f618_rst), .rdata(f618_rdata));
  assign f618_clk = clk;
  assign f618_rst = rst;
  // Bindings to f618

  // f620
  logic [0:0] f620_wen;
  logic [31:0] f620_wdata;
  logic [0:0] f620_clk;
  logic [0:0] f620_rst;
  logic [31:0] f620_rdata;
  sr_buffer_32_1 f620(.wen(f620_wen), .wdata(f620_wdata), .clk(f620_clk), .rst(f620_rst), .rdata(f620_rdata));
  assign f620_clk = clk;
  assign f620_rst = rst;
  // Bindings to f620

  // f622
  logic [0:0] f622_wen;
  logic [31:0] f622_wdata;
  logic [0:0] f622_clk;
  logic [0:0] f622_rst;
  logic [31:0] f622_rdata;
  sr_buffer_32_1 f622(.wen(f622_wen), .wdata(f622_wdata), .clk(f622_clk), .rst(f622_rst), .rdata(f622_rdata));
  assign f622_clk = clk;
  assign f622_rst = rst;
  // Bindings to f622

  // f624
  logic [0:0] f624_wen;
  logic [31:0] f624_wdata;
  logic [0:0] f624_clk;
  logic [0:0] f624_rst;
  logic [31:0] f624_rdata;
  sr_buffer_32_1 f624(.wen(f624_wen), .wdata(f624_wdata), .clk(f624_clk), .rst(f624_rst), .rdata(f624_rdata));
  assign f624_clk = clk;
  assign f624_rst = rst;
  // Bindings to f624

  // f626
  logic [0:0] f626_wen;
  logic [31:0] f626_wdata;
  logic [0:0] f626_clk;
  logic [0:0] f626_rst;
  logic [31:0] f626_rdata;
  sr_buffer_32_1 f626(.wen(f626_wen), .wdata(f626_wdata), .clk(f626_clk), .rst(f626_rst), .rdata(f626_rdata));
  assign f626_clk = clk;
  assign f626_rst = rst;
  // Bindings to f626

  // f628
  logic [0:0] f628_wen;
  logic [31:0] f628_wdata;
  logic [0:0] f628_clk;
  logic [0:0] f628_rst;
  logic [31:0] f628_rdata;
  sr_buffer_32_1 f628(.wen(f628_wen), .wdata(f628_wdata), .clk(f628_clk), .rst(f628_rst), .rdata(f628_rdata));
  assign f628_clk = clk;
  assign f628_rst = rst;
  // Bindings to f628

  // f630
  logic [0:0] f630_wen;
  logic [31:0] f630_wdata;
  logic [0:0] f630_clk;
  logic [0:0] f630_rst;
  logic [31:0] f630_rdata;
  sr_buffer_32_1 f630(.wen(f630_wen), .wdata(f630_wdata), .clk(f630_clk), .rst(f630_rst), .rdata(f630_rdata));
  assign f630_clk = clk;
  assign f630_rst = rst;
  // Bindings to f630

  // f632
  logic [0:0] f632_wen;
  logic [31:0] f632_wdata;
  logic [0:0] f632_clk;
  logic [0:0] f632_rst;
  logic [31:0] f632_rdata;
  sr_buffer_32_1 f632(.wen(f632_wen), .wdata(f632_wdata), .clk(f632_clk), .rst(f632_rst), .rdata(f632_rdata));
  assign f632_clk = clk;
  assign f632_rst = rst;
  // Bindings to f632

  // f634
  logic [0:0] f634_wen;
  logic [31:0] f634_wdata;
  logic [0:0] f634_clk;
  logic [0:0] f634_rst;
  logic [31:0] f634_rdata;
  sr_buffer_32_1 f634(.wen(f634_wen), .wdata(f634_wdata), .clk(f634_clk), .rst(f634_rst), .rdata(f634_rdata));
  assign f634_clk = clk;
  assign f634_rst = rst;
  // Bindings to f634

  // f636
  logic [0:0] f636_wen;
  logic [31:0] f636_wdata;
  logic [0:0] f636_clk;
  logic [0:0] f636_rst;
  logic [31:0] f636_rdata;
  sr_buffer_32_1 f636(.wen(f636_wen), .wdata(f636_wdata), .clk(f636_clk), .rst(f636_rst), .rdata(f636_rdata));
  assign f636_clk = clk;
  assign f636_rst = rst;
  // Bindings to f636

  // f638
  logic [0:0] f638_wen;
  logic [31:0] f638_wdata;
  logic [0:0] f638_clk;
  logic [0:0] f638_rst;
  logic [31:0] f638_rdata;
  sr_buffer_32_1 f638(.wen(f638_wen), .wdata(f638_wdata), .clk(f638_clk), .rst(f638_rst), .rdata(f638_rdata));
  assign f638_clk = clk;
  assign f638_rst = rst;
  // Bindings to f638

  // f640
  logic [0:0] f640_wen;
  logic [31:0] f640_wdata;
  logic [0:0] f640_clk;
  logic [0:0] f640_rst;
  logic [31:0] f640_rdata;
  sr_buffer_32_1 f640(.wen(f640_wen), .wdata(f640_wdata), .clk(f640_clk), .rst(f640_rst), .rdata(f640_rdata));
  assign f640_clk = clk;
  assign f640_rst = rst;
  // Bindings to f640

  // f642
  logic [0:0] f642_wen;
  logic [31:0] f642_wdata;
  logic [0:0] f642_clk;
  logic [0:0] f642_rst;
  logic [31:0] f642_rdata;
  sr_buffer_32_1 f642(.wen(f642_wen), .wdata(f642_wdata), .clk(f642_clk), .rst(f642_rst), .rdata(f642_rdata));
  assign f642_clk = clk;
  assign f642_rst = rst;
  // Bindings to f642

  // f644
  logic [0:0] f644_wen;
  logic [31:0] f644_wdata;
  logic [0:0] f644_clk;
  logic [0:0] f644_rst;
  logic [31:0] f644_rdata;
  sr_buffer_32_1 f644(.wen(f644_wen), .wdata(f644_wdata), .clk(f644_clk), .rst(f644_rst), .rdata(f644_rdata));
  assign f644_clk = clk;
  assign f644_rst = rst;
  // Bindings to f644

  // f646
  logic [0:0] f646_wen;
  logic [31:0] f646_wdata;
  logic [0:0] f646_clk;
  logic [0:0] f646_rst;
  logic [31:0] f646_rdata;
  sr_buffer_32_1 f646(.wen(f646_wen), .wdata(f646_wdata), .clk(f646_clk), .rst(f646_rst), .rdata(f646_rdata));
  assign f646_clk = clk;
  assign f646_rst = rst;
  // Bindings to f646

  // f648
  logic [0:0] f648_wen;
  logic [31:0] f648_wdata;
  logic [0:0] f648_clk;
  logic [0:0] f648_rst;
  logic [31:0] f648_rdata;
  sr_buffer_32_1 f648(.wen(f648_wen), .wdata(f648_wdata), .clk(f648_clk), .rst(f648_rst), .rdata(f648_rdata));
  assign f648_clk = clk;
  assign f648_rst = rst;
  // Bindings to f648

  // f650
  logic [0:0] f650_wen;
  logic [31:0] f650_wdata;
  logic [0:0] f650_clk;
  logic [0:0] f650_rst;
  logic [31:0] f650_rdata;
  sr_buffer_32_1 f650(.wen(f650_wen), .wdata(f650_wdata), .clk(f650_clk), .rst(f650_rst), .rdata(f650_rdata));
  assign f650_clk = clk;
  assign f650_rst = rst;
  // Bindings to f650

  // f652
  logic [0:0] f652_wen;
  logic [31:0] f652_wdata;
  logic [0:0] f652_clk;
  logic [0:0] f652_rst;
  logic [31:0] f652_rdata;
  sr_buffer_32_1 f652(.wen(f652_wen), .wdata(f652_wdata), .clk(f652_clk), .rst(f652_rst), .rdata(f652_rdata));
  assign f652_clk = clk;
  assign f652_rst = rst;
  // Bindings to f652

  // f654
  logic [0:0] f654_wen;
  logic [31:0] f654_wdata;
  logic [0:0] f654_clk;
  logic [0:0] f654_rst;
  logic [31:0] f654_rdata;
  sr_buffer_32_1 f654(.wen(f654_wen), .wdata(f654_wdata), .clk(f654_clk), .rst(f654_rst), .rdata(f654_rdata));
  assign f654_clk = clk;
  assign f654_rst = rst;
  // Bindings to f654

  // f656
  logic [0:0] f656_wen;
  logic [31:0] f656_wdata;
  logic [0:0] f656_clk;
  logic [0:0] f656_rst;
  logic [31:0] f656_rdata;
  sr_buffer_32_1 f656(.wen(f656_wen), .wdata(f656_wdata), .clk(f656_clk), .rst(f656_rst), .rdata(f656_rdata));
  assign f656_clk = clk;
  assign f656_rst = rst;
  // Bindings to f656

  // f658
  logic [0:0] f658_wen;
  logic [31:0] f658_wdata;
  logic [0:0] f658_clk;
  logic [0:0] f658_rst;
  logic [31:0] f658_rdata;
  sr_buffer_32_1 f658(.wen(f658_wen), .wdata(f658_wdata), .clk(f658_clk), .rst(f658_rst), .rdata(f658_rdata));
  assign f658_clk = clk;
  assign f658_rst = rst;
  // Bindings to f658

  // f660
  logic [0:0] f660_wen;
  logic [31:0] f660_wdata;
  logic [0:0] f660_clk;
  logic [0:0] f660_rst;
  logic [31:0] f660_rdata;
  sr_buffer_32_1 f660(.wen(f660_wen), .wdata(f660_wdata), .clk(f660_clk), .rst(f660_rst), .rdata(f660_rdata));
  assign f660_clk = clk;
  assign f660_rst = rst;
  // Bindings to f660

  // f662
  logic [0:0] f662_wen;
  logic [31:0] f662_wdata;
  logic [0:0] f662_clk;
  logic [0:0] f662_rst;
  logic [31:0] f662_rdata;
  sr_buffer_32_1 f662(.wen(f662_wen), .wdata(f662_wdata), .clk(f662_clk), .rst(f662_rst), .rdata(f662_rdata));
  assign f662_clk = clk;
  assign f662_rst = rst;
  // Bindings to f662

  // f664
  logic [0:0] f664_wen;
  logic [31:0] f664_wdata;
  logic [0:0] f664_clk;
  logic [0:0] f664_rst;
  logic [31:0] f664_rdata;
  sr_buffer_32_1 f664(.wen(f664_wen), .wdata(f664_wdata), .clk(f664_clk), .rst(f664_rst), .rdata(f664_rdata));
  assign f664_clk = clk;
  assign f664_rst = rst;
  // Bindings to f664

  // f666
  logic [0:0] f666_wen;
  logic [31:0] f666_wdata;
  logic [0:0] f666_clk;
  logic [0:0] f666_rst;
  logic [31:0] f666_rdata;
  sr_buffer_32_1 f666(.wen(f666_wen), .wdata(f666_wdata), .clk(f666_clk), .rst(f666_rst), .rdata(f666_rdata));
  assign f666_clk = clk;
  assign f666_rst = rst;
  // Bindings to f666

  // f668
  logic [0:0] f668_wen;
  logic [31:0] f668_wdata;
  logic [0:0] f668_clk;
  logic [0:0] f668_rst;
  logic [31:0] f668_rdata;
  sr_buffer_32_1 f668(.wen(f668_wen), .wdata(f668_wdata), .clk(f668_clk), .rst(f668_rst), .rdata(f668_rdata));
  assign f668_clk = clk;
  assign f668_rst = rst;
  // Bindings to f668

  // f670
  logic [0:0] f670_wen;
  logic [31:0] f670_wdata;
  logic [0:0] f670_clk;
  logic [0:0] f670_rst;
  logic [31:0] f670_rdata;
  sr_buffer_32_1 f670(.wen(f670_wen), .wdata(f670_wdata), .clk(f670_clk), .rst(f670_rst), .rdata(f670_rdata));
  assign f670_clk = clk;
  assign f670_rst = rst;
  // Bindings to f670

  // f672
  logic [0:0] f672_wen;
  logic [31:0] f672_wdata;
  logic [0:0] f672_clk;
  logic [0:0] f672_rst;
  logic [31:0] f672_rdata;
  sr_buffer_32_1 f672(.wen(f672_wen), .wdata(f672_wdata), .clk(f672_clk), .rst(f672_rst), .rdata(f672_rdata));
  assign f672_clk = clk;
  assign f672_rst = rst;
  // Bindings to f672

  // f674
  logic [0:0] f674_wen;
  logic [31:0] f674_wdata;
  logic [0:0] f674_clk;
  logic [0:0] f674_rst;
  logic [31:0] f674_rdata;
  sr_buffer_32_1 f674(.wen(f674_wen), .wdata(f674_wdata), .clk(f674_clk), .rst(f674_rst), .rdata(f674_rdata));
  assign f674_clk = clk;
  assign f674_rst = rst;
  // Bindings to f674

  // f676
  logic [0:0] f676_wen;
  logic [31:0] f676_wdata;
  logic [0:0] f676_clk;
  logic [0:0] f676_rst;
  logic [31:0] f676_rdata;
  sr_buffer_32_1 f676(.wen(f676_wen), .wdata(f676_wdata), .clk(f676_clk), .rst(f676_rst), .rdata(f676_rdata));
  assign f676_clk = clk;
  assign f676_rst = rst;
  // Bindings to f676

  // f678
  logic [0:0] f678_wen;
  logic [31:0] f678_wdata;
  logic [0:0] f678_clk;
  logic [0:0] f678_rst;
  logic [31:0] f678_rdata;
  sr_buffer_32_1 f678(.wen(f678_wen), .wdata(f678_wdata), .clk(f678_clk), .rst(f678_rst), .rdata(f678_rdata));
  assign f678_clk = clk;
  assign f678_rst = rst;
  // Bindings to f678

  // f680
  logic [0:0] f680_wen;
  logic [31:0] f680_wdata;
  logic [0:0] f680_clk;
  logic [0:0] f680_rst;
  logic [31:0] f680_rdata;
  sr_buffer_32_1 f680(.wen(f680_wen), .wdata(f680_wdata), .clk(f680_clk), .rst(f680_rst), .rdata(f680_rdata));
  assign f680_clk = clk;
  assign f680_rst = rst;
  // Bindings to f680

  // f682
  logic [0:0] f682_wen;
  logic [31:0] f682_wdata;
  logic [0:0] f682_clk;
  logic [0:0] f682_rst;
  logic [31:0] f682_rdata;
  sr_buffer_32_1 f682(.wen(f682_wen), .wdata(f682_wdata), .clk(f682_clk), .rst(f682_rst), .rdata(f682_rdata));
  assign f682_clk = clk;
  assign f682_rst = rst;
  // Bindings to f682

  // f684
  logic [0:0] f684_wen;
  logic [31:0] f684_wdata;
  logic [0:0] f684_clk;
  logic [0:0] f684_rst;
  logic [31:0] f684_rdata;
  sr_buffer_32_1 f684(.wen(f684_wen), .wdata(f684_wdata), .clk(f684_clk), .rst(f684_rst), .rdata(f684_rdata));
  assign f684_clk = clk;
  assign f684_rst = rst;
  // Bindings to f684

  // f686
  logic [0:0] f686_wen;
  logic [31:0] f686_wdata;
  logic [0:0] f686_clk;
  logic [0:0] f686_rst;
  logic [31:0] f686_rdata;
  sr_buffer_32_1 f686(.wen(f686_wen), .wdata(f686_wdata), .clk(f686_clk), .rst(f686_rst), .rdata(f686_rdata));
  assign f686_clk = clk;
  assign f686_rst = rst;
  // Bindings to f686

  // f688
  logic [0:0] f688_wen;
  logic [31:0] f688_wdata;
  logic [0:0] f688_clk;
  logic [0:0] f688_rst;
  logic [31:0] f688_rdata;
  sr_buffer_32_1 f688(.wen(f688_wen), .wdata(f688_wdata), .clk(f688_clk), .rst(f688_rst), .rdata(f688_rdata));
  assign f688_clk = clk;
  assign f688_rst = rst;
  // Bindings to f688

  // f690
  logic [0:0] f690_wen;
  logic [31:0] f690_wdata;
  logic [0:0] f690_clk;
  logic [0:0] f690_rst;
  logic [31:0] f690_rdata;
  sr_buffer_32_1 f690(.wen(f690_wen), .wdata(f690_wdata), .clk(f690_clk), .rst(f690_rst), .rdata(f690_rdata));
  assign f690_clk = clk;
  assign f690_rst = rst;
  // Bindings to f690

  // f692
  logic [0:0] f692_wen;
  logic [31:0] f692_wdata;
  logic [0:0] f692_clk;
  logic [0:0] f692_rst;
  logic [31:0] f692_rdata;
  sr_buffer_32_1 f692(.wen(f692_wen), .wdata(f692_wdata), .clk(f692_clk), .rst(f692_rst), .rdata(f692_rdata));
  assign f692_clk = clk;
  assign f692_rst = rst;
  // Bindings to f692

  // f694
  logic [0:0] f694_wen;
  logic [31:0] f694_wdata;
  logic [0:0] f694_clk;
  logic [0:0] f694_rst;
  logic [31:0] f694_rdata;
  sr_buffer_32_1 f694(.wen(f694_wen), .wdata(f694_wdata), .clk(f694_clk), .rst(f694_rst), .rdata(f694_rdata));
  assign f694_clk = clk;
  assign f694_rst = rst;
  // Bindings to f694

  // f696
  logic [0:0] f696_wen;
  logic [31:0] f696_wdata;
  logic [0:0] f696_clk;
  logic [0:0] f696_rst;
  logic [31:0] f696_rdata;
  sr_buffer_32_1 f696(.wen(f696_wen), .wdata(f696_wdata), .clk(f696_clk), .rst(f696_rst), .rdata(f696_rdata));
  assign f696_clk = clk;
  assign f696_rst = rst;
  // Bindings to f696

  // f698
  logic [0:0] f698_wen;
  logic [31:0] f698_wdata;
  logic [0:0] f698_clk;
  logic [0:0] f698_rst;
  logic [31:0] f698_rdata;
  sr_buffer_32_1 f698(.wen(f698_wen), .wdata(f698_wdata), .clk(f698_clk), .rst(f698_rst), .rdata(f698_rdata));
  assign f698_clk = clk;
  assign f698_rst = rst;
  // Bindings to f698

  // f700
  logic [0:0] f700_wen;
  logic [31:0] f700_wdata;
  logic [0:0] f700_clk;
  logic [0:0] f700_rst;
  logic [31:0] f700_rdata;
  sr_buffer_32_1 f700(.wen(f700_wen), .wdata(f700_wdata), .clk(f700_clk), .rst(f700_rst), .rdata(f700_rdata));
  assign f700_clk = clk;
  assign f700_rst = rst;
  // Bindings to f700

  // f702
  logic [0:0] f702_wen;
  logic [31:0] f702_wdata;
  logic [0:0] f702_clk;
  logic [0:0] f702_rst;
  logic [31:0] f702_rdata;
  sr_buffer_32_1 f702(.wen(f702_wen), .wdata(f702_wdata), .clk(f702_clk), .rst(f702_rst), .rdata(f702_rdata));
  assign f702_clk = clk;
  assign f702_rst = rst;
  // Bindings to f702

  // f704
  logic [0:0] f704_wen;
  logic [31:0] f704_wdata;
  logic [0:0] f704_clk;
  logic [0:0] f704_rst;
  logic [31:0] f704_rdata;
  sr_buffer_32_1 f704(.wen(f704_wen), .wdata(f704_wdata), .clk(f704_clk), .rst(f704_rst), .rdata(f704_rdata));
  assign f704_clk = clk;
  assign f704_rst = rst;
  // Bindings to f704

  // f706
  logic [0:0] f706_wen;
  logic [31:0] f706_wdata;
  logic [0:0] f706_clk;
  logic [0:0] f706_rst;
  logic [31:0] f706_rdata;
  sr_buffer_32_1 f706(.wen(f706_wen), .wdata(f706_wdata), .clk(f706_clk), .rst(f706_rst), .rdata(f706_rdata));
  assign f706_clk = clk;
  assign f706_rst = rst;
  // Bindings to f706

  // f708
  logic [0:0] f708_wen;
  logic [31:0] f708_wdata;
  logic [0:0] f708_clk;
  logic [0:0] f708_rst;
  logic [31:0] f708_rdata;
  sr_buffer_32_1 f708(.wen(f708_wen), .wdata(f708_wdata), .clk(f708_clk), .rst(f708_rst), .rdata(f708_rdata));
  assign f708_clk = clk;
  assign f708_rst = rst;
  // Bindings to f708

  // f710
  logic [0:0] f710_wen;
  logic [31:0] f710_wdata;
  logic [0:0] f710_clk;
  logic [0:0] f710_rst;
  logic [31:0] f710_rdata;
  sr_buffer_32_1 f710(.wen(f710_wen), .wdata(f710_wdata), .clk(f710_clk), .rst(f710_rst), .rdata(f710_rdata));
  assign f710_clk = clk;
  assign f710_rst = rst;
  // Bindings to f710

  // f712
  logic [0:0] f712_wen;
  logic [31:0] f712_wdata;
  logic [0:0] f712_clk;
  logic [0:0] f712_rst;
  logic [31:0] f712_rdata;
  sr_buffer_32_1 f712(.wen(f712_wen), .wdata(f712_wdata), .clk(f712_clk), .rst(f712_rst), .rdata(f712_rdata));
  assign f712_clk = clk;
  assign f712_rst = rst;
  // Bindings to f712

  // f714
  logic [0:0] f714_wen;
  logic [31:0] f714_wdata;
  logic [0:0] f714_clk;
  logic [0:0] f714_rst;
  logic [31:0] f714_rdata;
  sr_buffer_32_1 f714(.wen(f714_wen), .wdata(f714_wdata), .clk(f714_clk), .rst(f714_rst), .rdata(f714_rdata));
  assign f714_clk = clk;
  assign f714_rst = rst;
  // Bindings to f714

  // f716
  logic [0:0] f716_wen;
  logic [31:0] f716_wdata;
  logic [0:0] f716_clk;
  logic [0:0] f716_rst;
  logic [31:0] f716_rdata;
  sr_buffer_32_1 f716(.wen(f716_wen), .wdata(f716_wdata), .clk(f716_clk), .rst(f716_rst), .rdata(f716_rdata));
  assign f716_clk = clk;
  assign f716_rst = rst;
  // Bindings to f716

  // f718
  logic [0:0] f718_wen;
  logic [31:0] f718_wdata;
  logic [0:0] f718_clk;
  logic [0:0] f718_rst;
  logic [31:0] f718_rdata;
  sr_buffer_32_1 f718(.wen(f718_wen), .wdata(f718_wdata), .clk(f718_clk), .rst(f718_rst), .rdata(f718_rdata));
  assign f718_clk = clk;
  assign f718_rst = rst;
  // Bindings to f718

  // f720
  logic [0:0] f720_wen;
  logic [31:0] f720_wdata;
  logic [0:0] f720_clk;
  logic [0:0] f720_rst;
  logic [31:0] f720_rdata;
  sr_buffer_32_1 f720(.wen(f720_wen), .wdata(f720_wdata), .clk(f720_clk), .rst(f720_rst), .rdata(f720_rdata));
  assign f720_clk = clk;
  assign f720_rst = rst;
  // Bindings to f720

  // f722
  logic [0:0] f722_wen;
  logic [31:0] f722_wdata;
  logic [0:0] f722_clk;
  logic [0:0] f722_rst;
  logic [31:0] f722_rdata;
  sr_buffer_32_1 f722(.wen(f722_wen), .wdata(f722_wdata), .clk(f722_clk), .rst(f722_rst), .rdata(f722_rdata));
  assign f722_clk = clk;
  assign f722_rst = rst;
  // Bindings to f722

  // f724
  logic [0:0] f724_wen;
  logic [31:0] f724_wdata;
  logic [0:0] f724_clk;
  logic [0:0] f724_rst;
  logic [31:0] f724_rdata;
  sr_buffer_32_1 f724(.wen(f724_wen), .wdata(f724_wdata), .clk(f724_clk), .rst(f724_rst), .rdata(f724_rdata));
  assign f724_clk = clk;
  assign f724_rst = rst;
  // Bindings to f724

  // f726
  logic [0:0] f726_wen;
  logic [31:0] f726_wdata;
  logic [0:0] f726_clk;
  logic [0:0] f726_rst;
  logic [31:0] f726_rdata;
  sr_buffer_32_1 f726(.wen(f726_wen), .wdata(f726_wdata), .clk(f726_clk), .rst(f726_rst), .rdata(f726_rdata));
  assign f726_clk = clk;
  assign f726_rst = rst;
  // Bindings to f726

  // f728
  logic [0:0] f728_wen;
  logic [31:0] f728_wdata;
  logic [0:0] f728_clk;
  logic [0:0] f728_rst;
  logic [31:0] f728_rdata;
  sr_buffer_32_1 f728(.wen(f728_wen), .wdata(f728_wdata), .clk(f728_clk), .rst(f728_rst), .rdata(f728_rdata));
  assign f728_clk = clk;
  assign f728_rst = rst;
  // Bindings to f728

  // f730
  logic [0:0] f730_wen;
  logic [31:0] f730_wdata;
  logic [0:0] f730_clk;
  logic [0:0] f730_rst;
  logic [31:0] f730_rdata;
  sr_buffer_32_1 f730(.wen(f730_wen), .wdata(f730_wdata), .clk(f730_clk), .rst(f730_rst), .rdata(f730_rdata));
  assign f730_clk = clk;
  assign f730_rst = rst;
  // Bindings to f730

  // f732
  logic [0:0] f732_wen;
  logic [31:0] f732_wdata;
  logic [0:0] f732_clk;
  logic [0:0] f732_rst;
  logic [31:0] f732_rdata;
  sr_buffer_32_1 f732(.wen(f732_wen), .wdata(f732_wdata), .clk(f732_clk), .rst(f732_rst), .rdata(f732_rdata));
  assign f732_clk = clk;
  assign f732_rst = rst;
  // Bindings to f732

  // f734
  logic [0:0] f734_wen;
  logic [31:0] f734_wdata;
  logic [0:0] f734_clk;
  logic [0:0] f734_rst;
  logic [31:0] f734_rdata;
  sr_buffer_32_1 f734(.wen(f734_wen), .wdata(f734_wdata), .clk(f734_clk), .rst(f734_rst), .rdata(f734_rdata));
  assign f734_clk = clk;
  assign f734_rst = rst;
  // Bindings to f734

  // f736
  logic [0:0] f736_wen;
  logic [31:0] f736_wdata;
  logic [0:0] f736_clk;
  logic [0:0] f736_rst;
  logic [31:0] f736_rdata;
  sr_buffer_32_1 f736(.wen(f736_wen), .wdata(f736_wdata), .clk(f736_clk), .rst(f736_rst), .rdata(f736_rdata));
  assign f736_clk = clk;
  assign f736_rst = rst;
  // Bindings to f736

  // f738
  logic [0:0] f738_wen;
  logic [31:0] f738_wdata;
  logic [0:0] f738_clk;
  logic [0:0] f738_rst;
  logic [31:0] f738_rdata;
  sr_buffer_32_1 f738(.wen(f738_wen), .wdata(f738_wdata), .clk(f738_clk), .rst(f738_rst), .rdata(f738_rdata));
  assign f738_clk = clk;
  assign f738_rst = rst;
  // Bindings to f738

  // f740
  logic [0:0] f740_wen;
  logic [31:0] f740_wdata;
  logic [0:0] f740_clk;
  logic [0:0] f740_rst;
  logic [31:0] f740_rdata;
  sr_buffer_32_1 f740(.wen(f740_wen), .wdata(f740_wdata), .clk(f740_clk), .rst(f740_rst), .rdata(f740_rdata));
  assign f740_clk = clk;
  assign f740_rst = rst;
  // Bindings to f740

  // f742
  logic [0:0] f742_wen;
  logic [31:0] f742_wdata;
  logic [0:0] f742_clk;
  logic [0:0] f742_rst;
  logic [31:0] f742_rdata;
  sr_buffer_32_1 f742(.wen(f742_wen), .wdata(f742_wdata), .clk(f742_clk), .rst(f742_rst), .rdata(f742_rdata));
  assign f742_clk = clk;
  assign f742_rst = rst;
  // Bindings to f742

  // f744
  logic [0:0] f744_wen;
  logic [31:0] f744_wdata;
  logic [0:0] f744_clk;
  logic [0:0] f744_rst;
  logic [31:0] f744_rdata;
  sr_buffer_32_1 f744(.wen(f744_wen), .wdata(f744_wdata), .clk(f744_clk), .rst(f744_rst), .rdata(f744_rdata));
  assign f744_clk = clk;
  assign f744_rst = rst;
  // Bindings to f744

  // f746
  logic [0:0] f746_wen;
  logic [31:0] f746_wdata;
  logic [0:0] f746_clk;
  logic [0:0] f746_rst;
  logic [31:0] f746_rdata;
  sr_buffer_32_1 f746(.wen(f746_wen), .wdata(f746_wdata), .clk(f746_clk), .rst(f746_rst), .rdata(f746_rdata));
  assign f746_clk = clk;
  assign f746_rst = rst;
  // Bindings to f746

  // f748
  logic [0:0] f748_wen;
  logic [31:0] f748_wdata;
  logic [0:0] f748_clk;
  logic [0:0] f748_rst;
  logic [31:0] f748_rdata;
  sr_buffer_32_1 f748(.wen(f748_wen), .wdata(f748_wdata), .clk(f748_clk), .rst(f748_rst), .rdata(f748_rdata));
  assign f748_clk = clk;
  assign f748_rst = rst;
  // Bindings to f748

  // f750
  logic [0:0] f750_wen;
  logic [31:0] f750_wdata;
  logic [0:0] f750_clk;
  logic [0:0] f750_rst;
  logic [31:0] f750_rdata;
  sr_buffer_32_1 f750(.wen(f750_wen), .wdata(f750_wdata), .clk(f750_clk), .rst(f750_rst), .rdata(f750_rdata));
  assign f750_clk = clk;
  assign f750_rst = rst;
  // Bindings to f750

  // f752
  logic [0:0] f752_wen;
  logic [31:0] f752_wdata;
  logic [0:0] f752_clk;
  logic [0:0] f752_rst;
  logic [31:0] f752_rdata;
  sr_buffer_32_1 f752(.wen(f752_wen), .wdata(f752_wdata), .clk(f752_clk), .rst(f752_rst), .rdata(f752_rdata));
  assign f752_clk = clk;
  assign f752_rst = rst;
  // Bindings to f752

  // f754
  logic [0:0] f754_wen;
  logic [31:0] f754_wdata;
  logic [0:0] f754_clk;
  logic [0:0] f754_rst;
  logic [31:0] f754_rdata;
  sr_buffer_32_1 f754(.wen(f754_wen), .wdata(f754_wdata), .clk(f754_clk), .rst(f754_rst), .rdata(f754_rdata));
  assign f754_clk = clk;
  assign f754_rst = rst;
  // Bindings to f754

  // f756
  logic [0:0] f756_wen;
  logic [31:0] f756_wdata;
  logic [0:0] f756_clk;
  logic [0:0] f756_rst;
  logic [31:0] f756_rdata;
  sr_buffer_32_1 f756(.wen(f756_wen), .wdata(f756_wdata), .clk(f756_clk), .rst(f756_rst), .rdata(f756_rdata));
  assign f756_clk = clk;
  assign f756_rst = rst;
  // Bindings to f756

  // f758
  logic [0:0] f758_wen;
  logic [31:0] f758_wdata;
  logic [0:0] f758_clk;
  logic [0:0] f758_rst;
  logic [31:0] f758_rdata;
  sr_buffer_32_1 f758(.wen(f758_wen), .wdata(f758_wdata), .clk(f758_clk), .rst(f758_rst), .rdata(f758_rdata));
  assign f758_clk = clk;
  assign f758_rst = rst;
  // Bindings to f758

  // f760
  logic [0:0] f760_wen;
  logic [31:0] f760_wdata;
  logic [0:0] f760_clk;
  logic [0:0] f760_rst;
  logic [31:0] f760_rdata;
  sr_buffer_32_1 f760(.wen(f760_wen), .wdata(f760_wdata), .clk(f760_clk), .rst(f760_rst), .rdata(f760_rdata));
  assign f760_clk = clk;
  assign f760_rst = rst;
  // Bindings to f760

  // f762
  logic [0:0] f762_wen;
  logic [31:0] f762_wdata;
  logic [0:0] f762_clk;
  logic [0:0] f762_rst;
  logic [31:0] f762_rdata;
  sr_buffer_32_1 f762(.wen(f762_wen), .wdata(f762_wdata), .clk(f762_clk), .rst(f762_rst), .rdata(f762_rdata));
  assign f762_clk = clk;
  assign f762_rst = rst;
  // Bindings to f762

  // f764
  logic [0:0] f764_wen;
  logic [31:0] f764_wdata;
  logic [0:0] f764_clk;
  logic [0:0] f764_rst;
  logic [31:0] f764_rdata;
  sr_buffer_32_1 f764(.wen(f764_wen), .wdata(f764_wdata), .clk(f764_clk), .rst(f764_rst), .rdata(f764_rdata));
  assign f764_clk = clk;
  assign f764_rst = rst;
  // Bindings to f764

  // f766
  logic [0:0] f766_wen;
  logic [31:0] f766_wdata;
  logic [0:0] f766_clk;
  logic [0:0] f766_rst;
  logic [31:0] f766_rdata;
  sr_buffer_32_1 f766(.wen(f766_wen), .wdata(f766_wdata), .clk(f766_clk), .rst(f766_rst), .rdata(f766_rdata));
  assign f766_clk = clk;
  assign f766_rst = rst;
  // Bindings to f766

  // f768
  logic [0:0] f768_wen;
  logic [31:0] f768_wdata;
  logic [0:0] f768_clk;
  logic [0:0] f768_rst;
  logic [31:0] f768_rdata;
  sr_buffer_32_1 f768(.wen(f768_wen), .wdata(f768_wdata), .clk(f768_clk), .rst(f768_rst), .rdata(f768_rdata));
  assign f768_clk = clk;
  assign f768_rst = rst;
  // Bindings to f768

  // f770
  logic [0:0] f770_wen;
  logic [31:0] f770_wdata;
  logic [0:0] f770_clk;
  logic [0:0] f770_rst;
  logic [31:0] f770_rdata;
  sr_buffer_32_1 f770(.wen(f770_wen), .wdata(f770_wdata), .clk(f770_clk), .rst(f770_rst), .rdata(f770_rdata));
  assign f770_clk = clk;
  assign f770_rst = rst;
  // Bindings to f770

  // f772
  logic [0:0] f772_wen;
  logic [31:0] f772_wdata;
  logic [0:0] f772_clk;
  logic [0:0] f772_rst;
  logic [31:0] f772_rdata;
  sr_buffer_32_1 f772(.wen(f772_wen), .wdata(f772_wdata), .clk(f772_clk), .rst(f772_rst), .rdata(f772_rdata));
  assign f772_clk = clk;
  assign f772_rst = rst;
  // Bindings to f772

  // f774
  logic [0:0] f774_wen;
  logic [31:0] f774_wdata;
  logic [0:0] f774_clk;
  logic [0:0] f774_rst;
  logic [31:0] f774_rdata;
  sr_buffer_32_1 f774(.wen(f774_wen), .wdata(f774_wdata), .clk(f774_clk), .rst(f774_rst), .rdata(f774_rdata));
  assign f774_clk = clk;
  assign f774_rst = rst;
  // Bindings to f774

  // f776
  logic [0:0] f776_wen;
  logic [31:0] f776_wdata;
  logic [0:0] f776_clk;
  logic [0:0] f776_rst;
  logic [31:0] f776_rdata;
  sr_buffer_32_1 f776(.wen(f776_wen), .wdata(f776_wdata), .clk(f776_clk), .rst(f776_rst), .rdata(f776_rdata));
  assign f776_clk = clk;
  assign f776_rst = rst;
  // Bindings to f776

  // f778
  logic [0:0] f778_wen;
  logic [31:0] f778_wdata;
  logic [0:0] f778_clk;
  logic [0:0] f778_rst;
  logic [31:0] f778_rdata;
  sr_buffer_32_1 f778(.wen(f778_wen), .wdata(f778_wdata), .clk(f778_clk), .rst(f778_rst), .rdata(f778_rdata));
  assign f778_clk = clk;
  assign f778_rst = rst;
  // Bindings to f778

  // f780
  logic [0:0] f780_wen;
  logic [31:0] f780_wdata;
  logic [0:0] f780_clk;
  logic [0:0] f780_rst;
  logic [31:0] f780_rdata;
  sr_buffer_32_1 f780(.wen(f780_wen), .wdata(f780_wdata), .clk(f780_clk), .rst(f780_rst), .rdata(f780_rdata));
  assign f780_clk = clk;
  assign f780_rst = rst;
  // Bindings to f780

  // f782
  logic [0:0] f782_wen;
  logic [31:0] f782_wdata;
  logic [0:0] f782_clk;
  logic [0:0] f782_rst;
  logic [31:0] f782_rdata;
  sr_buffer_32_1 f782(.wen(f782_wen), .wdata(f782_wdata), .clk(f782_clk), .rst(f782_rst), .rdata(f782_rdata));
  assign f782_clk = clk;
  assign f782_rst = rst;
  // Bindings to f782

  // f784
  logic [0:0] f784_wen;
  logic [31:0] f784_wdata;
  logic [0:0] f784_clk;
  logic [0:0] f784_rst;
  logic [31:0] f784_rdata;
  sr_buffer_32_1 f784(.wen(f784_wen), .wdata(f784_wdata), .clk(f784_clk), .rst(f784_rst), .rdata(f784_rdata));
  assign f784_clk = clk;
  assign f784_rst = rst;
  // Bindings to f784

  // f786
  logic [0:0] f786_wen;
  logic [31:0] f786_wdata;
  logic [0:0] f786_clk;
  logic [0:0] f786_rst;
  logic [31:0] f786_rdata;
  sr_buffer_32_1 f786(.wen(f786_wen), .wdata(f786_wdata), .clk(f786_clk), .rst(f786_rst), .rdata(f786_rdata));
  assign f786_clk = clk;
  assign f786_rst = rst;
  // Bindings to f786

  // f788
  logic [0:0] f788_wen;
  logic [31:0] f788_wdata;
  logic [0:0] f788_clk;
  logic [0:0] f788_rst;
  logic [31:0] f788_rdata;
  sr_buffer_32_1 f788(.wen(f788_wen), .wdata(f788_wdata), .clk(f788_clk), .rst(f788_rst), .rdata(f788_rdata));
  assign f788_clk = clk;
  assign f788_rst = rst;
  // Bindings to f788

  // f790
  logic [0:0] f790_wen;
  logic [31:0] f790_wdata;
  logic [0:0] f790_clk;
  logic [0:0] f790_rst;
  logic [31:0] f790_rdata;
  sr_buffer_32_1 f790(.wen(f790_wen), .wdata(f790_wdata), .clk(f790_clk), .rst(f790_rst), .rdata(f790_rdata));
  assign f790_clk = clk;
  assign f790_rst = rst;
  // Bindings to f790

  // f792
  logic [0:0] f792_wen;
  logic [31:0] f792_wdata;
  logic [0:0] f792_clk;
  logic [0:0] f792_rst;
  logic [31:0] f792_rdata;
  sr_buffer_32_1 f792(.wen(f792_wen), .wdata(f792_wdata), .clk(f792_clk), .rst(f792_rst), .rdata(f792_rdata));
  assign f792_clk = clk;
  assign f792_rst = rst;
  // Bindings to f792

  // f794
  logic [0:0] f794_wen;
  logic [31:0] f794_wdata;
  logic [0:0] f794_clk;
  logic [0:0] f794_rst;
  logic [31:0] f794_rdata;
  sr_buffer_32_1 f794(.wen(f794_wen), .wdata(f794_wdata), .clk(f794_clk), .rst(f794_rst), .rdata(f794_rdata));
  assign f794_clk = clk;
  assign f794_rst = rst;
  // Bindings to f794

  // f796
  logic [0:0] f796_wen;
  logic [31:0] f796_wdata;
  logic [0:0] f796_clk;
  logic [0:0] f796_rst;
  logic [31:0] f796_rdata;
  sr_buffer_32_1 f796(.wen(f796_wen), .wdata(f796_wdata), .clk(f796_clk), .rst(f796_rst), .rdata(f796_rdata));
  assign f796_clk = clk;
  assign f796_rst = rst;
  // Bindings to f796

  // f798
  logic [0:0] f798_wen;
  logic [31:0] f798_wdata;
  logic [0:0] f798_clk;
  logic [0:0] f798_rst;
  logic [31:0] f798_rdata;
  sr_buffer_32_1 f798(.wen(f798_wen), .wdata(f798_wdata), .clk(f798_clk), .rst(f798_rst), .rdata(f798_rdata));
  assign f798_clk = clk;
  assign f798_rst = rst;
  // Bindings to f798

  // f800
  logic [0:0] f800_wen;
  logic [31:0] f800_wdata;
  logic [0:0] f800_clk;
  logic [0:0] f800_rst;
  logic [31:0] f800_rdata;
  sr_buffer_32_1 f800(.wen(f800_wen), .wdata(f800_wdata), .clk(f800_clk), .rst(f800_rst), .rdata(f800_rdata));
  assign f800_clk = clk;
  assign f800_rst = rst;
  // Bindings to f800

  // f802
  logic [0:0] f802_wen;
  logic [31:0] f802_wdata;
  logic [0:0] f802_clk;
  logic [0:0] f802_rst;
  logic [31:0] f802_rdata;
  sr_buffer_32_1 f802(.wen(f802_wen), .wdata(f802_wdata), .clk(f802_clk), .rst(f802_rst), .rdata(f802_rdata));
  assign f802_clk = clk;
  assign f802_rst = rst;
  // Bindings to f802

  // f804
  logic [0:0] f804_wen;
  logic [31:0] f804_wdata;
  logic [0:0] f804_clk;
  logic [0:0] f804_rst;
  logic [31:0] f804_rdata;
  sr_buffer_32_1 f804(.wen(f804_wen), .wdata(f804_wdata), .clk(f804_clk), .rst(f804_rst), .rdata(f804_rdata));
  assign f804_clk = clk;
  assign f804_rst = rst;
  // Bindings to f804

  // f806
  logic [0:0] f806_wen;
  logic [31:0] f806_wdata;
  logic [0:0] f806_clk;
  logic [0:0] f806_rst;
  logic [31:0] f806_rdata;
  sr_buffer_32_1 f806(.wen(f806_wen), .wdata(f806_wdata), .clk(f806_clk), .rst(f806_rst), .rdata(f806_rdata));
  assign f806_clk = clk;
  assign f806_rst = rst;
  // Bindings to f806

  // f808
  logic [0:0] f808_wen;
  logic [31:0] f808_wdata;
  logic [0:0] f808_clk;
  logic [0:0] f808_rst;
  logic [31:0] f808_rdata;
  sr_buffer_32_1 f808(.wen(f808_wen), .wdata(f808_wdata), .clk(f808_clk), .rst(f808_rst), .rdata(f808_rdata));
  assign f808_clk = clk;
  assign f808_rst = rst;
  // Bindings to f808

  // f810
  logic [0:0] f810_wen;
  logic [31:0] f810_wdata;
  logic [0:0] f810_clk;
  logic [0:0] f810_rst;
  logic [31:0] f810_rdata;
  sr_buffer_32_1 f810(.wen(f810_wen), .wdata(f810_wdata), .clk(f810_clk), .rst(f810_rst), .rdata(f810_rdata));
  assign f810_clk = clk;
  assign f810_rst = rst;
  // Bindings to f810

  // f812
  logic [0:0] f812_wen;
  logic [31:0] f812_wdata;
  logic [0:0] f812_clk;
  logic [0:0] f812_rst;
  logic [31:0] f812_rdata;
  sr_buffer_32_1 f812(.wen(f812_wen), .wdata(f812_wdata), .clk(f812_clk), .rst(f812_rst), .rdata(f812_rdata));
  assign f812_clk = clk;
  assign f812_rst = rst;
  // Bindings to f812

  // f814
  logic [0:0] f814_wen;
  logic [31:0] f814_wdata;
  logic [0:0] f814_clk;
  logic [0:0] f814_rst;
  logic [31:0] f814_rdata;
  sr_buffer_32_1 f814(.wen(f814_wen), .wdata(f814_wdata), .clk(f814_clk), .rst(f814_rst), .rdata(f814_rdata));
  assign f814_clk = clk;
  assign f814_rst = rst;
  // Bindings to f814

  // f816
  logic [0:0] f816_wen;
  logic [31:0] f816_wdata;
  logic [0:0] f816_clk;
  logic [0:0] f816_rst;
  logic [31:0] f816_rdata;
  sr_buffer_32_1 f816(.wen(f816_wen), .wdata(f816_wdata), .clk(f816_clk), .rst(f816_rst), .rdata(f816_rdata));
  assign f816_clk = clk;
  assign f816_rst = rst;
  // Bindings to f816

  // f818
  logic [0:0] f818_wen;
  logic [31:0] f818_wdata;
  logic [0:0] f818_clk;
  logic [0:0] f818_rst;
  logic [31:0] f818_rdata;
  sr_buffer_32_1 f818(.wen(f818_wen), .wdata(f818_wdata), .clk(f818_clk), .rst(f818_rst), .rdata(f818_rdata));
  assign f818_clk = clk;
  assign f818_rst = rst;
  // Bindings to f818

  // f820
  logic [0:0] f820_wen;
  logic [31:0] f820_wdata;
  logic [0:0] f820_clk;
  logic [0:0] f820_rst;
  logic [31:0] f820_rdata;
  sr_buffer_32_1 f820(.wen(f820_wen), .wdata(f820_wdata), .clk(f820_clk), .rst(f820_rst), .rdata(f820_rdata));
  assign f820_clk = clk;
  assign f820_rst = rst;
  // Bindings to f820

  // f822
  logic [0:0] f822_wen;
  logic [31:0] f822_wdata;
  logic [0:0] f822_clk;
  logic [0:0] f822_rst;
  logic [31:0] f822_rdata;
  sr_buffer_32_1 f822(.wen(f822_wen), .wdata(f822_wdata), .clk(f822_clk), .rst(f822_rst), .rdata(f822_rdata));
  assign f822_clk = clk;
  assign f822_rst = rst;
  // Bindings to f822

  // f824
  logic [0:0] f824_wen;
  logic [31:0] f824_wdata;
  logic [0:0] f824_clk;
  logic [0:0] f824_rst;
  logic [31:0] f824_rdata;
  sr_buffer_32_1 f824(.wen(f824_wen), .wdata(f824_wdata), .clk(f824_clk), .rst(f824_rst), .rdata(f824_rdata));
  assign f824_clk = clk;
  assign f824_rst = rst;
  // Bindings to f824

  // f826
  logic [0:0] f826_wen;
  logic [31:0] f826_wdata;
  logic [0:0] f826_clk;
  logic [0:0] f826_rst;
  logic [31:0] f826_rdata;
  sr_buffer_32_1 f826(.wen(f826_wen), .wdata(f826_wdata), .clk(f826_clk), .rst(f826_rst), .rdata(f826_rdata));
  assign f826_clk = clk;
  assign f826_rst = rst;
  // Bindings to f826

  // f828
  logic [0:0] f828_wen;
  logic [31:0] f828_wdata;
  logic [0:0] f828_clk;
  logic [0:0] f828_rst;
  logic [31:0] f828_rdata;
  sr_buffer_32_1 f828(.wen(f828_wen), .wdata(f828_wdata), .clk(f828_clk), .rst(f828_rst), .rdata(f828_rdata));
  assign f828_clk = clk;
  assign f828_rst = rst;
  // Bindings to f828

  // f830
  logic [0:0] f830_wen;
  logic [31:0] f830_wdata;
  logic [0:0] f830_clk;
  logic [0:0] f830_rst;
  logic [31:0] f830_rdata;
  sr_buffer_32_1 f830(.wen(f830_wen), .wdata(f830_wdata), .clk(f830_clk), .rst(f830_rst), .rdata(f830_rdata));
  assign f830_clk = clk;
  assign f830_rst = rst;
  // Bindings to f830

  // f832
  logic [0:0] f832_wen;
  logic [31:0] f832_wdata;
  logic [0:0] f832_clk;
  logic [0:0] f832_rst;
  logic [31:0] f832_rdata;
  sr_buffer_32_1 f832(.wen(f832_wen), .wdata(f832_wdata), .clk(f832_clk), .rst(f832_rst), .rdata(f832_rdata));
  assign f832_clk = clk;
  assign f832_rst = rst;
  // Bindings to f832

  // f834
  logic [0:0] f834_wen;
  logic [31:0] f834_wdata;
  logic [0:0] f834_clk;
  logic [0:0] f834_rst;
  logic [31:0] f834_rdata;
  sr_buffer_32_1 f834(.wen(f834_wen), .wdata(f834_wdata), .clk(f834_clk), .rst(f834_rst), .rdata(f834_rdata));
  assign f834_clk = clk;
  assign f834_rst = rst;
  // Bindings to f834

  // f836
  logic [0:0] f836_wen;
  logic [31:0] f836_wdata;
  logic [0:0] f836_clk;
  logic [0:0] f836_rst;
  logic [31:0] f836_rdata;
  sr_buffer_32_1 f836(.wen(f836_wen), .wdata(f836_wdata), .clk(f836_clk), .rst(f836_rst), .rdata(f836_rdata));
  assign f836_clk = clk;
  assign f836_rst = rst;
  // Bindings to f836

  // f838
  logic [0:0] f838_wen;
  logic [31:0] f838_wdata;
  logic [0:0] f838_clk;
  logic [0:0] f838_rst;
  logic [31:0] f838_rdata;
  sr_buffer_32_1 f838(.wen(f838_wen), .wdata(f838_wdata), .clk(f838_clk), .rst(f838_rst), .rdata(f838_rdata));
  assign f838_clk = clk;
  assign f838_rst = rst;
  // Bindings to f838

  // f840
  logic [0:0] f840_wen;
  logic [31:0] f840_wdata;
  logic [0:0] f840_clk;
  logic [0:0] f840_rst;
  logic [31:0] f840_rdata;
  sr_buffer_32_1 f840(.wen(f840_wen), .wdata(f840_wdata), .clk(f840_clk), .rst(f840_rst), .rdata(f840_rdata));
  assign f840_clk = clk;
  assign f840_rst = rst;
  // Bindings to f840

  // f842
  logic [0:0] f842_wen;
  logic [31:0] f842_wdata;
  logic [0:0] f842_clk;
  logic [0:0] f842_rst;
  logic [31:0] f842_rdata;
  sr_buffer_32_1 f842(.wen(f842_wen), .wdata(f842_wdata), .clk(f842_clk), .rst(f842_rst), .rdata(f842_rdata));
  assign f842_clk = clk;
  assign f842_rst = rst;
  // Bindings to f842

  // f844
  logic [0:0] f844_wen;
  logic [31:0] f844_wdata;
  logic [0:0] f844_clk;
  logic [0:0] f844_rst;
  logic [31:0] f844_rdata;
  sr_buffer_32_1 f844(.wen(f844_wen), .wdata(f844_wdata), .clk(f844_clk), .rst(f844_rst), .rdata(f844_rdata));
  assign f844_clk = clk;
  assign f844_rst = rst;
  // Bindings to f844

  // f846
  logic [0:0] f846_wen;
  logic [31:0] f846_wdata;
  logic [0:0] f846_clk;
  logic [0:0] f846_rst;
  logic [31:0] f846_rdata;
  sr_buffer_32_1 f846(.wen(f846_wen), .wdata(f846_wdata), .clk(f846_clk), .rst(f846_rst), .rdata(f846_rdata));
  assign f846_clk = clk;
  assign f846_rst = rst;
  // Bindings to f846

  // f848
  logic [0:0] f848_wen;
  logic [31:0] f848_wdata;
  logic [0:0] f848_clk;
  logic [0:0] f848_rst;
  logic [31:0] f848_rdata;
  sr_buffer_32_1 f848(.wen(f848_wen), .wdata(f848_wdata), .clk(f848_clk), .rst(f848_rst), .rdata(f848_rdata));
  assign f848_clk = clk;
  assign f848_rst = rst;
  // Bindings to f848

  // f850
  logic [0:0] f850_wen;
  logic [31:0] f850_wdata;
  logic [0:0] f850_clk;
  logic [0:0] f850_rst;
  logic [31:0] f850_rdata;
  sr_buffer_32_1 f850(.wen(f850_wen), .wdata(f850_wdata), .clk(f850_clk), .rst(f850_rst), .rdata(f850_rdata));
  assign f850_clk = clk;
  assign f850_rst = rst;
  // Bindings to f850

  // f852
  logic [0:0] f852_wen;
  logic [31:0] f852_wdata;
  logic [0:0] f852_clk;
  logic [0:0] f852_rst;
  logic [31:0] f852_rdata;
  sr_buffer_32_1 f852(.wen(f852_wen), .wdata(f852_wdata), .clk(f852_clk), .rst(f852_rst), .rdata(f852_rdata));
  assign f852_clk = clk;
  assign f852_rst = rst;
  // Bindings to f852

  // f854
  logic [0:0] f854_wen;
  logic [31:0] f854_wdata;
  logic [0:0] f854_clk;
  logic [0:0] f854_rst;
  logic [31:0] f854_rdata;
  sr_buffer_32_1 f854(.wen(f854_wen), .wdata(f854_wdata), .clk(f854_clk), .rst(f854_rst), .rdata(f854_rdata));
  assign f854_clk = clk;
  assign f854_rst = rst;
  // Bindings to f854

  // f856
  logic [0:0] f856_wen;
  logic [31:0] f856_wdata;
  logic [0:0] f856_clk;
  logic [0:0] f856_rst;
  logic [31:0] f856_rdata;
  sr_buffer_32_1 f856(.wen(f856_wen), .wdata(f856_wdata), .clk(f856_clk), .rst(f856_rst), .rdata(f856_rdata));
  assign f856_clk = clk;
  assign f856_rst = rst;
  // Bindings to f856

  // f858
  logic [0:0] f858_wen;
  logic [31:0] f858_wdata;
  logic [0:0] f858_clk;
  logic [0:0] f858_rst;
  logic [31:0] f858_rdata;
  sr_buffer_32_1 f858(.wen(f858_wen), .wdata(f858_wdata), .clk(f858_clk), .rst(f858_rst), .rdata(f858_rdata));
  assign f858_clk = clk;
  assign f858_rst = rst;
  // Bindings to f858

  // f860
  logic [0:0] f860_wen;
  logic [31:0] f860_wdata;
  logic [0:0] f860_clk;
  logic [0:0] f860_rst;
  logic [31:0] f860_rdata;
  sr_buffer_32_1 f860(.wen(f860_wen), .wdata(f860_wdata), .clk(f860_clk), .rst(f860_rst), .rdata(f860_rdata));
  assign f860_clk = clk;
  assign f860_rst = rst;
  // Bindings to f860

  // f862
  logic [0:0] f862_wen;
  logic [31:0] f862_wdata;
  logic [0:0] f862_clk;
  logic [0:0] f862_rst;
  logic [31:0] f862_rdata;
  sr_buffer_32_1 f862(.wen(f862_wen), .wdata(f862_wdata), .clk(f862_clk), .rst(f862_rst), .rdata(f862_rdata));
  assign f862_clk = clk;
  assign f862_rst = rst;
  // Bindings to f862

  // f864
  logic [0:0] f864_wen;
  logic [31:0] f864_wdata;
  logic [0:0] f864_clk;
  logic [0:0] f864_rst;
  logic [31:0] f864_rdata;
  sr_buffer_32_1 f864(.wen(f864_wen), .wdata(f864_wdata), .clk(f864_clk), .rst(f864_rst), .rdata(f864_rdata));
  assign f864_clk = clk;
  assign f864_rst = rst;
  // Bindings to f864

  // f866
  logic [0:0] f866_wen;
  logic [31:0] f866_wdata;
  logic [0:0] f866_clk;
  logic [0:0] f866_rst;
  logic [31:0] f866_rdata;
  sr_buffer_32_1 f866(.wen(f866_wen), .wdata(f866_wdata), .clk(f866_clk), .rst(f866_rst), .rdata(f866_rdata));
  assign f866_clk = clk;
  assign f866_rst = rst;
  // Bindings to f866

  // f868
  logic [0:0] f868_wen;
  logic [31:0] f868_wdata;
  logic [0:0] f868_clk;
  logic [0:0] f868_rst;
  logic [31:0] f868_rdata;
  sr_buffer_32_1 f868(.wen(f868_wen), .wdata(f868_wdata), .clk(f868_clk), .rst(f868_rst), .rdata(f868_rdata));
  assign f868_clk = clk;
  assign f868_rst = rst;
  // Bindings to f868

  // f870
  logic [0:0] f870_wen;
  logic [31:0] f870_wdata;
  logic [0:0] f870_clk;
  logic [0:0] f870_rst;
  logic [31:0] f870_rdata;
  sr_buffer_32_1 f870(.wen(f870_wen), .wdata(f870_wdata), .clk(f870_clk), .rst(f870_rst), .rdata(f870_rdata));
  assign f870_clk = clk;
  assign f870_rst = rst;
  // Bindings to f870

  // f872
  logic [0:0] f872_wen;
  logic [31:0] f872_wdata;
  logic [0:0] f872_clk;
  logic [0:0] f872_rst;
  logic [31:0] f872_rdata;
  sr_buffer_32_1 f872(.wen(f872_wen), .wdata(f872_wdata), .clk(f872_clk), .rst(f872_rst), .rdata(f872_rdata));
  assign f872_clk = clk;
  assign f872_rst = rst;
  // Bindings to f872

  // f874
  logic [0:0] f874_wen;
  logic [31:0] f874_wdata;
  logic [0:0] f874_clk;
  logic [0:0] f874_rst;
  logic [31:0] f874_rdata;
  sr_buffer_32_1 f874(.wen(f874_wen), .wdata(f874_wdata), .clk(f874_clk), .rst(f874_rst), .rdata(f874_rdata));
  assign f874_clk = clk;
  assign f874_rst = rst;
  // Bindings to f874

  // f876
  logic [0:0] f876_wen;
  logic [31:0] f876_wdata;
  logic [0:0] f876_clk;
  logic [0:0] f876_rst;
  logic [31:0] f876_rdata;
  sr_buffer_32_1 f876(.wen(f876_wen), .wdata(f876_wdata), .clk(f876_clk), .rst(f876_rst), .rdata(f876_rdata));
  assign f876_clk = clk;
  assign f876_rst = rst;
  // Bindings to f876

  // f878
  logic [0:0] f878_wen;
  logic [31:0] f878_wdata;
  logic [0:0] f878_clk;
  logic [0:0] f878_rst;
  logic [31:0] f878_rdata;
  sr_buffer_32_1 f878(.wen(f878_wen), .wdata(f878_wdata), .clk(f878_clk), .rst(f878_rst), .rdata(f878_rdata));
  assign f878_clk = clk;
  assign f878_rst = rst;
  // Bindings to f878

  // f880
  logic [0:0] f880_wen;
  logic [31:0] f880_wdata;
  logic [0:0] f880_clk;
  logic [0:0] f880_rst;
  logic [31:0] f880_rdata;
  sr_buffer_32_1 f880(.wen(f880_wen), .wdata(f880_wdata), .clk(f880_clk), .rst(f880_rst), .rdata(f880_rdata));
  assign f880_clk = clk;
  assign f880_rst = rst;
  // Bindings to f880

  // f882
  logic [0:0] f882_wen;
  logic [31:0] f882_wdata;
  logic [0:0] f882_clk;
  logic [0:0] f882_rst;
  logic [31:0] f882_rdata;
  sr_buffer_32_1 f882(.wen(f882_wen), .wdata(f882_wdata), .clk(f882_clk), .rst(f882_rst), .rdata(f882_rdata));
  assign f882_clk = clk;
  assign f882_rst = rst;
  // Bindings to f882

  // f884
  logic [0:0] f884_wen;
  logic [31:0] f884_wdata;
  logic [0:0] f884_clk;
  logic [0:0] f884_rst;
  logic [31:0] f884_rdata;
  sr_buffer_32_1 f884(.wen(f884_wen), .wdata(f884_wdata), .clk(f884_clk), .rst(f884_rst), .rdata(f884_rdata));
  assign f884_clk = clk;
  assign f884_rst = rst;
  // Bindings to f884

  // f886
  logic [0:0] f886_wen;
  logic [31:0] f886_wdata;
  logic [0:0] f886_clk;
  logic [0:0] f886_rst;
  logic [31:0] f886_rdata;
  sr_buffer_32_1 f886(.wen(f886_wen), .wdata(f886_wdata), .clk(f886_clk), .rst(f886_rst), .rdata(f886_rdata));
  assign f886_clk = clk;
  assign f886_rst = rst;
  // Bindings to f886

  // f888
  logic [0:0] f888_wen;
  logic [31:0] f888_wdata;
  logic [0:0] f888_clk;
  logic [0:0] f888_rst;
  logic [31:0] f888_rdata;
  sr_buffer_32_1 f888(.wen(f888_wen), .wdata(f888_wdata), .clk(f888_clk), .rst(f888_rst), .rdata(f888_rdata));
  assign f888_clk = clk;
  assign f888_rst = rst;
  // Bindings to f888

  // f890
  logic [0:0] f890_wen;
  logic [31:0] f890_wdata;
  logic [0:0] f890_clk;
  logic [0:0] f890_rst;
  logic [31:0] f890_rdata;
  sr_buffer_32_1 f890(.wen(f890_wen), .wdata(f890_wdata), .clk(f890_clk), .rst(f890_rst), .rdata(f890_rdata));
  assign f890_clk = clk;
  assign f890_rst = rst;
  // Bindings to f890

  // f892
  logic [0:0] f892_wen;
  logic [31:0] f892_wdata;
  logic [0:0] f892_clk;
  logic [0:0] f892_rst;
  logic [31:0] f892_rdata;
  sr_buffer_32_1 f892(.wen(f892_wen), .wdata(f892_wdata), .clk(f892_clk), .rst(f892_rst), .rdata(f892_rdata));
  assign f892_clk = clk;
  assign f892_rst = rst;
  // Bindings to f892

  // f894
  logic [0:0] f894_wen;
  logic [31:0] f894_wdata;
  logic [0:0] f894_clk;
  logic [0:0] f894_rst;
  logic [31:0] f894_rdata;
  sr_buffer_32_1 f894(.wen(f894_wen), .wdata(f894_wdata), .clk(f894_clk), .rst(f894_rst), .rdata(f894_rdata));
  assign f894_clk = clk;
  assign f894_rst = rst;
  // Bindings to f894

  // f896
  logic [0:0] f896_wen;
  logic [31:0] f896_wdata;
  logic [0:0] f896_clk;
  logic [0:0] f896_rst;
  logic [31:0] f896_rdata;
  sr_buffer_32_1 f896(.wen(f896_wen), .wdata(f896_wdata), .clk(f896_clk), .rst(f896_rst), .rdata(f896_rdata));
  assign f896_clk = clk;
  assign f896_rst = rst;
  // Bindings to f896

  // f898
  logic [0:0] f898_wen;
  logic [31:0] f898_wdata;
  logic [0:0] f898_clk;
  logic [0:0] f898_rst;
  logic [31:0] f898_rdata;
  sr_buffer_32_1 f898(.wen(f898_wen), .wdata(f898_wdata), .clk(f898_clk), .rst(f898_rst), .rdata(f898_rdata));
  assign f898_clk = clk;
  assign f898_rst = rst;
  // Bindings to f898

  // f900
  logic [0:0] f900_wen;
  logic [31:0] f900_wdata;
  logic [0:0] f900_clk;
  logic [0:0] f900_rst;
  logic [31:0] f900_rdata;
  sr_buffer_32_1 f900(.wen(f900_wen), .wdata(f900_wdata), .clk(f900_clk), .rst(f900_rst), .rdata(f900_rdata));
  assign f900_clk = clk;
  assign f900_rst = rst;
  // Bindings to f900

  // f902
  logic [0:0] f902_wen;
  logic [31:0] f902_wdata;
  logic [0:0] f902_clk;
  logic [0:0] f902_rst;
  logic [31:0] f902_rdata;
  sr_buffer_32_1 f902(.wen(f902_wen), .wdata(f902_wdata), .clk(f902_clk), .rst(f902_rst), .rdata(f902_rdata));
  assign f902_clk = clk;
  assign f902_rst = rst;
  // Bindings to f902

  // f904
  logic [0:0] f904_wen;
  logic [31:0] f904_wdata;
  logic [0:0] f904_clk;
  logic [0:0] f904_rst;
  logic [31:0] f904_rdata;
  sr_buffer_32_1 f904(.wen(f904_wen), .wdata(f904_wdata), .clk(f904_clk), .rst(f904_rst), .rdata(f904_rdata));
  assign f904_clk = clk;
  assign f904_rst = rst;
  // Bindings to f904

  // f906
  logic [0:0] f906_wen;
  logic [31:0] f906_wdata;
  logic [0:0] f906_clk;
  logic [0:0] f906_rst;
  logic [31:0] f906_rdata;
  sr_buffer_32_1 f906(.wen(f906_wen), .wdata(f906_wdata), .clk(f906_clk), .rst(f906_rst), .rdata(f906_rdata));
  assign f906_clk = clk;
  assign f906_rst = rst;
  // Bindings to f906

  // f908
  logic [0:0] f908_wen;
  logic [31:0] f908_wdata;
  logic [0:0] f908_clk;
  logic [0:0] f908_rst;
  logic [31:0] f908_rdata;
  sr_buffer_32_1 f908(.wen(f908_wen), .wdata(f908_wdata), .clk(f908_clk), .rst(f908_rst), .rdata(f908_rdata));
  assign f908_clk = clk;
  assign f908_rst = rst;
  // Bindings to f908

  // f910
  logic [0:0] f910_wen;
  logic [31:0] f910_wdata;
  logic [0:0] f910_clk;
  logic [0:0] f910_rst;
  logic [31:0] f910_rdata;
  sr_buffer_32_1 f910(.wen(f910_wen), .wdata(f910_wdata), .clk(f910_clk), .rst(f910_rst), .rdata(f910_rdata));
  assign f910_clk = clk;
  assign f910_rst = rst;
  // Bindings to f910

  // f912
  logic [0:0] f912_wen;
  logic [31:0] f912_wdata;
  logic [0:0] f912_clk;
  logic [0:0] f912_rst;
  logic [31:0] f912_rdata;
  sr_buffer_32_1 f912(.wen(f912_wen), .wdata(f912_wdata), .clk(f912_clk), .rst(f912_rst), .rdata(f912_rdata));
  assign f912_clk = clk;
  assign f912_rst = rst;
  // Bindings to f912

  // f914
  logic [0:0] f914_wen;
  logic [31:0] f914_wdata;
  logic [0:0] f914_clk;
  logic [0:0] f914_rst;
  logic [31:0] f914_rdata;
  sr_buffer_32_1 f914(.wen(f914_wen), .wdata(f914_wdata), .clk(f914_clk), .rst(f914_rst), .rdata(f914_rdata));
  assign f914_clk = clk;
  assign f914_rst = rst;
  // Bindings to f914

  // f916
  logic [0:0] f916_wen;
  logic [31:0] f916_wdata;
  logic [0:0] f916_clk;
  logic [0:0] f916_rst;
  logic [31:0] f916_rdata;
  sr_buffer_32_1 f916(.wen(f916_wen), .wdata(f916_wdata), .clk(f916_clk), .rst(f916_rst), .rdata(f916_rdata));
  assign f916_clk = clk;
  assign f916_rst = rst;
  // Bindings to f916

  // f918
  logic [0:0] f918_wen;
  logic [31:0] f918_wdata;
  logic [0:0] f918_clk;
  logic [0:0] f918_rst;
  logic [31:0] f918_rdata;
  sr_buffer_32_1 f918(.wen(f918_wen), .wdata(f918_wdata), .clk(f918_clk), .rst(f918_rst), .rdata(f918_rdata));
  assign f918_clk = clk;
  assign f918_rst = rst;
  // Bindings to f918

  // f920
  logic [0:0] f920_wen;
  logic [31:0] f920_wdata;
  logic [0:0] f920_clk;
  logic [0:0] f920_rst;
  logic [31:0] f920_rdata;
  sr_buffer_32_1 f920(.wen(f920_wen), .wdata(f920_wdata), .clk(f920_clk), .rst(f920_rst), .rdata(f920_rdata));
  assign f920_clk = clk;
  assign f920_rst = rst;
  // Bindings to f920

  // f922
  logic [0:0] f922_wen;
  logic [31:0] f922_wdata;
  logic [0:0] f922_clk;
  logic [0:0] f922_rst;
  logic [31:0] f922_rdata;
  sr_buffer_32_1 f922(.wen(f922_wen), .wdata(f922_wdata), .clk(f922_clk), .rst(f922_rst), .rdata(f922_rdata));
  assign f922_clk = clk;
  assign f922_rst = rst;
  // Bindings to f922

  // f924
  logic [0:0] f924_wen;
  logic [31:0] f924_wdata;
  logic [0:0] f924_clk;
  logic [0:0] f924_rst;
  logic [31:0] f924_rdata;
  sr_buffer_32_1 f924(.wen(f924_wen), .wdata(f924_wdata), .clk(f924_clk), .rst(f924_rst), .rdata(f924_rdata));
  assign f924_clk = clk;
  assign f924_rst = rst;
  // Bindings to f924

  // f926
  logic [0:0] f926_wen;
  logic [31:0] f926_wdata;
  logic [0:0] f926_clk;
  logic [0:0] f926_rst;
  logic [31:0] f926_rdata;
  sr_buffer_32_1 f926(.wen(f926_wen), .wdata(f926_wdata), .clk(f926_clk), .rst(f926_rst), .rdata(f926_rdata));
  assign f926_clk = clk;
  assign f926_rst = rst;
  // Bindings to f926

  // f928
  logic [0:0] f928_wen;
  logic [31:0] f928_wdata;
  logic [0:0] f928_clk;
  logic [0:0] f928_rst;
  logic [31:0] f928_rdata;
  sr_buffer_32_1 f928(.wen(f928_wen), .wdata(f928_wdata), .clk(f928_clk), .rst(f928_rst), .rdata(f928_rdata));
  assign f928_clk = clk;
  assign f928_rst = rst;
  // Bindings to f928

  // f930
  logic [0:0] f930_wen;
  logic [31:0] f930_wdata;
  logic [0:0] f930_clk;
  logic [0:0] f930_rst;
  logic [31:0] f930_rdata;
  sr_buffer_32_1 f930(.wen(f930_wen), .wdata(f930_wdata), .clk(f930_clk), .rst(f930_rst), .rdata(f930_rdata));
  assign f930_clk = clk;
  assign f930_rst = rst;
  // Bindings to f930

  // f932
  logic [0:0] f932_wen;
  logic [31:0] f932_wdata;
  logic [0:0] f932_clk;
  logic [0:0] f932_rst;
  logic [31:0] f932_rdata;
  sr_buffer_32_1 f932(.wen(f932_wen), .wdata(f932_wdata), .clk(f932_clk), .rst(f932_rst), .rdata(f932_rdata));
  assign f932_clk = clk;
  assign f932_rst = rst;
  // Bindings to f932

  // f934
  logic [0:0] f934_wen;
  logic [31:0] f934_wdata;
  logic [0:0] f934_clk;
  logic [0:0] f934_rst;
  logic [31:0] f934_rdata;
  sr_buffer_32_1 f934(.wen(f934_wen), .wdata(f934_wdata), .clk(f934_clk), .rst(f934_rst), .rdata(f934_rdata));
  assign f934_clk = clk;
  assign f934_rst = rst;
  // Bindings to f934

  // f936
  logic [0:0] f936_wen;
  logic [31:0] f936_wdata;
  logic [0:0] f936_clk;
  logic [0:0] f936_rst;
  logic [31:0] f936_rdata;
  sr_buffer_32_1 f936(.wen(f936_wen), .wdata(f936_wdata), .clk(f936_clk), .rst(f936_rst), .rdata(f936_rdata));
  assign f936_clk = clk;
  assign f936_rst = rst;
  // Bindings to f936

  // f938
  logic [0:0] f938_wen;
  logic [31:0] f938_wdata;
  logic [0:0] f938_clk;
  logic [0:0] f938_rst;
  logic [31:0] f938_rdata;
  sr_buffer_32_1 f938(.wen(f938_wen), .wdata(f938_wdata), .clk(f938_clk), .rst(f938_rst), .rdata(f938_rdata));
  assign f938_clk = clk;
  assign f938_rst = rst;
  // Bindings to f938

  // f940
  logic [0:0] f940_wen;
  logic [31:0] f940_wdata;
  logic [0:0] f940_clk;
  logic [0:0] f940_rst;
  logic [31:0] f940_rdata;
  sr_buffer_32_1 f940(.wen(f940_wen), .wdata(f940_wdata), .clk(f940_clk), .rst(f940_rst), .rdata(f940_rdata));
  assign f940_clk = clk;
  assign f940_rst = rst;
  // Bindings to f940

  // f942
  logic [0:0] f942_wen;
  logic [31:0] f942_wdata;
  logic [0:0] f942_clk;
  logic [0:0] f942_rst;
  logic [31:0] f942_rdata;
  sr_buffer_32_1 f942(.wen(f942_wen), .wdata(f942_wdata), .clk(f942_clk), .rst(f942_rst), .rdata(f942_rdata));
  assign f942_clk = clk;
  assign f942_rst = rst;
  // Bindings to f942

  // f944
  logic [0:0] f944_wen;
  logic [31:0] f944_wdata;
  logic [0:0] f944_clk;
  logic [0:0] f944_rst;
  logic [31:0] f944_rdata;
  sr_buffer_32_1 f944(.wen(f944_wen), .wdata(f944_wdata), .clk(f944_clk), .rst(f944_rst), .rdata(f944_rdata));
  assign f944_clk = clk;
  assign f944_rst = rst;
  // Bindings to f944

  // f946
  logic [0:0] f946_wen;
  logic [31:0] f946_wdata;
  logic [0:0] f946_clk;
  logic [0:0] f946_rst;
  logic [31:0] f946_rdata;
  sr_buffer_32_1 f946(.wen(f946_wen), .wdata(f946_wdata), .clk(f946_clk), .rst(f946_rst), .rdata(f946_rdata));
  assign f946_clk = clk;
  assign f946_rst = rst;
  // Bindings to f946

  // f948
  logic [0:0] f948_wen;
  logic [31:0] f948_wdata;
  logic [0:0] f948_clk;
  logic [0:0] f948_rst;
  logic [31:0] f948_rdata;
  sr_buffer_32_1 f948(.wen(f948_wen), .wdata(f948_wdata), .clk(f948_clk), .rst(f948_rst), .rdata(f948_rdata));
  assign f948_clk = clk;
  assign f948_rst = rst;
  // Bindings to f948

  // f950
  logic [0:0] f950_wen;
  logic [31:0] f950_wdata;
  logic [0:0] f950_clk;
  logic [0:0] f950_rst;
  logic [31:0] f950_rdata;
  sr_buffer_32_1 f950(.wen(f950_wen), .wdata(f950_wdata), .clk(f950_clk), .rst(f950_rst), .rdata(f950_rdata));
  assign f950_clk = clk;
  assign f950_rst = rst;
  // Bindings to f950

  // f952
  logic [0:0] f952_wen;
  logic [31:0] f952_wdata;
  logic [0:0] f952_clk;
  logic [0:0] f952_rst;
  logic [31:0] f952_rdata;
  sr_buffer_32_1 f952(.wen(f952_wen), .wdata(f952_wdata), .clk(f952_clk), .rst(f952_rst), .rdata(f952_rdata));
  assign f952_clk = clk;
  assign f952_rst = rst;
  // Bindings to f952

  // f954
  logic [0:0] f954_wen;
  logic [31:0] f954_wdata;
  logic [0:0] f954_clk;
  logic [0:0] f954_rst;
  logic [31:0] f954_rdata;
  sr_buffer_32_1 f954(.wen(f954_wen), .wdata(f954_wdata), .clk(f954_clk), .rst(f954_rst), .rdata(f954_rdata));
  assign f954_clk = clk;
  assign f954_rst = rst;
  // Bindings to f954

  // f956
  logic [0:0] f956_wen;
  logic [31:0] f956_wdata;
  logic [0:0] f956_clk;
  logic [0:0] f956_rst;
  logic [31:0] f956_rdata;
  sr_buffer_32_1 f956(.wen(f956_wen), .wdata(f956_wdata), .clk(f956_clk), .rst(f956_rst), .rdata(f956_rdata));
  assign f956_clk = clk;
  assign f956_rst = rst;
  // Bindings to f956

  // f958
  logic [0:0] f958_wen;
  logic [31:0] f958_wdata;
  logic [0:0] f958_clk;
  logic [0:0] f958_rst;
  logic [31:0] f958_rdata;
  sr_buffer_32_1 f958(.wen(f958_wen), .wdata(f958_wdata), .clk(f958_clk), .rst(f958_rst), .rdata(f958_rdata));
  assign f958_clk = clk;
  assign f958_rst = rst;
  // Bindings to f958

  // f960
  logic [0:0] f960_wen;
  logic [31:0] f960_wdata;
  logic [0:0] f960_clk;
  logic [0:0] f960_rst;
  logic [31:0] f960_rdata;
  sr_buffer_32_1 f960(.wen(f960_wen), .wdata(f960_wdata), .clk(f960_clk), .rst(f960_rst), .rdata(f960_rdata));
  assign f960_clk = clk;
  assign f960_rst = rst;
  // Bindings to f960

  // f962
  logic [0:0] f962_wen;
  logic [31:0] f962_wdata;
  logic [0:0] f962_clk;
  logic [0:0] f962_rst;
  logic [31:0] f962_rdata;
  sr_buffer_32_1 f962(.wen(f962_wen), .wdata(f962_wdata), .clk(f962_clk), .rst(f962_rst), .rdata(f962_rdata));
  assign f962_clk = clk;
  assign f962_rst = rst;
  // Bindings to f962

  // f964
  logic [0:0] f964_wen;
  logic [31:0] f964_wdata;
  logic [0:0] f964_clk;
  logic [0:0] f964_rst;
  logic [31:0] f964_rdata;
  sr_buffer_32_1 f964(.wen(f964_wen), .wdata(f964_wdata), .clk(f964_clk), .rst(f964_rst), .rdata(f964_rdata));
  assign f964_clk = clk;
  assign f964_rst = rst;
  // Bindings to f964

  // f966
  logic [0:0] f966_wen;
  logic [31:0] f966_wdata;
  logic [0:0] f966_clk;
  logic [0:0] f966_rst;
  logic [31:0] f966_rdata;
  sr_buffer_32_1 f966(.wen(f966_wen), .wdata(f966_wdata), .clk(f966_clk), .rst(f966_rst), .rdata(f966_rdata));
  assign f966_clk = clk;
  assign f966_rst = rst;
  // Bindings to f966

  // f968
  logic [0:0] f968_wen;
  logic [31:0] f968_wdata;
  logic [0:0] f968_clk;
  logic [0:0] f968_rst;
  logic [31:0] f968_rdata;
  sr_buffer_32_1 f968(.wen(f968_wen), .wdata(f968_wdata), .clk(f968_clk), .rst(f968_rst), .rdata(f968_rdata));
  assign f968_clk = clk;
  assign f968_rst = rst;
  // Bindings to f968

  // f970
  logic [0:0] f970_wen;
  logic [31:0] f970_wdata;
  logic [0:0] f970_clk;
  logic [0:0] f970_rst;
  logic [31:0] f970_rdata;
  sr_buffer_32_1 f970(.wen(f970_wen), .wdata(f970_wdata), .clk(f970_clk), .rst(f970_rst), .rdata(f970_rdata));
  assign f970_clk = clk;
  assign f970_rst = rst;
  // Bindings to f970

  // f972
  logic [0:0] f972_wen;
  logic [31:0] f972_wdata;
  logic [0:0] f972_clk;
  logic [0:0] f972_rst;
  logic [31:0] f972_rdata;
  sr_buffer_32_1 f972(.wen(f972_wen), .wdata(f972_wdata), .clk(f972_clk), .rst(f972_rst), .rdata(f972_rdata));
  assign f972_clk = clk;
  assign f972_rst = rst;
  // Bindings to f972

  // f974
  logic [0:0] f974_wen;
  logic [31:0] f974_wdata;
  logic [0:0] f974_clk;
  logic [0:0] f974_rst;
  logic [31:0] f974_rdata;
  sr_buffer_32_1 f974(.wen(f974_wen), .wdata(f974_wdata), .clk(f974_clk), .rst(f974_rst), .rdata(f974_rdata));
  assign f974_clk = clk;
  assign f974_rst = rst;
  // Bindings to f974

  // f976
  logic [0:0] f976_wen;
  logic [31:0] f976_wdata;
  logic [0:0] f976_clk;
  logic [0:0] f976_rst;
  logic [31:0] f976_rdata;
  sr_buffer_32_1 f976(.wen(f976_wen), .wdata(f976_wdata), .clk(f976_clk), .rst(f976_rst), .rdata(f976_rdata));
  assign f976_clk = clk;
  assign f976_rst = rst;
  // Bindings to f976

  // f978
  logic [0:0] f978_wen;
  logic [31:0] f978_wdata;
  logic [0:0] f978_clk;
  logic [0:0] f978_rst;
  logic [31:0] f978_rdata;
  sr_buffer_32_1 f978(.wen(f978_wen), .wdata(f978_wdata), .clk(f978_clk), .rst(f978_rst), .rdata(f978_rdata));
  assign f978_clk = clk;
  assign f978_rst = rst;
  // Bindings to f978

  // f980
  logic [0:0] f980_wen;
  logic [31:0] f980_wdata;
  logic [0:0] f980_clk;
  logic [0:0] f980_rst;
  logic [31:0] f980_rdata;
  sr_buffer_32_1 f980(.wen(f980_wen), .wdata(f980_wdata), .clk(f980_clk), .rst(f980_rst), .rdata(f980_rdata));
  assign f980_clk = clk;
  assign f980_rst = rst;
  // Bindings to f980

  // f982
  logic [0:0] f982_wen;
  logic [31:0] f982_wdata;
  logic [0:0] f982_clk;
  logic [0:0] f982_rst;
  logic [31:0] f982_rdata;
  sr_buffer_32_1 f982(.wen(f982_wen), .wdata(f982_wdata), .clk(f982_clk), .rst(f982_rst), .rdata(f982_rdata));
  assign f982_clk = clk;
  assign f982_rst = rst;
  // Bindings to f982

  // f984
  logic [0:0] f984_wen;
  logic [31:0] f984_wdata;
  logic [0:0] f984_clk;
  logic [0:0] f984_rst;
  logic [31:0] f984_rdata;
  sr_buffer_32_1 f984(.wen(f984_wen), .wdata(f984_wdata), .clk(f984_clk), .rst(f984_rst), .rdata(f984_rdata));
  assign f984_clk = clk;
  assign f984_rst = rst;
  // Bindings to f984

  // f986
  logic [0:0] f986_wen;
  logic [31:0] f986_wdata;
  logic [0:0] f986_clk;
  logic [0:0] f986_rst;
  logic [31:0] f986_rdata;
  sr_buffer_32_1 f986(.wen(f986_wen), .wdata(f986_wdata), .clk(f986_clk), .rst(f986_rst), .rdata(f986_rdata));
  assign f986_clk = clk;
  assign f986_rst = rst;
  // Bindings to f986

  // f988
  logic [0:0] f988_wen;
  logic [31:0] f988_wdata;
  logic [0:0] f988_clk;
  logic [0:0] f988_rst;
  logic [31:0] f988_rdata;
  sr_buffer_32_1 f988(.wen(f988_wen), .wdata(f988_wdata), .clk(f988_clk), .rst(f988_rst), .rdata(f988_rdata));
  assign f988_clk = clk;
  assign f988_rst = rst;
  // Bindings to f988

  // f990
  logic [0:0] f990_wen;
  logic [31:0] f990_wdata;
  logic [0:0] f990_clk;
  logic [0:0] f990_rst;
  logic [31:0] f990_rdata;
  sr_buffer_32_1 f990(.wen(f990_wen), .wdata(f990_wdata), .clk(f990_clk), .rst(f990_rst), .rdata(f990_rdata));
  assign f990_clk = clk;
  assign f990_rst = rst;
  // Bindings to f990

  // f992
  logic [0:0] f992_wen;
  logic [31:0] f992_wdata;
  logic [0:0] f992_clk;
  logic [0:0] f992_rst;
  logic [31:0] f992_rdata;
  sr_buffer_32_1 f992(.wen(f992_wen), .wdata(f992_wdata), .clk(f992_clk), .rst(f992_rst), .rdata(f992_rdata));
  assign f992_clk = clk;
  assign f992_rst = rst;
  // Bindings to f992

  // f994
  logic [0:0] f994_wen;
  logic [31:0] f994_wdata;
  logic [0:0] f994_clk;
  logic [0:0] f994_rst;
  logic [31:0] f994_rdata;
  sr_buffer_32_1 f994(.wen(f994_wen), .wdata(f994_wdata), .clk(f994_clk), .rst(f994_rst), .rdata(f994_rdata));
  assign f994_clk = clk;
  assign f994_rst = rst;
  // Bindings to f994

  // f996
  logic [0:0] f996_wen;
  logic [31:0] f996_wdata;
  logic [0:0] f996_clk;
  logic [0:0] f996_rst;
  logic [31:0] f996_rdata;
  sr_buffer_32_1 f996(.wen(f996_wen), .wdata(f996_wdata), .clk(f996_clk), .rst(f996_rst), .rdata(f996_rdata));
  assign f996_clk = clk;
  assign f996_rst = rst;
  // Bindings to f996

  // f998
  logic [0:0] f998_wen;
  logic [31:0] f998_wdata;
  logic [0:0] f998_clk;
  logic [0:0] f998_rst;
  logic [31:0] f998_rdata;
  sr_buffer_32_1 f998(.wen(f998_wen), .wdata(f998_wdata), .clk(f998_clk), .rst(f998_rst), .rdata(f998_rdata));
  assign f998_clk = clk;
  assign f998_rst = rst;
  // Bindings to f998

  // f1000
  logic [0:0] f1000_wen;
  logic [31:0] f1000_wdata;
  logic [0:0] f1000_clk;
  logic [0:0] f1000_rst;
  logic [31:0] f1000_rdata;
  sr_buffer_32_1 f1000(.wen(f1000_wen), .wdata(f1000_wdata), .clk(f1000_clk), .rst(f1000_rst), .rdata(f1000_rdata));
  assign f1000_clk = clk;
  assign f1000_rst = rst;
  // Bindings to f1000

  // f1002
  logic [0:0] f1002_wen;
  logic [31:0] f1002_wdata;
  logic [0:0] f1002_clk;
  logic [0:0] f1002_rst;
  logic [31:0] f1002_rdata;
  sr_buffer_32_1 f1002(.wen(f1002_wen), .wdata(f1002_wdata), .clk(f1002_clk), .rst(f1002_rst), .rdata(f1002_rdata));
  assign f1002_clk = clk;
  assign f1002_rst = rst;
  // Bindings to f1002

  // f1004
  logic [0:0] f1004_wen;
  logic [31:0] f1004_wdata;
  logic [0:0] f1004_clk;
  logic [0:0] f1004_rst;
  logic [31:0] f1004_rdata;
  sr_buffer_32_1 f1004(.wen(f1004_wen), .wdata(f1004_wdata), .clk(f1004_clk), .rst(f1004_rst), .rdata(f1004_rdata));
  assign f1004_clk = clk;
  assign f1004_rst = rst;
  // Bindings to f1004

  // f1006
  logic [0:0] f1006_wen;
  logic [31:0] f1006_wdata;
  logic [0:0] f1006_clk;
  logic [0:0] f1006_rst;
  logic [31:0] f1006_rdata;
  sr_buffer_32_1 f1006(.wen(f1006_wen), .wdata(f1006_wdata), .clk(f1006_clk), .rst(f1006_rst), .rdata(f1006_rdata));
  assign f1006_clk = clk;
  assign f1006_rst = rst;
  // Bindings to f1006

  // f1008
  logic [0:0] f1008_wen;
  logic [31:0] f1008_wdata;
  logic [0:0] f1008_clk;
  logic [0:0] f1008_rst;
  logic [31:0] f1008_rdata;
  sr_buffer_32_1 f1008(.wen(f1008_wen), .wdata(f1008_wdata), .clk(f1008_clk), .rst(f1008_rst), .rdata(f1008_rdata));
  assign f1008_clk = clk;
  assign f1008_rst = rst;
  // Bindings to f1008

  // f1010
  logic [0:0] f1010_wen;
  logic [31:0] f1010_wdata;
  logic [0:0] f1010_clk;
  logic [0:0] f1010_rst;
  logic [31:0] f1010_rdata;
  sr_buffer_32_1 f1010(.wen(f1010_wen), .wdata(f1010_wdata), .clk(f1010_clk), .rst(f1010_rst), .rdata(f1010_rdata));
  assign f1010_clk = clk;
  assign f1010_rst = rst;
  // Bindings to f1010

  // f1012
  logic [0:0] f1012_wen;
  logic [31:0] f1012_wdata;
  logic [0:0] f1012_clk;
  logic [0:0] f1012_rst;
  logic [31:0] f1012_rdata;
  sr_buffer_32_1 f1012(.wen(f1012_wen), .wdata(f1012_wdata), .clk(f1012_clk), .rst(f1012_rst), .rdata(f1012_rdata));
  assign f1012_clk = clk;
  assign f1012_rst = rst;
  // Bindings to f1012

  // f1014
  logic [0:0] f1014_wen;
  logic [31:0] f1014_wdata;
  logic [0:0] f1014_clk;
  logic [0:0] f1014_rst;
  logic [31:0] f1014_rdata;
  sr_buffer_32_1 f1014(.wen(f1014_wen), .wdata(f1014_wdata), .clk(f1014_clk), .rst(f1014_rst), .rdata(f1014_rdata));
  assign f1014_clk = clk;
  assign f1014_rst = rst;
  // Bindings to f1014

  // f1016
  logic [0:0] f1016_wen;
  logic [31:0] f1016_wdata;
  logic [0:0] f1016_clk;
  logic [0:0] f1016_rst;
  logic [31:0] f1016_rdata;
  sr_buffer_32_1 f1016(.wen(f1016_wen), .wdata(f1016_wdata), .clk(f1016_clk), .rst(f1016_rst), .rdata(f1016_rdata));
  assign f1016_clk = clk;
  assign f1016_rst = rst;
  // Bindings to f1016

  // f1018
  logic [0:0] f1018_wen;
  logic [31:0] f1018_wdata;
  logic [0:0] f1018_clk;
  logic [0:0] f1018_rst;
  logic [31:0] f1018_rdata;
  sr_buffer_32_1 f1018(.wen(f1018_wen), .wdata(f1018_wdata), .clk(f1018_clk), .rst(f1018_rst), .rdata(f1018_rdata));
  assign f1018_clk = clk;
  assign f1018_rst = rst;
  // Bindings to f1018

  // f1020
  logic [0:0] f1020_wen;
  logic [31:0] f1020_wdata;
  logic [0:0] f1020_clk;
  logic [0:0] f1020_rst;
  logic [31:0] f1020_rdata;
  sr_buffer_32_1 f1020(.wen(f1020_wen), .wdata(f1020_wdata), .clk(f1020_clk), .rst(f1020_rst), .rdata(f1020_rdata));
  assign f1020_clk = clk;
  assign f1020_rst = rst;
  // Bindings to f1020

  // f1022
  logic [0:0] f1022_wen;
  logic [31:0] f1022_wdata;
  logic [0:0] f1022_clk;
  logic [0:0] f1022_rst;
  logic [31:0] f1022_rdata;
  sr_buffer_32_1 f1022(.wen(f1022_wen), .wdata(f1022_wdata), .clk(f1022_clk), .rst(f1022_rst), .rdata(f1022_rdata));
  assign f1022_clk = clk;
  assign f1022_rst = rst;
  // Bindings to f1022

  // f1024
  logic [0:0] f1024_wen;
  logic [31:0] f1024_wdata;
  logic [0:0] f1024_clk;
  logic [0:0] f1024_rst;
  logic [31:0] f1024_rdata;
  sr_buffer_32_1 f1024(.wen(f1024_wen), .wdata(f1024_wdata), .clk(f1024_clk), .rst(f1024_rst), .rdata(f1024_rdata));
  assign f1024_clk = clk;
  assign f1024_rst = rst;
  // Bindings to f1024

  // f1026
  logic [0:0] f1026_wen;
  logic [31:0] f1026_wdata;
  logic [0:0] f1026_clk;
  logic [0:0] f1026_rst;
  logic [31:0] f1026_rdata;
  sr_buffer_32_1 f1026(.wen(f1026_wen), .wdata(f1026_wdata), .clk(f1026_clk), .rst(f1026_rst), .rdata(f1026_rdata));
  assign f1026_clk = clk;
  assign f1026_rst = rst;
  // Bindings to f1026

  // f1028
  logic [0:0] f1028_wen;
  logic [31:0] f1028_wdata;
  logic [0:0] f1028_clk;
  logic [0:0] f1028_rst;
  logic [31:0] f1028_rdata;
  sr_buffer_32_1 f1028(.wen(f1028_wen), .wdata(f1028_wdata), .clk(f1028_clk), .rst(f1028_rst), .rdata(f1028_rdata));
  assign f1028_clk = clk;
  assign f1028_rst = rst;
  // Bindings to f1028

  // f1030
  logic [0:0] f1030_wen;
  logic [31:0] f1030_wdata;
  logic [0:0] f1030_clk;
  logic [0:0] f1030_rst;
  logic [31:0] f1030_rdata;
  sr_buffer_32_1 f1030(.wen(f1030_wen), .wdata(f1030_wdata), .clk(f1030_clk), .rst(f1030_rst), .rdata(f1030_rdata));
  assign f1030_clk = clk;
  assign f1030_rst = rst;
  // Bindings to f1030

  // f1032
  logic [0:0] f1032_wen;
  logic [31:0] f1032_wdata;
  logic [0:0] f1032_clk;
  logic [0:0] f1032_rst;
  logic [31:0] f1032_rdata;
  sr_buffer_32_1 f1032(.wen(f1032_wen), .wdata(f1032_wdata), .clk(f1032_clk), .rst(f1032_rst), .rdata(f1032_rdata));
  assign f1032_clk = clk;
  assign f1032_rst = rst;
  // Bindings to f1032

  // f1034
  logic [0:0] f1034_wen;
  logic [31:0] f1034_wdata;
  logic [0:0] f1034_clk;
  logic [0:0] f1034_rst;
  logic [31:0] f1034_rdata;
  sr_buffer_32_1 f1034(.wen(f1034_wen), .wdata(f1034_wdata), .clk(f1034_clk), .rst(f1034_rst), .rdata(f1034_rdata));
  assign f1034_clk = clk;
  assign f1034_rst = rst;
  // Bindings to f1034

  // f1036
  logic [0:0] f1036_wen;
  logic [31:0] f1036_wdata;
  logic [0:0] f1036_clk;
  logic [0:0] f1036_rst;
  logic [31:0] f1036_rdata;
  sr_buffer_32_1 f1036(.wen(f1036_wen), .wdata(f1036_wdata), .clk(f1036_clk), .rst(f1036_rst), .rdata(f1036_rdata));
  assign f1036_clk = clk;
  assign f1036_rst = rst;
  // Bindings to f1036

  // f1038
  logic [0:0] f1038_wen;
  logic [31:0] f1038_wdata;
  logic [0:0] f1038_clk;
  logic [0:0] f1038_rst;
  logic [31:0] f1038_rdata;
  sr_buffer_32_1 f1038(.wen(f1038_wen), .wdata(f1038_wdata), .clk(f1038_clk), .rst(f1038_rst), .rdata(f1038_rdata));
  assign f1038_clk = clk;
  assign f1038_rst = rst;
  // Bindings to f1038

  // f1040
  logic [0:0] f1040_wen;
  logic [31:0] f1040_wdata;
  logic [0:0] f1040_clk;
  logic [0:0] f1040_rst;
  logic [31:0] f1040_rdata;
  sr_buffer_32_1 f1040(.wen(f1040_wen), .wdata(f1040_wdata), .clk(f1040_clk), .rst(f1040_rst), .rdata(f1040_rdata));
  assign f1040_clk = clk;
  assign f1040_rst = rst;
  // Bindings to f1040

  // f1042
  logic [0:0] f1042_wen;
  logic [31:0] f1042_wdata;
  logic [0:0] f1042_clk;
  logic [0:0] f1042_rst;
  logic [31:0] f1042_rdata;
  sr_buffer_32_1 f1042(.wen(f1042_wen), .wdata(f1042_wdata), .clk(f1042_clk), .rst(f1042_rst), .rdata(f1042_rdata));
  assign f1042_clk = clk;
  assign f1042_rst = rst;
  // Bindings to f1042

  // f1044
  logic [0:0] f1044_wen;
  logic [31:0] f1044_wdata;
  logic [0:0] f1044_clk;
  logic [0:0] f1044_rst;
  logic [31:0] f1044_rdata;
  sr_buffer_32_1 f1044(.wen(f1044_wen), .wdata(f1044_wdata), .clk(f1044_clk), .rst(f1044_rst), .rdata(f1044_rdata));
  assign f1044_clk = clk;
  assign f1044_rst = rst;
  // Bindings to f1044

  // f1046
  logic [0:0] f1046_wen;
  logic [31:0] f1046_wdata;
  logic [0:0] f1046_clk;
  logic [0:0] f1046_rst;
  logic [31:0] f1046_rdata;
  sr_buffer_32_1 f1046(.wen(f1046_wen), .wdata(f1046_wdata), .clk(f1046_clk), .rst(f1046_rst), .rdata(f1046_rdata));
  assign f1046_clk = clk;
  assign f1046_rst = rst;
  // Bindings to f1046

  // f1048
  logic [0:0] f1048_wen;
  logic [31:0] f1048_wdata;
  logic [0:0] f1048_clk;
  logic [0:0] f1048_rst;
  logic [31:0] f1048_rdata;
  sr_buffer_32_1 f1048(.wen(f1048_wen), .wdata(f1048_wdata), .clk(f1048_clk), .rst(f1048_rst), .rdata(f1048_rdata));
  assign f1048_clk = clk;
  assign f1048_rst = rst;
  // Bindings to f1048

  // f1050
  logic [0:0] f1050_wen;
  logic [31:0] f1050_wdata;
  logic [0:0] f1050_clk;
  logic [0:0] f1050_rst;
  logic [31:0] f1050_rdata;
  sr_buffer_32_1 f1050(.wen(f1050_wen), .wdata(f1050_wdata), .clk(f1050_clk), .rst(f1050_rst), .rdata(f1050_rdata));
  assign f1050_clk = clk;
  assign f1050_rst = rst;
  // Bindings to f1050

  // f1052
  logic [0:0] f1052_wen;
  logic [31:0] f1052_wdata;
  logic [0:0] f1052_clk;
  logic [0:0] f1052_rst;
  logic [31:0] f1052_rdata;
  sr_buffer_32_1 f1052(.wen(f1052_wen), .wdata(f1052_wdata), .clk(f1052_clk), .rst(f1052_rst), .rdata(f1052_rdata));
  assign f1052_clk = clk;
  assign f1052_rst = rst;
  // Bindings to f1052

  // f1054
  logic [0:0] f1054_wen;
  logic [31:0] f1054_wdata;
  logic [0:0] f1054_clk;
  logic [0:0] f1054_rst;
  logic [31:0] f1054_rdata;
  sr_buffer_32_1 f1054(.wen(f1054_wen), .wdata(f1054_wdata), .clk(f1054_clk), .rst(f1054_rst), .rdata(f1054_rdata));
  assign f1054_clk = clk;
  assign f1054_rst = rst;
  // Bindings to f1054

  // f1056
  logic [0:0] f1056_wen;
  logic [31:0] f1056_wdata;
  logic [0:0] f1056_clk;
  logic [0:0] f1056_rst;
  logic [31:0] f1056_rdata;
  sr_buffer_32_1 f1056(.wen(f1056_wen), .wdata(f1056_wdata), .clk(f1056_clk), .rst(f1056_rst), .rdata(f1056_rdata));
  assign f1056_clk = clk;
  assign f1056_rst = rst;
  // Bindings to f1056

  // f1058
  logic [0:0] f1058_wen;
  logic [31:0] f1058_wdata;
  logic [0:0] f1058_clk;
  logic [0:0] f1058_rst;
  logic [31:0] f1058_rdata;
  sr_buffer_32_1 f1058(.wen(f1058_wen), .wdata(f1058_wdata), .clk(f1058_clk), .rst(f1058_rst), .rdata(f1058_rdata));
  assign f1058_clk = clk;
  assign f1058_rst = rst;
  // Bindings to f1058

  // f1060
  logic [0:0] f1060_wen;
  logic [31:0] f1060_wdata;
  logic [0:0] f1060_clk;
  logic [0:0] f1060_rst;
  logic [31:0] f1060_rdata;
  sr_buffer_32_1 f1060(.wen(f1060_wen), .wdata(f1060_wdata), .clk(f1060_clk), .rst(f1060_rst), .rdata(f1060_rdata));
  assign f1060_clk = clk;
  assign f1060_rst = rst;
  // Bindings to f1060

  // f1062
  logic [0:0] f1062_wen;
  logic [31:0] f1062_wdata;
  logic [0:0] f1062_clk;
  logic [0:0] f1062_rst;
  logic [31:0] f1062_rdata;
  sr_buffer_32_1 f1062(.wen(f1062_wen), .wdata(f1062_wdata), .clk(f1062_clk), .rst(f1062_rst), .rdata(f1062_rdata));
  assign f1062_clk = clk;
  assign f1062_rst = rst;
  // Bindings to f1062

  // f1064
  logic [0:0] f1064_wen;
  logic [31:0] f1064_wdata;
  logic [0:0] f1064_clk;
  logic [0:0] f1064_rst;
  logic [31:0] f1064_rdata;
  sr_buffer_32_1 f1064(.wen(f1064_wen), .wdata(f1064_wdata), .clk(f1064_clk), .rst(f1064_rst), .rdata(f1064_rdata));
  assign f1064_clk = clk;
  assign f1064_rst = rst;
  // Bindings to f1064

  // f1066
  logic [0:0] f1066_wen;
  logic [31:0] f1066_wdata;
  logic [0:0] f1066_clk;
  logic [0:0] f1066_rst;
  logic [31:0] f1066_rdata;
  sr_buffer_32_1 f1066(.wen(f1066_wen), .wdata(f1066_wdata), .clk(f1066_clk), .rst(f1066_rst), .rdata(f1066_rdata));
  assign f1066_clk = clk;
  assign f1066_rst = rst;
  // Bindings to f1066

  // f1068
  logic [0:0] f1068_wen;
  logic [31:0] f1068_wdata;
  logic [0:0] f1068_clk;
  logic [0:0] f1068_rst;
  logic [31:0] f1068_rdata;
  sr_buffer_32_1 f1068(.wen(f1068_wen), .wdata(f1068_wdata), .clk(f1068_clk), .rst(f1068_rst), .rdata(f1068_rdata));
  assign f1068_clk = clk;
  assign f1068_rst = rst;
  // Bindings to f1068

  // f1070
  logic [0:0] f1070_wen;
  logic [31:0] f1070_wdata;
  logic [0:0] f1070_clk;
  logic [0:0] f1070_rst;
  logic [31:0] f1070_rdata;
  sr_buffer_32_1 f1070(.wen(f1070_wen), .wdata(f1070_wdata), .clk(f1070_clk), .rst(f1070_rst), .rdata(f1070_rdata));
  assign f1070_clk = clk;
  assign f1070_rst = rst;
  // Bindings to f1070

  // f1072
  logic [0:0] f1072_wen;
  logic [31:0] f1072_wdata;
  logic [0:0] f1072_clk;
  logic [0:0] f1072_rst;
  logic [31:0] f1072_rdata;
  sr_buffer_32_1 f1072(.wen(f1072_wen), .wdata(f1072_wdata), .clk(f1072_clk), .rst(f1072_rst), .rdata(f1072_rdata));
  assign f1072_clk = clk;
  assign f1072_rst = rst;
  // Bindings to f1072

  // f1074
  logic [0:0] f1074_wen;
  logic [31:0] f1074_wdata;
  logic [0:0] f1074_clk;
  logic [0:0] f1074_rst;
  logic [31:0] f1074_rdata;
  sr_buffer_32_1 f1074(.wen(f1074_wen), .wdata(f1074_wdata), .clk(f1074_clk), .rst(f1074_rst), .rdata(f1074_rdata));
  assign f1074_clk = clk;
  assign f1074_rst = rst;
  // Bindings to f1074

  // f1076
  logic [0:0] f1076_wen;
  logic [31:0] f1076_wdata;
  logic [0:0] f1076_clk;
  logic [0:0] f1076_rst;
  logic [31:0] f1076_rdata;
  sr_buffer_32_1 f1076(.wen(f1076_wen), .wdata(f1076_wdata), .clk(f1076_clk), .rst(f1076_rst), .rdata(f1076_rdata));
  assign f1076_clk = clk;
  assign f1076_rst = rst;
  // Bindings to f1076

  // f1078
  logic [0:0] f1078_wen;
  logic [31:0] f1078_wdata;
  logic [0:0] f1078_clk;
  logic [0:0] f1078_rst;
  logic [31:0] f1078_rdata;
  sr_buffer_32_1 f1078(.wen(f1078_wen), .wdata(f1078_wdata), .clk(f1078_clk), .rst(f1078_rst), .rdata(f1078_rdata));
  assign f1078_clk = clk;
  assign f1078_rst = rst;
  // Bindings to f1078

  // f1080
  logic [0:0] f1080_wen;
  logic [31:0] f1080_wdata;
  logic [0:0] f1080_clk;
  logic [0:0] f1080_rst;
  logic [31:0] f1080_rdata;
  sr_buffer_32_1 f1080(.wen(f1080_wen), .wdata(f1080_wdata), .clk(f1080_clk), .rst(f1080_rst), .rdata(f1080_rdata));
  assign f1080_clk = clk;
  assign f1080_rst = rst;
  // Bindings to f1080

  // f1082
  logic [0:0] f1082_wen;
  logic [31:0] f1082_wdata;
  logic [0:0] f1082_clk;
  logic [0:0] f1082_rst;
  logic [31:0] f1082_rdata;
  sr_buffer_32_1 f1082(.wen(f1082_wen), .wdata(f1082_wdata), .clk(f1082_clk), .rst(f1082_rst), .rdata(f1082_rdata));
  assign f1082_clk = clk;
  assign f1082_rst = rst;
  // Bindings to f1082

  // f1084
  logic [0:0] f1084_wen;
  logic [31:0] f1084_wdata;
  logic [0:0] f1084_clk;
  logic [0:0] f1084_rst;
  logic [31:0] f1084_rdata;
  sr_buffer_32_1 f1084(.wen(f1084_wen), .wdata(f1084_wdata), .clk(f1084_clk), .rst(f1084_rst), .rdata(f1084_rdata));
  assign f1084_clk = clk;
  assign f1084_rst = rst;
  // Bindings to f1084

  // f1086
  logic [0:0] f1086_wen;
  logic [31:0] f1086_wdata;
  logic [0:0] f1086_clk;
  logic [0:0] f1086_rst;
  logic [31:0] f1086_rdata;
  sr_buffer_32_1 f1086(.wen(f1086_wen), .wdata(f1086_wdata), .clk(f1086_clk), .rst(f1086_rst), .rdata(f1086_rdata));
  assign f1086_clk = clk;
  assign f1086_rst = rst;
  // Bindings to f1086

  // f1088
  logic [0:0] f1088_wen;
  logic [31:0] f1088_wdata;
  logic [0:0] f1088_clk;
  logic [0:0] f1088_rst;
  logic [31:0] f1088_rdata;
  sr_buffer_32_1 f1088(.wen(f1088_wen), .wdata(f1088_wdata), .clk(f1088_clk), .rst(f1088_rst), .rdata(f1088_rdata));
  assign f1088_clk = clk;
  assign f1088_rst = rst;
  // Bindings to f1088

  // f1090
  logic [0:0] f1090_wen;
  logic [31:0] f1090_wdata;
  logic [0:0] f1090_clk;
  logic [0:0] f1090_rst;
  logic [31:0] f1090_rdata;
  sr_buffer_32_1 f1090(.wen(f1090_wen), .wdata(f1090_wdata), .clk(f1090_clk), .rst(f1090_rst), .rdata(f1090_rdata));
  assign f1090_clk = clk;
  assign f1090_rst = rst;
  // Bindings to f1090

  // f1092
  logic [0:0] f1092_wen;
  logic [31:0] f1092_wdata;
  logic [0:0] f1092_clk;
  logic [0:0] f1092_rst;
  logic [31:0] f1092_rdata;
  sr_buffer_32_1 f1092(.wen(f1092_wen), .wdata(f1092_wdata), .clk(f1092_clk), .rst(f1092_rst), .rdata(f1092_rdata));
  assign f1092_clk = clk;
  assign f1092_rst = rst;
  // Bindings to f1092

  // f1094
  logic [0:0] f1094_wen;
  logic [31:0] f1094_wdata;
  logic [0:0] f1094_clk;
  logic [0:0] f1094_rst;
  logic [31:0] f1094_rdata;
  sr_buffer_32_1 f1094(.wen(f1094_wen), .wdata(f1094_wdata), .clk(f1094_clk), .rst(f1094_rst), .rdata(f1094_rdata));
  assign f1094_clk = clk;
  assign f1094_rst = rst;
  // Bindings to f1094

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f1096
  logic [0:0] f1096_wen;
  logic [31:0] f1096_wdata;
  logic [0:0] f1096_clk;
  logic [0:0] f1096_rst;
  logic [31:0] f1096_rdata;
  sr_buffer_32_1 f1096(.wen(f1096_wen), .wdata(f1096_wdata), .clk(f1096_clk), .rst(f1096_rst), .rdata(f1096_rdata));
  assign f1096_clk = clk;
  assign f1096_rst = rst;
  // Bindings to f1096

  // f1098
  logic [0:0] f1098_wen;
  logic [31:0] f1098_wdata;
  logic [0:0] f1098_clk;
  logic [0:0] f1098_rst;
  logic [31:0] f1098_rdata;
  sr_buffer_32_1 f1098(.wen(f1098_wen), .wdata(f1098_wdata), .clk(f1098_clk), .rst(f1098_rst), .rdata(f1098_rdata));
  assign f1098_clk = clk;
  assign f1098_rst = rst;
  // Bindings to f1098

  // f1100
  logic [0:0] f1100_wen;
  logic [31:0] f1100_wdata;
  logic [0:0] f1100_clk;
  logic [0:0] f1100_rst;
  logic [31:0] f1100_rdata;
  sr_buffer_32_1 f1100(.wen(f1100_wen), .wdata(f1100_wdata), .clk(f1100_clk), .rst(f1100_rst), .rdata(f1100_rdata));
  assign f1100_clk = clk;
  assign f1100_rst = rst;
  // Bindings to f1100

  // f1102
  logic [0:0] f1102_wen;
  logic [31:0] f1102_wdata;
  logic [0:0] f1102_clk;
  logic [0:0] f1102_rst;
  logic [31:0] f1102_rdata;
  sr_buffer_32_1 f1102(.wen(f1102_wen), .wdata(f1102_wdata), .clk(f1102_clk), .rst(f1102_rst), .rdata(f1102_rdata));
  assign f1102_clk = clk;
  assign f1102_rst = rst;
  // Bindings to f1102

  // f1104
  logic [0:0] f1104_wen;
  logic [31:0] f1104_wdata;
  logic [0:0] f1104_clk;
  logic [0:0] f1104_rst;
  logic [31:0] f1104_rdata;
  sr_buffer_32_1 f1104(.wen(f1104_wen), .wdata(f1104_wdata), .clk(f1104_clk), .rst(f1104_rst), .rdata(f1104_rdata));
  assign f1104_clk = clk;
  assign f1104_rst = rst;
  // Bindings to f1104

  // f1106
  logic [0:0] f1106_wen;
  logic [31:0] f1106_wdata;
  logic [0:0] f1106_clk;
  logic [0:0] f1106_rst;
  logic [31:0] f1106_rdata;
  sr_buffer_32_1 f1106(.wen(f1106_wen), .wdata(f1106_wdata), .clk(f1106_clk), .rst(f1106_rst), .rdata(f1106_rdata));
  assign f1106_clk = clk;
  assign f1106_rst = rst;
  // Bindings to f1106

  // f1108
  logic [0:0] f1108_wen;
  logic [31:0] f1108_wdata;
  logic [0:0] f1108_clk;
  logic [0:0] f1108_rst;
  logic [31:0] f1108_rdata;
  sr_buffer_32_1 f1108(.wen(f1108_wen), .wdata(f1108_wdata), .clk(f1108_clk), .rst(f1108_rst), .rdata(f1108_rdata));
  assign f1108_clk = clk;
  assign f1108_rst = rst;
  // Bindings to f1108

  // f1110
  logic [0:0] f1110_wen;
  logic [31:0] f1110_wdata;
  logic [0:0] f1110_clk;
  logic [0:0] f1110_rst;
  logic [31:0] f1110_rdata;
  sr_buffer_32_1 f1110(.wen(f1110_wen), .wdata(f1110_wdata), .clk(f1110_clk), .rst(f1110_rst), .rdata(f1110_rdata));
  assign f1110_clk = clk;
  assign f1110_rst = rst;
  // Bindings to f1110

  // f1112
  logic [0:0] f1112_wen;
  logic [31:0] f1112_wdata;
  logic [0:0] f1112_clk;
  logic [0:0] f1112_rst;
  logic [31:0] f1112_rdata;
  sr_buffer_32_1 f1112(.wen(f1112_wen), .wdata(f1112_wdata), .clk(f1112_clk), .rst(f1112_rst), .rdata(f1112_rdata));
  assign f1112_clk = clk;
  assign f1112_rst = rst;
  // Bindings to f1112

  // f1114
  logic [0:0] f1114_wen;
  logic [31:0] f1114_wdata;
  logic [0:0] f1114_clk;
  logic [0:0] f1114_rst;
  logic [31:0] f1114_rdata;
  sr_buffer_32_1 f1114(.wen(f1114_wen), .wdata(f1114_wdata), .clk(f1114_clk), .rst(f1114_rst), .rdata(f1114_rdata));
  assign f1114_clk = clk;
  assign f1114_rst = rst;
  // Bindings to f1114

  // f1116
  logic [0:0] f1116_wen;
  logic [31:0] f1116_wdata;
  logic [0:0] f1116_clk;
  logic [0:0] f1116_rst;
  logic [31:0] f1116_rdata;
  sr_buffer_32_1 f1116(.wen(f1116_wen), .wdata(f1116_wdata), .clk(f1116_clk), .rst(f1116_rst), .rdata(f1116_rdata));
  assign f1116_clk = clk;
  assign f1116_rst = rst;
  // Bindings to f1116

  // f1118
  logic [0:0] f1118_wen;
  logic [31:0] f1118_wdata;
  logic [0:0] f1118_clk;
  logic [0:0] f1118_rst;
  logic [31:0] f1118_rdata;
  sr_buffer_32_1 f1118(.wen(f1118_wen), .wdata(f1118_wdata), .clk(f1118_clk), .rst(f1118_rst), .rdata(f1118_rdata));
  assign f1118_clk = clk;
  assign f1118_rst = rst;
  // Bindings to f1118

  // f1120
  logic [0:0] f1120_wen;
  logic [31:0] f1120_wdata;
  logic [0:0] f1120_clk;
  logic [0:0] f1120_rst;
  logic [31:0] f1120_rdata;
  sr_buffer_32_1 f1120(.wen(f1120_wen), .wdata(f1120_wdata), .clk(f1120_clk), .rst(f1120_rst), .rdata(f1120_rdata));
  assign f1120_clk = clk;
  assign f1120_rst = rst;
  // Bindings to f1120

  // f1122
  logic [0:0] f1122_wen;
  logic [31:0] f1122_wdata;
  logic [0:0] f1122_clk;
  logic [0:0] f1122_rst;
  logic [31:0] f1122_rdata;
  sr_buffer_32_1 f1122(.wen(f1122_wen), .wdata(f1122_wdata), .clk(f1122_clk), .rst(f1122_rst), .rdata(f1122_rdata));
  assign f1122_clk = clk;
  assign f1122_rst = rst;
  // Bindings to f1122

  // f1124
  logic [0:0] f1124_wen;
  logic [31:0] f1124_wdata;
  logic [0:0] f1124_clk;
  logic [0:0] f1124_rst;
  logic [31:0] f1124_rdata;
  sr_buffer_32_1 f1124(.wen(f1124_wen), .wdata(f1124_wdata), .clk(f1124_clk), .rst(f1124_rst), .rdata(f1124_rdata));
  assign f1124_clk = clk;
  assign f1124_rst = rst;
  // Bindings to f1124

  // f1126
  logic [0:0] f1126_wen;
  logic [31:0] f1126_wdata;
  logic [0:0] f1126_clk;
  logic [0:0] f1126_rst;
  logic [31:0] f1126_rdata;
  sr_buffer_32_1 f1126(.wen(f1126_wen), .wdata(f1126_wdata), .clk(f1126_clk), .rst(f1126_rst), .rdata(f1126_rdata));
  assign f1126_clk = clk;
  assign f1126_rst = rst;
  // Bindings to f1126

  // f1128
  logic [0:0] f1128_wen;
  logic [31:0] f1128_wdata;
  logic [0:0] f1128_clk;
  logic [0:0] f1128_rst;
  logic [31:0] f1128_rdata;
  sr_buffer_32_1 f1128(.wen(f1128_wen), .wdata(f1128_wdata), .clk(f1128_clk), .rst(f1128_rst), .rdata(f1128_rdata));
  assign f1128_clk = clk;
  assign f1128_rst = rst;
  // Bindings to f1128

  // f1130
  logic [0:0] f1130_wen;
  logic [31:0] f1130_wdata;
  logic [0:0] f1130_clk;
  logic [0:0] f1130_rst;
  logic [31:0] f1130_rdata;
  sr_buffer_32_1 f1130(.wen(f1130_wen), .wdata(f1130_wdata), .clk(f1130_clk), .rst(f1130_rst), .rdata(f1130_rdata));
  assign f1130_clk = clk;
  assign f1130_rst = rst;
  // Bindings to f1130

  // f1132
  logic [0:0] f1132_wen;
  logic [31:0] f1132_wdata;
  logic [0:0] f1132_clk;
  logic [0:0] f1132_rst;
  logic [31:0] f1132_rdata;
  sr_buffer_32_1 f1132(.wen(f1132_wen), .wdata(f1132_wdata), .clk(f1132_clk), .rst(f1132_rst), .rdata(f1132_rdata));
  assign f1132_clk = clk;
  assign f1132_rst = rst;
  // Bindings to f1132

  // f1134
  logic [0:0] f1134_wen;
  logic [31:0] f1134_wdata;
  logic [0:0] f1134_clk;
  logic [0:0] f1134_rst;
  logic [31:0] f1134_rdata;
  sr_buffer_32_1 f1134(.wen(f1134_wen), .wdata(f1134_wdata), .clk(f1134_clk), .rst(f1134_rst), .rdata(f1134_rdata));
  assign f1134_clk = clk;
  assign f1134_rst = rst;
  // Bindings to f1134

  // f1136
  logic [0:0] f1136_wen;
  logic [31:0] f1136_wdata;
  logic [0:0] f1136_clk;
  logic [0:0] f1136_rst;
  logic [31:0] f1136_rdata;
  sr_buffer_32_1 f1136(.wen(f1136_wen), .wdata(f1136_wdata), .clk(f1136_clk), .rst(f1136_rst), .rdata(f1136_rdata));
  assign f1136_clk = clk;
  assign f1136_rst = rst;
  // Bindings to f1136

  // f1138
  logic [0:0] f1138_wen;
  logic [31:0] f1138_wdata;
  logic [0:0] f1138_clk;
  logic [0:0] f1138_rst;
  logic [31:0] f1138_rdata;
  sr_buffer_32_1 f1138(.wen(f1138_wen), .wdata(f1138_wdata), .clk(f1138_clk), .rst(f1138_rst), .rdata(f1138_rdata));
  assign f1138_clk = clk;
  assign f1138_rst = rst;
  // Bindings to f1138

  // f1140
  logic [0:0] f1140_wen;
  logic [31:0] f1140_wdata;
  logic [0:0] f1140_clk;
  logic [0:0] f1140_rst;
  logic [31:0] f1140_rdata;
  sr_buffer_32_1 f1140(.wen(f1140_wen), .wdata(f1140_wdata), .clk(f1140_clk), .rst(f1140_rst), .rdata(f1140_rdata));
  assign f1140_clk = clk;
  assign f1140_rst = rst;
  // Bindings to f1140

  // f1142
  logic [0:0] f1142_wen;
  logic [31:0] f1142_wdata;
  logic [0:0] f1142_clk;
  logic [0:0] f1142_rst;
  logic [31:0] f1142_rdata;
  sr_buffer_32_1 f1142(.wen(f1142_wen), .wdata(f1142_wdata), .clk(f1142_clk), .rst(f1142_rst), .rdata(f1142_rdata));
  assign f1142_clk = clk;
  assign f1142_rst = rst;
  // Bindings to f1142

  // f1144
  logic [0:0] f1144_wen;
  logic [31:0] f1144_wdata;
  logic [0:0] f1144_clk;
  logic [0:0] f1144_rst;
  logic [31:0] f1144_rdata;
  sr_buffer_32_1 f1144(.wen(f1144_wen), .wdata(f1144_wdata), .clk(f1144_clk), .rst(f1144_rst), .rdata(f1144_rdata));
  assign f1144_clk = clk;
  assign f1144_rst = rst;
  // Bindings to f1144

  // f1146
  logic [0:0] f1146_wen;
  logic [31:0] f1146_wdata;
  logic [0:0] f1146_clk;
  logic [0:0] f1146_rst;
  logic [31:0] f1146_rdata;
  sr_buffer_32_1 f1146(.wen(f1146_wen), .wdata(f1146_wdata), .clk(f1146_clk), .rst(f1146_rst), .rdata(f1146_rdata));
  assign f1146_clk = clk;
  assign f1146_rst = rst;
  // Bindings to f1146

  // f1148
  logic [0:0] f1148_wen;
  logic [31:0] f1148_wdata;
  logic [0:0] f1148_clk;
  logic [0:0] f1148_rst;
  logic [31:0] f1148_rdata;
  sr_buffer_32_1 f1148(.wen(f1148_wen), .wdata(f1148_wdata), .clk(f1148_clk), .rst(f1148_rst), .rdata(f1148_rdata));
  assign f1148_clk = clk;
  assign f1148_rst = rst;
  // Bindings to f1148

  // f1150
  logic [0:0] f1150_wen;
  logic [31:0] f1150_wdata;
  logic [0:0] f1150_clk;
  logic [0:0] f1150_rst;
  logic [31:0] f1150_rdata;
  sr_buffer_32_1 f1150(.wen(f1150_wen), .wdata(f1150_wdata), .clk(f1150_clk), .rst(f1150_rst), .rdata(f1150_rdata));
  assign f1150_clk = clk;
  assign f1150_rst = rst;
  // Bindings to f1150

  // f1152
  logic [0:0] f1152_wen;
  logic [31:0] f1152_wdata;
  logic [0:0] f1152_clk;
  logic [0:0] f1152_rst;
  logic [31:0] f1152_rdata;
  sr_buffer_32_1 f1152(.wen(f1152_wen), .wdata(f1152_wdata), .clk(f1152_clk), .rst(f1152_rst), .rdata(f1152_rdata));
  assign f1152_clk = clk;
  assign f1152_rst = rst;
  // Bindings to f1152

  // f1154
  logic [0:0] f1154_wen;
  logic [31:0] f1154_wdata;
  logic [0:0] f1154_clk;
  logic [0:0] f1154_rst;
  logic [31:0] f1154_rdata;
  sr_buffer_32_1 f1154(.wen(f1154_wen), .wdata(f1154_wdata), .clk(f1154_clk), .rst(f1154_rst), .rdata(f1154_rdata));
  assign f1154_clk = clk;
  assign f1154_rst = rst;
  // Bindings to f1154

  // f1156
  logic [0:0] f1156_wen;
  logic [31:0] f1156_wdata;
  logic [0:0] f1156_clk;
  logic [0:0] f1156_rst;
  logic [31:0] f1156_rdata;
  sr_buffer_32_1 f1156(.wen(f1156_wen), .wdata(f1156_wdata), .clk(f1156_clk), .rst(f1156_rst), .rdata(f1156_rdata));
  assign f1156_clk = clk;
  assign f1156_rst = rst;
  // Bindings to f1156

  // f1158
  logic [0:0] f1158_wen;
  logic [31:0] f1158_wdata;
  logic [0:0] f1158_clk;
  logic [0:0] f1158_rst;
  logic [31:0] f1158_rdata;
  sr_buffer_32_1 f1158(.wen(f1158_wen), .wdata(f1158_wdata), .clk(f1158_clk), .rst(f1158_rst), .rdata(f1158_rdata));
  assign f1158_clk = clk;
  assign f1158_rst = rst;
  // Bindings to f1158

  // f1160
  logic [0:0] f1160_wen;
  logic [31:0] f1160_wdata;
  logic [0:0] f1160_clk;
  logic [0:0] f1160_rst;
  logic [31:0] f1160_rdata;
  sr_buffer_32_1 f1160(.wen(f1160_wen), .wdata(f1160_wdata), .clk(f1160_clk), .rst(f1160_rst), .rdata(f1160_rdata));
  assign f1160_clk = clk;
  assign f1160_rst = rst;
  // Bindings to f1160

  // f1162
  logic [0:0] f1162_wen;
  logic [31:0] f1162_wdata;
  logic [0:0] f1162_clk;
  logic [0:0] f1162_rst;
  logic [31:0] f1162_rdata;
  sr_buffer_32_1 f1162(.wen(f1162_wen), .wdata(f1162_wdata), .clk(f1162_clk), .rst(f1162_rst), .rdata(f1162_rdata));
  assign f1162_clk = clk;
  assign f1162_rst = rst;
  // Bindings to f1162

  // f1164
  logic [0:0] f1164_wen;
  logic [31:0] f1164_wdata;
  logic [0:0] f1164_clk;
  logic [0:0] f1164_rst;
  logic [31:0] f1164_rdata;
  sr_buffer_32_1 f1164(.wen(f1164_wen), .wdata(f1164_wdata), .clk(f1164_clk), .rst(f1164_rst), .rdata(f1164_rdata));
  assign f1164_clk = clk;
  assign f1164_rst = rst;
  // Bindings to f1164

  // f1166
  logic [0:0] f1166_wen;
  logic [31:0] f1166_wdata;
  logic [0:0] f1166_clk;
  logic [0:0] f1166_rst;
  logic [31:0] f1166_rdata;
  sr_buffer_32_1 f1166(.wen(f1166_wen), .wdata(f1166_wdata), .clk(f1166_clk), .rst(f1166_rst), .rdata(f1166_rdata));
  assign f1166_clk = clk;
  assign f1166_rst = rst;
  // Bindings to f1166

  // f1168
  logic [0:0] f1168_wen;
  logic [31:0] f1168_wdata;
  logic [0:0] f1168_clk;
  logic [0:0] f1168_rst;
  logic [31:0] f1168_rdata;
  sr_buffer_32_1 f1168(.wen(f1168_wen), .wdata(f1168_wdata), .clk(f1168_clk), .rst(f1168_rst), .rdata(f1168_rdata));
  assign f1168_clk = clk;
  assign f1168_rst = rst;
  // Bindings to f1168

  // f1170
  logic [0:0] f1170_wen;
  logic [31:0] f1170_wdata;
  logic [0:0] f1170_clk;
  logic [0:0] f1170_rst;
  logic [31:0] f1170_rdata;
  sr_buffer_32_1 f1170(.wen(f1170_wen), .wdata(f1170_wdata), .clk(f1170_clk), .rst(f1170_rst), .rdata(f1170_rdata));
  assign f1170_clk = clk;
  assign f1170_rst = rst;
  // Bindings to f1170

  // f1172
  logic [0:0] f1172_wen;
  logic [31:0] f1172_wdata;
  logic [0:0] f1172_clk;
  logic [0:0] f1172_rst;
  logic [31:0] f1172_rdata;
  sr_buffer_32_1 f1172(.wen(f1172_wen), .wdata(f1172_wdata), .clk(f1172_clk), .rst(f1172_rst), .rdata(f1172_rdata));
  assign f1172_clk = clk;
  assign f1172_rst = rst;
  // Bindings to f1172

  // f1174
  logic [0:0] f1174_wen;
  logic [31:0] f1174_wdata;
  logic [0:0] f1174_clk;
  logic [0:0] f1174_rst;
  logic [31:0] f1174_rdata;
  sr_buffer_32_1 f1174(.wen(f1174_wen), .wdata(f1174_wdata), .clk(f1174_clk), .rst(f1174_rst), .rdata(f1174_rdata));
  assign f1174_clk = clk;
  assign f1174_rst = rst;
  // Bindings to f1174

  // f1176
  logic [0:0] f1176_wen;
  logic [31:0] f1176_wdata;
  logic [0:0] f1176_clk;
  logic [0:0] f1176_rst;
  logic [31:0] f1176_rdata;
  sr_buffer_32_1 f1176(.wen(f1176_wen), .wdata(f1176_wdata), .clk(f1176_clk), .rst(f1176_rst), .rdata(f1176_rdata));
  assign f1176_clk = clk;
  assign f1176_rst = rst;
  // Bindings to f1176

  // f1178
  logic [0:0] f1178_wen;
  logic [31:0] f1178_wdata;
  logic [0:0] f1178_clk;
  logic [0:0] f1178_rst;
  logic [31:0] f1178_rdata;
  sr_buffer_32_1 f1178(.wen(f1178_wen), .wdata(f1178_wdata), .clk(f1178_clk), .rst(f1178_rst), .rdata(f1178_rdata));
  assign f1178_clk = clk;
  assign f1178_rst = rst;
  // Bindings to f1178

  // f1180
  logic [0:0] f1180_wen;
  logic [31:0] f1180_wdata;
  logic [0:0] f1180_clk;
  logic [0:0] f1180_rst;
  logic [31:0] f1180_rdata;
  sr_buffer_32_1 f1180(.wen(f1180_wen), .wdata(f1180_wdata), .clk(f1180_clk), .rst(f1180_rst), .rdata(f1180_rdata));
  assign f1180_clk = clk;
  assign f1180_rst = rst;
  // Bindings to f1180

  // f1182
  logic [0:0] f1182_wen;
  logic [31:0] f1182_wdata;
  logic [0:0] f1182_clk;
  logic [0:0] f1182_rst;
  logic [31:0] f1182_rdata;
  sr_buffer_32_1 f1182(.wen(f1182_wen), .wdata(f1182_wdata), .clk(f1182_clk), .rst(f1182_rst), .rdata(f1182_rdata));
  assign f1182_clk = clk;
  assign f1182_rst = rst;
  // Bindings to f1182

  // f1184
  logic [0:0] f1184_wen;
  logic [31:0] f1184_wdata;
  logic [0:0] f1184_clk;
  logic [0:0] f1184_rst;
  logic [31:0] f1184_rdata;
  sr_buffer_32_1 f1184(.wen(f1184_wen), .wdata(f1184_wdata), .clk(f1184_clk), .rst(f1184_rst), .rdata(f1184_rdata));
  assign f1184_clk = clk;
  assign f1184_rst = rst;
  // Bindings to f1184

  // f1186
  logic [0:0] f1186_wen;
  logic [31:0] f1186_wdata;
  logic [0:0] f1186_clk;
  logic [0:0] f1186_rst;
  logic [31:0] f1186_rdata;
  sr_buffer_32_1 f1186(.wen(f1186_wen), .wdata(f1186_wdata), .clk(f1186_clk), .rst(f1186_rst), .rdata(f1186_rdata));
  assign f1186_clk = clk;
  assign f1186_rst = rst;
  // Bindings to f1186

  // f1188
  logic [0:0] f1188_wen;
  logic [31:0] f1188_wdata;
  logic [0:0] f1188_clk;
  logic [0:0] f1188_rst;
  logic [31:0] f1188_rdata;
  sr_buffer_32_1 f1188(.wen(f1188_wen), .wdata(f1188_wdata), .clk(f1188_clk), .rst(f1188_rst), .rdata(f1188_rdata));
  assign f1188_clk = clk;
  assign f1188_rst = rst;
  // Bindings to f1188

  // f1190
  logic [0:0] f1190_wen;
  logic [31:0] f1190_wdata;
  logic [0:0] f1190_clk;
  logic [0:0] f1190_rst;
  logic [31:0] f1190_rdata;
  sr_buffer_32_1 f1190(.wen(f1190_wen), .wdata(f1190_wdata), .clk(f1190_clk), .rst(f1190_rst), .rdata(f1190_rdata));
  assign f1190_clk = clk;
  assign f1190_rst = rst;
  // Bindings to f1190

  // f1192
  logic [0:0] f1192_wen;
  logic [31:0] f1192_wdata;
  logic [0:0] f1192_clk;
  logic [0:0] f1192_rst;
  logic [31:0] f1192_rdata;
  sr_buffer_32_1 f1192(.wen(f1192_wen), .wdata(f1192_wdata), .clk(f1192_clk), .rst(f1192_rst), .rdata(f1192_rdata));
  assign f1192_clk = clk;
  assign f1192_rst = rst;
  // Bindings to f1192

  // f1194
  logic [0:0] f1194_wen;
  logic [31:0] f1194_wdata;
  logic [0:0] f1194_clk;
  logic [0:0] f1194_rst;
  logic [31:0] f1194_rdata;
  sr_buffer_32_1 f1194(.wen(f1194_wen), .wdata(f1194_wdata), .clk(f1194_clk), .rst(f1194_rst), .rdata(f1194_rdata));
  assign f1194_clk = clk;
  assign f1194_rst = rst;
  // Bindings to f1194

  // f1196
  logic [0:0] f1196_wen;
  logic [31:0] f1196_wdata;
  logic [0:0] f1196_clk;
  logic [0:0] f1196_rst;
  logic [31:0] f1196_rdata;
  sr_buffer_32_1 f1196(.wen(f1196_wen), .wdata(f1196_wdata), .clk(f1196_clk), .rst(f1196_rst), .rdata(f1196_rdata));
  assign f1196_clk = clk;
  assign f1196_rst = rst;
  // Bindings to f1196

  // f1198
  logic [0:0] f1198_wen;
  logic [31:0] f1198_wdata;
  logic [0:0] f1198_clk;
  logic [0:0] f1198_rst;
  logic [31:0] f1198_rdata;
  sr_buffer_32_1 f1198(.wen(f1198_wen), .wdata(f1198_wdata), .clk(f1198_clk), .rst(f1198_rst), .rdata(f1198_rdata));
  assign f1198_clk = clk;
  assign f1198_rst = rst;
  // Bindings to f1198

  // f1200
  logic [0:0] f1200_wen;
  logic [31:0] f1200_wdata;
  logic [0:0] f1200_clk;
  logic [0:0] f1200_rst;
  logic [31:0] f1200_rdata;
  sr_buffer_32_1 f1200(.wen(f1200_wen), .wdata(f1200_wdata), .clk(f1200_clk), .rst(f1200_rst), .rdata(f1200_rdata));
  assign f1200_clk = clk;
  assign f1200_rst = rst;
  // Bindings to f1200

  // f1202
  logic [0:0] f1202_wen;
  logic [31:0] f1202_wdata;
  logic [0:0] f1202_clk;
  logic [0:0] f1202_rst;
  logic [31:0] f1202_rdata;
  sr_buffer_32_1 f1202(.wen(f1202_wen), .wdata(f1202_wdata), .clk(f1202_clk), .rst(f1202_rst), .rdata(f1202_rdata));
  assign f1202_clk = clk;
  assign f1202_rst = rst;
  // Bindings to f1202

  // f1204
  logic [0:0] f1204_wen;
  logic [31:0] f1204_wdata;
  logic [0:0] f1204_clk;
  logic [0:0] f1204_rst;
  logic [31:0] f1204_rdata;
  sr_buffer_32_1 f1204(.wen(f1204_wen), .wdata(f1204_wdata), .clk(f1204_clk), .rst(f1204_rst), .rdata(f1204_rdata));
  assign f1204_clk = clk;
  assign f1204_rst = rst;
  // Bindings to f1204

  // f1206
  logic [0:0] f1206_wen;
  logic [31:0] f1206_wdata;
  logic [0:0] f1206_clk;
  logic [0:0] f1206_rst;
  logic [31:0] f1206_rdata;
  sr_buffer_32_1 f1206(.wen(f1206_wen), .wdata(f1206_wdata), .clk(f1206_clk), .rst(f1206_rst), .rdata(f1206_rdata));
  assign f1206_clk = clk;
  assign f1206_rst = rst;
  // Bindings to f1206

  // f1208
  logic [0:0] f1208_wen;
  logic [31:0] f1208_wdata;
  logic [0:0] f1208_clk;
  logic [0:0] f1208_rst;
  logic [31:0] f1208_rdata;
  sr_buffer_32_1 f1208(.wen(f1208_wen), .wdata(f1208_wdata), .clk(f1208_clk), .rst(f1208_rst), .rdata(f1208_rdata));
  assign f1208_clk = clk;
  assign f1208_rst = rst;
  // Bindings to f1208

  // f1210
  logic [0:0] f1210_wen;
  logic [31:0] f1210_wdata;
  logic [0:0] f1210_clk;
  logic [0:0] f1210_rst;
  logic [31:0] f1210_rdata;
  sr_buffer_32_1 f1210(.wen(f1210_wen), .wdata(f1210_wdata), .clk(f1210_clk), .rst(f1210_rst), .rdata(f1210_rdata));
  assign f1210_clk = clk;
  assign f1210_rst = rst;
  // Bindings to f1210

  // f1212
  logic [0:0] f1212_wen;
  logic [31:0] f1212_wdata;
  logic [0:0] f1212_clk;
  logic [0:0] f1212_rst;
  logic [31:0] f1212_rdata;
  sr_buffer_32_1 f1212(.wen(f1212_wen), .wdata(f1212_wdata), .clk(f1212_clk), .rst(f1212_rst), .rdata(f1212_rdata));
  assign f1212_clk = clk;
  assign f1212_rst = rst;
  // Bindings to f1212

  // f1214
  logic [0:0] f1214_wen;
  logic [31:0] f1214_wdata;
  logic [0:0] f1214_clk;
  logic [0:0] f1214_rst;
  logic [31:0] f1214_rdata;
  sr_buffer_32_1 f1214(.wen(f1214_wen), .wdata(f1214_wdata), .clk(f1214_clk), .rst(f1214_rst), .rdata(f1214_rdata));
  assign f1214_clk = clk;
  assign f1214_rst = rst;
  // Bindings to f1214

  // f1216
  logic [0:0] f1216_wen;
  logic [31:0] f1216_wdata;
  logic [0:0] f1216_clk;
  logic [0:0] f1216_rst;
  logic [31:0] f1216_rdata;
  sr_buffer_32_1 f1216(.wen(f1216_wen), .wdata(f1216_wdata), .clk(f1216_clk), .rst(f1216_rst), .rdata(f1216_rdata));
  assign f1216_clk = clk;
  assign f1216_rst = rst;
  // Bindings to f1216

  // f1218
  logic [0:0] f1218_wen;
  logic [31:0] f1218_wdata;
  logic [0:0] f1218_clk;
  logic [0:0] f1218_rst;
  logic [31:0] f1218_rdata;
  sr_buffer_32_1 f1218(.wen(f1218_wen), .wdata(f1218_wdata), .clk(f1218_clk), .rst(f1218_rst), .rdata(f1218_rdata));
  assign f1218_clk = clk;
  assign f1218_rst = rst;
  // Bindings to f1218

  // f1220
  logic [0:0] f1220_wen;
  logic [31:0] f1220_wdata;
  logic [0:0] f1220_clk;
  logic [0:0] f1220_rst;
  logic [31:0] f1220_rdata;
  sr_buffer_32_1 f1220(.wen(f1220_wen), .wdata(f1220_wdata), .clk(f1220_clk), .rst(f1220_rst), .rdata(f1220_rdata));
  assign f1220_clk = clk;
  assign f1220_rst = rst;
  // Bindings to f1220

  // f1222
  logic [0:0] f1222_wen;
  logic [31:0] f1222_wdata;
  logic [0:0] f1222_clk;
  logic [0:0] f1222_rst;
  logic [31:0] f1222_rdata;
  sr_buffer_32_1 f1222(.wen(f1222_wen), .wdata(f1222_wdata), .clk(f1222_clk), .rst(f1222_rst), .rdata(f1222_rdata));
  assign f1222_clk = clk;
  assign f1222_rst = rst;
  // Bindings to f1222

  // f1224
  logic [0:0] f1224_wen;
  logic [31:0] f1224_wdata;
  logic [0:0] f1224_clk;
  logic [0:0] f1224_rst;
  logic [31:0] f1224_rdata;
  sr_buffer_32_1 f1224(.wen(f1224_wen), .wdata(f1224_wdata), .clk(f1224_clk), .rst(f1224_rst), .rdata(f1224_rdata));
  assign f1224_clk = clk;
  assign f1224_rst = rst;
  // Bindings to f1224

  // f1226
  logic [0:0] f1226_wen;
  logic [31:0] f1226_wdata;
  logic [0:0] f1226_clk;
  logic [0:0] f1226_rst;
  logic [31:0] f1226_rdata;
  sr_buffer_32_1 f1226(.wen(f1226_wen), .wdata(f1226_wdata), .clk(f1226_clk), .rst(f1226_rst), .rdata(f1226_rdata));
  assign f1226_clk = clk;
  assign f1226_rst = rst;
  // Bindings to f1226

  // f1228
  logic [0:0] f1228_wen;
  logic [31:0] f1228_wdata;
  logic [0:0] f1228_clk;
  logic [0:0] f1228_rst;
  logic [31:0] f1228_rdata;
  sr_buffer_32_1 f1228(.wen(f1228_wen), .wdata(f1228_wdata), .clk(f1228_clk), .rst(f1228_rst), .rdata(f1228_rdata));
  assign f1228_clk = clk;
  assign f1228_rst = rst;
  // Bindings to f1228

  // f1230
  logic [0:0] f1230_wen;
  logic [31:0] f1230_wdata;
  logic [0:0] f1230_clk;
  logic [0:0] f1230_rst;
  logic [31:0] f1230_rdata;
  sr_buffer_32_1 f1230(.wen(f1230_wen), .wdata(f1230_wdata), .clk(f1230_clk), .rst(f1230_rst), .rdata(f1230_rdata));
  assign f1230_clk = clk;
  assign f1230_rst = rst;
  // Bindings to f1230

  // f1232
  logic [0:0] f1232_wen;
  logic [31:0] f1232_wdata;
  logic [0:0] f1232_clk;
  logic [0:0] f1232_rst;
  logic [31:0] f1232_rdata;
  sr_buffer_32_1 f1232(.wen(f1232_wen), .wdata(f1232_wdata), .clk(f1232_clk), .rst(f1232_rst), .rdata(f1232_rdata));
  assign f1232_clk = clk;
  assign f1232_rst = rst;
  // Bindings to f1232

  // f1234
  logic [0:0] f1234_wen;
  logic [31:0] f1234_wdata;
  logic [0:0] f1234_clk;
  logic [0:0] f1234_rst;
  logic [31:0] f1234_rdata;
  sr_buffer_32_1 f1234(.wen(f1234_wen), .wdata(f1234_wdata), .clk(f1234_clk), .rst(f1234_rst), .rdata(f1234_rdata));
  assign f1234_clk = clk;
  assign f1234_rst = rst;
  // Bindings to f1234

  // f1236
  logic [0:0] f1236_wen;
  logic [31:0] f1236_wdata;
  logic [0:0] f1236_clk;
  logic [0:0] f1236_rst;
  logic [31:0] f1236_rdata;
  sr_buffer_32_1 f1236(.wen(f1236_wen), .wdata(f1236_wdata), .clk(f1236_clk), .rst(f1236_rst), .rdata(f1236_rdata));
  assign f1236_clk = clk;
  assign f1236_rst = rst;
  // Bindings to f1236

  // f1238
  logic [0:0] f1238_wen;
  logic [31:0] f1238_wdata;
  logic [0:0] f1238_clk;
  logic [0:0] f1238_rst;
  logic [31:0] f1238_rdata;
  sr_buffer_32_1 f1238(.wen(f1238_wen), .wdata(f1238_wdata), .clk(f1238_clk), .rst(f1238_rst), .rdata(f1238_rdata));
  assign f1238_clk = clk;
  assign f1238_rst = rst;
  // Bindings to f1238

  // f1240
  logic [0:0] f1240_wen;
  logic [31:0] f1240_wdata;
  logic [0:0] f1240_clk;
  logic [0:0] f1240_rst;
  logic [31:0] f1240_rdata;
  sr_buffer_32_1 f1240(.wen(f1240_wen), .wdata(f1240_wdata), .clk(f1240_clk), .rst(f1240_rst), .rdata(f1240_rdata));
  assign f1240_clk = clk;
  assign f1240_rst = rst;
  // Bindings to f1240

  // f1242
  logic [0:0] f1242_wen;
  logic [31:0] f1242_wdata;
  logic [0:0] f1242_clk;
  logic [0:0] f1242_rst;
  logic [31:0] f1242_rdata;
  sr_buffer_32_1 f1242(.wen(f1242_wen), .wdata(f1242_wdata), .clk(f1242_clk), .rst(f1242_rst), .rdata(f1242_rdata));
  assign f1242_clk = clk;
  assign f1242_rst = rst;
  // Bindings to f1242

  // f1244
  logic [0:0] f1244_wen;
  logic [31:0] f1244_wdata;
  logic [0:0] f1244_clk;
  logic [0:0] f1244_rst;
  logic [31:0] f1244_rdata;
  sr_buffer_32_1 f1244(.wen(f1244_wen), .wdata(f1244_wdata), .clk(f1244_clk), .rst(f1244_rst), .rdata(f1244_rdata));
  assign f1244_clk = clk;
  assign f1244_rst = rst;
  // Bindings to f1244

  // f1246
  logic [0:0] f1246_wen;
  logic [31:0] f1246_wdata;
  logic [0:0] f1246_clk;
  logic [0:0] f1246_rst;
  logic [31:0] f1246_rdata;
  sr_buffer_32_1 f1246(.wen(f1246_wen), .wdata(f1246_wdata), .clk(f1246_clk), .rst(f1246_rst), .rdata(f1246_rdata));
  assign f1246_clk = clk;
  assign f1246_rst = rst;
  // Bindings to f1246

  // f1248
  logic [0:0] f1248_wen;
  logic [31:0] f1248_wdata;
  logic [0:0] f1248_clk;
  logic [0:0] f1248_rst;
  logic [31:0] f1248_rdata;
  sr_buffer_32_1 f1248(.wen(f1248_wen), .wdata(f1248_wdata), .clk(f1248_clk), .rst(f1248_rst), .rdata(f1248_rdata));
  assign f1248_clk = clk;
  assign f1248_rst = rst;
  // Bindings to f1248



endmodule


module in_wire_final_merged_1_update_0_write_wdata(output [31:0] final_merged_1_update_0_write_wdata);

endmodule


module in_wire_final_merged_0_update_0_read_dummy(output [31:0] final_merged_0_update_0_read_dummy);

endmodule


module out_wire_final_merged_0_update_0_read_rdata(input [31:0] final_merged_0_update_0_read_rdata);

endmodule


module final_merged_2_final_merged_2_update_0_write0_to_final_merged_1_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f314
  logic [0:0] f314_wen;
  logic [31:0] f314_wdata;
  logic [0:0] f314_clk;
  logic [0:0] f314_rst;
  logic [31:0] f314_rdata;
  sr_buffer_32_1 f314(.wen(f314_wen), .wdata(f314_wdata), .clk(f314_clk), .rst(f314_rst), .rdata(f314_rdata));
  assign f314_clk = clk;
  assign f314_rst = rst;
  // Bindings to f314

  // f316
  logic [0:0] f316_wen;
  logic [31:0] f316_wdata;
  logic [0:0] f316_clk;
  logic [0:0] f316_rst;
  logic [31:0] f316_rdata;
  sr_buffer_32_1 f316(.wen(f316_wen), .wdata(f316_wdata), .clk(f316_clk), .rst(f316_rst), .rdata(f316_rdata));
  assign f316_clk = clk;
  assign f316_rst = rst;
  // Bindings to f316

  // f318
  logic [0:0] f318_wen;
  logic [31:0] f318_wdata;
  logic [0:0] f318_clk;
  logic [0:0] f318_rst;
  logic [31:0] f318_rdata;
  sr_buffer_32_1 f318(.wen(f318_wen), .wdata(f318_wdata), .clk(f318_clk), .rst(f318_rst), .rdata(f318_rdata));
  assign f318_clk = clk;
  assign f318_rst = rst;
  // Bindings to f318

  // f320
  logic [0:0] f320_wen;
  logic [31:0] f320_wdata;
  logic [0:0] f320_clk;
  logic [0:0] f320_rst;
  logic [31:0] f320_rdata;
  sr_buffer_32_1 f320(.wen(f320_wen), .wdata(f320_wdata), .clk(f320_clk), .rst(f320_rst), .rdata(f320_rdata));
  assign f320_clk = clk;
  assign f320_rst = rst;
  // Bindings to f320

  // f322
  logic [0:0] f322_wen;
  logic [31:0] f322_wdata;
  logic [0:0] f322_clk;
  logic [0:0] f322_rst;
  logic [31:0] f322_rdata;
  sr_buffer_32_1 f322(.wen(f322_wen), .wdata(f322_wdata), .clk(f322_clk), .rst(f322_rst), .rdata(f322_rdata));
  assign f322_clk = clk;
  assign f322_rst = rst;
  // Bindings to f322

  // f324
  logic [0:0] f324_wen;
  logic [31:0] f324_wdata;
  logic [0:0] f324_clk;
  logic [0:0] f324_rst;
  logic [31:0] f324_rdata;
  sr_buffer_32_1 f324(.wen(f324_wen), .wdata(f324_wdata), .clk(f324_clk), .rst(f324_rst), .rdata(f324_rdata));
  assign f324_clk = clk;
  assign f324_rst = rst;
  // Bindings to f324

  // f326
  logic [0:0] f326_wen;
  logic [31:0] f326_wdata;
  logic [0:0] f326_clk;
  logic [0:0] f326_rst;
  logic [31:0] f326_rdata;
  sr_buffer_32_1 f326(.wen(f326_wen), .wdata(f326_wdata), .clk(f326_clk), .rst(f326_rst), .rdata(f326_rdata));
  assign f326_clk = clk;
  assign f326_rst = rst;
  // Bindings to f326

  // f328
  logic [0:0] f328_wen;
  logic [31:0] f328_wdata;
  logic [0:0] f328_clk;
  logic [0:0] f328_rst;
  logic [31:0] f328_rdata;
  sr_buffer_32_1 f328(.wen(f328_wen), .wdata(f328_wdata), .clk(f328_clk), .rst(f328_rst), .rdata(f328_rdata));
  assign f328_clk = clk;
  assign f328_rst = rst;
  // Bindings to f328

  // f330
  logic [0:0] f330_wen;
  logic [31:0] f330_wdata;
  logic [0:0] f330_clk;
  logic [0:0] f330_rst;
  logic [31:0] f330_rdata;
  sr_buffer_32_1 f330(.wen(f330_wen), .wdata(f330_wdata), .clk(f330_clk), .rst(f330_rst), .rdata(f330_rdata));
  assign f330_clk = clk;
  assign f330_rst = rst;
  // Bindings to f330

  // f332
  logic [0:0] f332_wen;
  logic [31:0] f332_wdata;
  logic [0:0] f332_clk;
  logic [0:0] f332_rst;
  logic [31:0] f332_rdata;
  sr_buffer_32_1 f332(.wen(f332_wen), .wdata(f332_wdata), .clk(f332_clk), .rst(f332_rst), .rdata(f332_rdata));
  assign f332_clk = clk;
  assign f332_rst = rst;
  // Bindings to f332

  // f334
  logic [0:0] f334_wen;
  logic [31:0] f334_wdata;
  logic [0:0] f334_clk;
  logic [0:0] f334_rst;
  logic [31:0] f334_rdata;
  sr_buffer_32_1 f334(.wen(f334_wen), .wdata(f334_wdata), .clk(f334_clk), .rst(f334_rst), .rdata(f334_rdata));
  assign f334_clk = clk;
  assign f334_rst = rst;
  // Bindings to f334

  // f336
  logic [0:0] f336_wen;
  logic [31:0] f336_wdata;
  logic [0:0] f336_clk;
  logic [0:0] f336_rst;
  logic [31:0] f336_rdata;
  sr_buffer_32_1 f336(.wen(f336_wen), .wdata(f336_wdata), .clk(f336_clk), .rst(f336_rst), .rdata(f336_rdata));
  assign f336_clk = clk;
  assign f336_rst = rst;
  // Bindings to f336

  // f338
  logic [0:0] f338_wen;
  logic [31:0] f338_wdata;
  logic [0:0] f338_clk;
  logic [0:0] f338_rst;
  logic [31:0] f338_rdata;
  sr_buffer_32_1 f338(.wen(f338_wen), .wdata(f338_wdata), .clk(f338_clk), .rst(f338_rst), .rdata(f338_rdata));
  assign f338_clk = clk;
  assign f338_rst = rst;
  // Bindings to f338

  // f340
  logic [0:0] f340_wen;
  logic [31:0] f340_wdata;
  logic [0:0] f340_clk;
  logic [0:0] f340_rst;
  logic [31:0] f340_rdata;
  sr_buffer_32_1 f340(.wen(f340_wen), .wdata(f340_wdata), .clk(f340_clk), .rst(f340_rst), .rdata(f340_rdata));
  assign f340_clk = clk;
  assign f340_rst = rst;
  // Bindings to f340

  // f342
  logic [0:0] f342_wen;
  logic [31:0] f342_wdata;
  logic [0:0] f342_clk;
  logic [0:0] f342_rst;
  logic [31:0] f342_rdata;
  sr_buffer_32_1 f342(.wen(f342_wen), .wdata(f342_wdata), .clk(f342_clk), .rst(f342_rst), .rdata(f342_rdata));
  assign f342_clk = clk;
  assign f342_rst = rst;
  // Bindings to f342

  // f344
  logic [0:0] f344_wen;
  logic [31:0] f344_wdata;
  logic [0:0] f344_clk;
  logic [0:0] f344_rst;
  logic [31:0] f344_rdata;
  sr_buffer_32_1 f344(.wen(f344_wen), .wdata(f344_wdata), .clk(f344_clk), .rst(f344_rst), .rdata(f344_rdata));
  assign f344_clk = clk;
  assign f344_rst = rst;
  // Bindings to f344

  // f346
  logic [0:0] f346_wen;
  logic [31:0] f346_wdata;
  logic [0:0] f346_clk;
  logic [0:0] f346_rst;
  logic [31:0] f346_rdata;
  sr_buffer_32_1 f346(.wen(f346_wen), .wdata(f346_wdata), .clk(f346_clk), .rst(f346_rst), .rdata(f346_rdata));
  assign f346_clk = clk;
  assign f346_rst = rst;
  // Bindings to f346

  // f348
  logic [0:0] f348_wen;
  logic [31:0] f348_wdata;
  logic [0:0] f348_clk;
  logic [0:0] f348_rst;
  logic [31:0] f348_rdata;
  sr_buffer_32_1 f348(.wen(f348_wen), .wdata(f348_wdata), .clk(f348_clk), .rst(f348_rst), .rdata(f348_rdata));
  assign f348_clk = clk;
  assign f348_rst = rst;
  // Bindings to f348

  // f350
  logic [0:0] f350_wen;
  logic [31:0] f350_wdata;
  logic [0:0] f350_clk;
  logic [0:0] f350_rst;
  logic [31:0] f350_rdata;
  sr_buffer_32_1 f350(.wen(f350_wen), .wdata(f350_wdata), .clk(f350_clk), .rst(f350_rst), .rdata(f350_rdata));
  assign f350_clk = clk;
  assign f350_rst = rst;
  // Bindings to f350

  // f352
  logic [0:0] f352_wen;
  logic [31:0] f352_wdata;
  logic [0:0] f352_clk;
  logic [0:0] f352_rst;
  logic [31:0] f352_rdata;
  sr_buffer_32_1 f352(.wen(f352_wen), .wdata(f352_wdata), .clk(f352_clk), .rst(f352_rst), .rdata(f352_rdata));
  assign f352_clk = clk;
  assign f352_rst = rst;
  // Bindings to f352

  // f354
  logic [0:0] f354_wen;
  logic [31:0] f354_wdata;
  logic [0:0] f354_clk;
  logic [0:0] f354_rst;
  logic [31:0] f354_rdata;
  sr_buffer_32_1 f354(.wen(f354_wen), .wdata(f354_wdata), .clk(f354_clk), .rst(f354_rst), .rdata(f354_rdata));
  assign f354_clk = clk;
  assign f354_rst = rst;
  // Bindings to f354

  // f356
  logic [0:0] f356_wen;
  logic [31:0] f356_wdata;
  logic [0:0] f356_clk;
  logic [0:0] f356_rst;
  logic [31:0] f356_rdata;
  sr_buffer_32_1 f356(.wen(f356_wen), .wdata(f356_wdata), .clk(f356_clk), .rst(f356_rst), .rdata(f356_rdata));
  assign f356_clk = clk;
  assign f356_rst = rst;
  // Bindings to f356

  // f358
  logic [0:0] f358_wen;
  logic [31:0] f358_wdata;
  logic [0:0] f358_clk;
  logic [0:0] f358_rst;
  logic [31:0] f358_rdata;
  sr_buffer_32_1 f358(.wen(f358_wen), .wdata(f358_wdata), .clk(f358_clk), .rst(f358_rst), .rdata(f358_rdata));
  assign f358_clk = clk;
  assign f358_rst = rst;
  // Bindings to f358

  // f360
  logic [0:0] f360_wen;
  logic [31:0] f360_wdata;
  logic [0:0] f360_clk;
  logic [0:0] f360_rst;
  logic [31:0] f360_rdata;
  sr_buffer_32_1 f360(.wen(f360_wen), .wdata(f360_wdata), .clk(f360_clk), .rst(f360_rst), .rdata(f360_rdata));
  assign f360_clk = clk;
  assign f360_rst = rst;
  // Bindings to f360

  // f362
  logic [0:0] f362_wen;
  logic [31:0] f362_wdata;
  logic [0:0] f362_clk;
  logic [0:0] f362_rst;
  logic [31:0] f362_rdata;
  sr_buffer_32_1 f362(.wen(f362_wen), .wdata(f362_wdata), .clk(f362_clk), .rst(f362_rst), .rdata(f362_rdata));
  assign f362_clk = clk;
  assign f362_rst = rst;
  // Bindings to f362

  // f364
  logic [0:0] f364_wen;
  logic [31:0] f364_wdata;
  logic [0:0] f364_clk;
  logic [0:0] f364_rst;
  logic [31:0] f364_rdata;
  sr_buffer_32_1 f364(.wen(f364_wen), .wdata(f364_wdata), .clk(f364_clk), .rst(f364_rst), .rdata(f364_rdata));
  assign f364_clk = clk;
  assign f364_rst = rst;
  // Bindings to f364

  // f366
  logic [0:0] f366_wen;
  logic [31:0] f366_wdata;
  logic [0:0] f366_clk;
  logic [0:0] f366_rst;
  logic [31:0] f366_rdata;
  sr_buffer_32_1 f366(.wen(f366_wen), .wdata(f366_wdata), .clk(f366_clk), .rst(f366_rst), .rdata(f366_rdata));
  assign f366_clk = clk;
  assign f366_rst = rst;
  // Bindings to f366

  // f368
  logic [0:0] f368_wen;
  logic [31:0] f368_wdata;
  logic [0:0] f368_clk;
  logic [0:0] f368_rst;
  logic [31:0] f368_rdata;
  sr_buffer_32_1 f368(.wen(f368_wen), .wdata(f368_wdata), .clk(f368_clk), .rst(f368_rst), .rdata(f368_rdata));
  assign f368_clk = clk;
  assign f368_rst = rst;
  // Bindings to f368

  // f370
  logic [0:0] f370_wen;
  logic [31:0] f370_wdata;
  logic [0:0] f370_clk;
  logic [0:0] f370_rst;
  logic [31:0] f370_rdata;
  sr_buffer_32_1 f370(.wen(f370_wen), .wdata(f370_wdata), .clk(f370_clk), .rst(f370_rst), .rdata(f370_rdata));
  assign f370_clk = clk;
  assign f370_rst = rst;
  // Bindings to f370

  // f372
  logic [0:0] f372_wen;
  logic [31:0] f372_wdata;
  logic [0:0] f372_clk;
  logic [0:0] f372_rst;
  logic [31:0] f372_rdata;
  sr_buffer_32_1 f372(.wen(f372_wen), .wdata(f372_wdata), .clk(f372_clk), .rst(f372_rst), .rdata(f372_rdata));
  assign f372_clk = clk;
  assign f372_rst = rst;
  // Bindings to f372

  // f374
  logic [0:0] f374_wen;
  logic [31:0] f374_wdata;
  logic [0:0] f374_clk;
  logic [0:0] f374_rst;
  logic [31:0] f374_rdata;
  sr_buffer_32_1 f374(.wen(f374_wen), .wdata(f374_wdata), .clk(f374_clk), .rst(f374_rst), .rdata(f374_rdata));
  assign f374_clk = clk;
  assign f374_rst = rst;
  // Bindings to f374

  // f376
  logic [0:0] f376_wen;
  logic [31:0] f376_wdata;
  logic [0:0] f376_clk;
  logic [0:0] f376_rst;
  logic [31:0] f376_rdata;
  sr_buffer_32_1 f376(.wen(f376_wen), .wdata(f376_wdata), .clk(f376_clk), .rst(f376_rst), .rdata(f376_rdata));
  assign f376_clk = clk;
  assign f376_rst = rst;
  // Bindings to f376

  // f378
  logic [0:0] f378_wen;
  logic [31:0] f378_wdata;
  logic [0:0] f378_clk;
  logic [0:0] f378_rst;
  logic [31:0] f378_rdata;
  sr_buffer_32_1 f378(.wen(f378_wen), .wdata(f378_wdata), .clk(f378_clk), .rst(f378_rst), .rdata(f378_rdata));
  assign f378_clk = clk;
  assign f378_rst = rst;
  // Bindings to f378

  // f380
  logic [0:0] f380_wen;
  logic [31:0] f380_wdata;
  logic [0:0] f380_clk;
  logic [0:0] f380_rst;
  logic [31:0] f380_rdata;
  sr_buffer_32_1 f380(.wen(f380_wen), .wdata(f380_wdata), .clk(f380_clk), .rst(f380_rst), .rdata(f380_rdata));
  assign f380_clk = clk;
  assign f380_rst = rst;
  // Bindings to f380

  // f382
  logic [0:0] f382_wen;
  logic [31:0] f382_wdata;
  logic [0:0] f382_clk;
  logic [0:0] f382_rst;
  logic [31:0] f382_rdata;
  sr_buffer_32_1 f382(.wen(f382_wen), .wdata(f382_wdata), .clk(f382_clk), .rst(f382_rst), .rdata(f382_rdata));
  assign f382_clk = clk;
  assign f382_rst = rst;
  // Bindings to f382

  // f384
  logic [0:0] f384_wen;
  logic [31:0] f384_wdata;
  logic [0:0] f384_clk;
  logic [0:0] f384_rst;
  logic [31:0] f384_rdata;
  sr_buffer_32_1 f384(.wen(f384_wen), .wdata(f384_wdata), .clk(f384_clk), .rst(f384_rst), .rdata(f384_rdata));
  assign f384_clk = clk;
  assign f384_rst = rst;
  // Bindings to f384

  // f386
  logic [0:0] f386_wen;
  logic [31:0] f386_wdata;
  logic [0:0] f386_clk;
  logic [0:0] f386_rst;
  logic [31:0] f386_rdata;
  sr_buffer_32_1 f386(.wen(f386_wen), .wdata(f386_wdata), .clk(f386_clk), .rst(f386_rst), .rdata(f386_rdata));
  assign f386_clk = clk;
  assign f386_rst = rst;
  // Bindings to f386

  // f388
  logic [0:0] f388_wen;
  logic [31:0] f388_wdata;
  logic [0:0] f388_clk;
  logic [0:0] f388_rst;
  logic [31:0] f388_rdata;
  sr_buffer_32_1 f388(.wen(f388_wen), .wdata(f388_wdata), .clk(f388_clk), .rst(f388_rst), .rdata(f388_rdata));
  assign f388_clk = clk;
  assign f388_rst = rst;
  // Bindings to f388

  // f390
  logic [0:0] f390_wen;
  logic [31:0] f390_wdata;
  logic [0:0] f390_clk;
  logic [0:0] f390_rst;
  logic [31:0] f390_rdata;
  sr_buffer_32_1 f390(.wen(f390_wen), .wdata(f390_wdata), .clk(f390_clk), .rst(f390_rst), .rdata(f390_rdata));
  assign f390_clk = clk;
  assign f390_rst = rst;
  // Bindings to f390

  // f392
  logic [0:0] f392_wen;
  logic [31:0] f392_wdata;
  logic [0:0] f392_clk;
  logic [0:0] f392_rst;
  logic [31:0] f392_rdata;
  sr_buffer_32_1 f392(.wen(f392_wen), .wdata(f392_wdata), .clk(f392_clk), .rst(f392_rst), .rdata(f392_rdata));
  assign f392_clk = clk;
  assign f392_rst = rst;
  // Bindings to f392

  // f394
  logic [0:0] f394_wen;
  logic [31:0] f394_wdata;
  logic [0:0] f394_clk;
  logic [0:0] f394_rst;
  logic [31:0] f394_rdata;
  sr_buffer_32_1 f394(.wen(f394_wen), .wdata(f394_wdata), .clk(f394_clk), .rst(f394_rst), .rdata(f394_rdata));
  assign f394_clk = clk;
  assign f394_rst = rst;
  // Bindings to f394

  // f396
  logic [0:0] f396_wen;
  logic [31:0] f396_wdata;
  logic [0:0] f396_clk;
  logic [0:0] f396_rst;
  logic [31:0] f396_rdata;
  sr_buffer_32_1 f396(.wen(f396_wen), .wdata(f396_wdata), .clk(f396_clk), .rst(f396_rst), .rdata(f396_rdata));
  assign f396_clk = clk;
  assign f396_rst = rst;
  // Bindings to f396

  // f398
  logic [0:0] f398_wen;
  logic [31:0] f398_wdata;
  logic [0:0] f398_clk;
  logic [0:0] f398_rst;
  logic [31:0] f398_rdata;
  sr_buffer_32_1 f398(.wen(f398_wen), .wdata(f398_wdata), .clk(f398_clk), .rst(f398_rst), .rdata(f398_rdata));
  assign f398_clk = clk;
  assign f398_rst = rst;
  // Bindings to f398

  // f400
  logic [0:0] f400_wen;
  logic [31:0] f400_wdata;
  logic [0:0] f400_clk;
  logic [0:0] f400_rst;
  logic [31:0] f400_rdata;
  sr_buffer_32_1 f400(.wen(f400_wen), .wdata(f400_wdata), .clk(f400_clk), .rst(f400_rst), .rdata(f400_rdata));
  assign f400_clk = clk;
  assign f400_rst = rst;
  // Bindings to f400

  // f402
  logic [0:0] f402_wen;
  logic [31:0] f402_wdata;
  logic [0:0] f402_clk;
  logic [0:0] f402_rst;
  logic [31:0] f402_rdata;
  sr_buffer_32_1 f402(.wen(f402_wen), .wdata(f402_wdata), .clk(f402_clk), .rst(f402_rst), .rdata(f402_rdata));
  assign f402_clk = clk;
  assign f402_rst = rst;
  // Bindings to f402

  // f404
  logic [0:0] f404_wen;
  logic [31:0] f404_wdata;
  logic [0:0] f404_clk;
  logic [0:0] f404_rst;
  logic [31:0] f404_rdata;
  sr_buffer_32_1 f404(.wen(f404_wen), .wdata(f404_wdata), .clk(f404_clk), .rst(f404_rst), .rdata(f404_rdata));
  assign f404_clk = clk;
  assign f404_rst = rst;
  // Bindings to f404

  // f406
  logic [0:0] f406_wen;
  logic [31:0] f406_wdata;
  logic [0:0] f406_clk;
  logic [0:0] f406_rst;
  logic [31:0] f406_rdata;
  sr_buffer_32_1 f406(.wen(f406_wen), .wdata(f406_wdata), .clk(f406_clk), .rst(f406_rst), .rdata(f406_rdata));
  assign f406_clk = clk;
  assign f406_rst = rst;
  // Bindings to f406

  // f408
  logic [0:0] f408_wen;
  logic [31:0] f408_wdata;
  logic [0:0] f408_clk;
  logic [0:0] f408_rst;
  logic [31:0] f408_rdata;
  sr_buffer_32_1 f408(.wen(f408_wen), .wdata(f408_wdata), .clk(f408_clk), .rst(f408_rst), .rdata(f408_rdata));
  assign f408_clk = clk;
  assign f408_rst = rst;
  // Bindings to f408

  // f410
  logic [0:0] f410_wen;
  logic [31:0] f410_wdata;
  logic [0:0] f410_clk;
  logic [0:0] f410_rst;
  logic [31:0] f410_rdata;
  sr_buffer_32_1 f410(.wen(f410_wen), .wdata(f410_wdata), .clk(f410_clk), .rst(f410_rst), .rdata(f410_rdata));
  assign f410_clk = clk;
  assign f410_rst = rst;
  // Bindings to f410

  // f412
  logic [0:0] f412_wen;
  logic [31:0] f412_wdata;
  logic [0:0] f412_clk;
  logic [0:0] f412_rst;
  logic [31:0] f412_rdata;
  sr_buffer_32_1 f412(.wen(f412_wen), .wdata(f412_wdata), .clk(f412_clk), .rst(f412_rst), .rdata(f412_rdata));
  assign f412_clk = clk;
  assign f412_rst = rst;
  // Bindings to f412

  // f414
  logic [0:0] f414_wen;
  logic [31:0] f414_wdata;
  logic [0:0] f414_clk;
  logic [0:0] f414_rst;
  logic [31:0] f414_rdata;
  sr_buffer_32_1 f414(.wen(f414_wen), .wdata(f414_wdata), .clk(f414_clk), .rst(f414_rst), .rdata(f414_rdata));
  assign f414_clk = clk;
  assign f414_rst = rst;
  // Bindings to f414

  // f416
  logic [0:0] f416_wen;
  logic [31:0] f416_wdata;
  logic [0:0] f416_clk;
  logic [0:0] f416_rst;
  logic [31:0] f416_rdata;
  sr_buffer_32_1 f416(.wen(f416_wen), .wdata(f416_wdata), .clk(f416_clk), .rst(f416_rst), .rdata(f416_rdata));
  assign f416_clk = clk;
  assign f416_rst = rst;
  // Bindings to f416

  // f418
  logic [0:0] f418_wen;
  logic [31:0] f418_wdata;
  logic [0:0] f418_clk;
  logic [0:0] f418_rst;
  logic [31:0] f418_rdata;
  sr_buffer_32_1 f418(.wen(f418_wen), .wdata(f418_wdata), .clk(f418_clk), .rst(f418_rst), .rdata(f418_rdata));
  assign f418_clk = clk;
  assign f418_rst = rst;
  // Bindings to f418

  // f420
  logic [0:0] f420_wen;
  logic [31:0] f420_wdata;
  logic [0:0] f420_clk;
  logic [0:0] f420_rst;
  logic [31:0] f420_rdata;
  sr_buffer_32_1 f420(.wen(f420_wen), .wdata(f420_wdata), .clk(f420_clk), .rst(f420_rst), .rdata(f420_rdata));
  assign f420_clk = clk;
  assign f420_rst = rst;
  // Bindings to f420

  // f422
  logic [0:0] f422_wen;
  logic [31:0] f422_wdata;
  logic [0:0] f422_clk;
  logic [0:0] f422_rst;
  logic [31:0] f422_rdata;
  sr_buffer_32_1 f422(.wen(f422_wen), .wdata(f422_wdata), .clk(f422_clk), .rst(f422_rst), .rdata(f422_rdata));
  assign f422_clk = clk;
  assign f422_rst = rst;
  // Bindings to f422

  // f424
  logic [0:0] f424_wen;
  logic [31:0] f424_wdata;
  logic [0:0] f424_clk;
  logic [0:0] f424_rst;
  logic [31:0] f424_rdata;
  sr_buffer_32_1 f424(.wen(f424_wen), .wdata(f424_wdata), .clk(f424_clk), .rst(f424_rst), .rdata(f424_rdata));
  assign f424_clk = clk;
  assign f424_rst = rst;
  // Bindings to f424

  // f426
  logic [0:0] f426_wen;
  logic [31:0] f426_wdata;
  logic [0:0] f426_clk;
  logic [0:0] f426_rst;
  logic [31:0] f426_rdata;
  sr_buffer_32_1 f426(.wen(f426_wen), .wdata(f426_wdata), .clk(f426_clk), .rst(f426_rst), .rdata(f426_rdata));
  assign f426_clk = clk;
  assign f426_rst = rst;
  // Bindings to f426

  // f428
  logic [0:0] f428_wen;
  logic [31:0] f428_wdata;
  logic [0:0] f428_clk;
  logic [0:0] f428_rst;
  logic [31:0] f428_rdata;
  sr_buffer_32_1 f428(.wen(f428_wen), .wdata(f428_wdata), .clk(f428_clk), .rst(f428_rst), .rdata(f428_rdata));
  assign f428_clk = clk;
  assign f428_rst = rst;
  // Bindings to f428

  // f430
  logic [0:0] f430_wen;
  logic [31:0] f430_wdata;
  logic [0:0] f430_clk;
  logic [0:0] f430_rst;
  logic [31:0] f430_rdata;
  sr_buffer_32_1 f430(.wen(f430_wen), .wdata(f430_wdata), .clk(f430_clk), .rst(f430_rst), .rdata(f430_rdata));
  assign f430_clk = clk;
  assign f430_rst = rst;
  // Bindings to f430

  // f432
  logic [0:0] f432_wen;
  logic [31:0] f432_wdata;
  logic [0:0] f432_clk;
  logic [0:0] f432_rst;
  logic [31:0] f432_rdata;
  sr_buffer_32_1 f432(.wen(f432_wen), .wdata(f432_wdata), .clk(f432_clk), .rst(f432_rst), .rdata(f432_rdata));
  assign f432_clk = clk;
  assign f432_rst = rst;
  // Bindings to f432

  // f434
  logic [0:0] f434_wen;
  logic [31:0] f434_wdata;
  logic [0:0] f434_clk;
  logic [0:0] f434_rst;
  logic [31:0] f434_rdata;
  sr_buffer_32_1 f434(.wen(f434_wen), .wdata(f434_wdata), .clk(f434_clk), .rst(f434_rst), .rdata(f434_rdata));
  assign f434_clk = clk;
  assign f434_rst = rst;
  // Bindings to f434

  // f436
  logic [0:0] f436_wen;
  logic [31:0] f436_wdata;
  logic [0:0] f436_clk;
  logic [0:0] f436_rst;
  logic [31:0] f436_rdata;
  sr_buffer_32_1 f436(.wen(f436_wen), .wdata(f436_wdata), .clk(f436_clk), .rst(f436_rst), .rdata(f436_rdata));
  assign f436_clk = clk;
  assign f436_rst = rst;
  // Bindings to f436

  // f438
  logic [0:0] f438_wen;
  logic [31:0] f438_wdata;
  logic [0:0] f438_clk;
  logic [0:0] f438_rst;
  logic [31:0] f438_rdata;
  sr_buffer_32_1 f438(.wen(f438_wen), .wdata(f438_wdata), .clk(f438_clk), .rst(f438_rst), .rdata(f438_rdata));
  assign f438_clk = clk;
  assign f438_rst = rst;
  // Bindings to f438

  // f440
  logic [0:0] f440_wen;
  logic [31:0] f440_wdata;
  logic [0:0] f440_clk;
  logic [0:0] f440_rst;
  logic [31:0] f440_rdata;
  sr_buffer_32_1 f440(.wen(f440_wen), .wdata(f440_wdata), .clk(f440_clk), .rst(f440_rst), .rdata(f440_rdata));
  assign f440_clk = clk;
  assign f440_rst = rst;
  // Bindings to f440

  // f442
  logic [0:0] f442_wen;
  logic [31:0] f442_wdata;
  logic [0:0] f442_clk;
  logic [0:0] f442_rst;
  logic [31:0] f442_rdata;
  sr_buffer_32_1 f442(.wen(f442_wen), .wdata(f442_wdata), .clk(f442_clk), .rst(f442_rst), .rdata(f442_rdata));
  assign f442_clk = clk;
  assign f442_rst = rst;
  // Bindings to f442

  // f444
  logic [0:0] f444_wen;
  logic [31:0] f444_wdata;
  logic [0:0] f444_clk;
  logic [0:0] f444_rst;
  logic [31:0] f444_rdata;
  sr_buffer_32_1 f444(.wen(f444_wen), .wdata(f444_wdata), .clk(f444_clk), .rst(f444_rst), .rdata(f444_rdata));
  assign f444_clk = clk;
  assign f444_rst = rst;
  // Bindings to f444

  // f446
  logic [0:0] f446_wen;
  logic [31:0] f446_wdata;
  logic [0:0] f446_clk;
  logic [0:0] f446_rst;
  logic [31:0] f446_rdata;
  sr_buffer_32_1 f446(.wen(f446_wen), .wdata(f446_wdata), .clk(f446_clk), .rst(f446_rst), .rdata(f446_rdata));
  assign f446_clk = clk;
  assign f446_rst = rst;
  // Bindings to f446

  // f448
  logic [0:0] f448_wen;
  logic [31:0] f448_wdata;
  logic [0:0] f448_clk;
  logic [0:0] f448_rst;
  logic [31:0] f448_rdata;
  sr_buffer_32_1 f448(.wen(f448_wen), .wdata(f448_wdata), .clk(f448_clk), .rst(f448_rst), .rdata(f448_rdata));
  assign f448_clk = clk;
  assign f448_rst = rst;
  // Bindings to f448

  // f450
  logic [0:0] f450_wen;
  logic [31:0] f450_wdata;
  logic [0:0] f450_clk;
  logic [0:0] f450_rst;
  logic [31:0] f450_rdata;
  sr_buffer_32_1 f450(.wen(f450_wen), .wdata(f450_wdata), .clk(f450_clk), .rst(f450_rst), .rdata(f450_rdata));
  assign f450_clk = clk;
  assign f450_rst = rst;
  // Bindings to f450

  // f452
  logic [0:0] f452_wen;
  logic [31:0] f452_wdata;
  logic [0:0] f452_clk;
  logic [0:0] f452_rst;
  logic [31:0] f452_rdata;
  sr_buffer_32_1 f452(.wen(f452_wen), .wdata(f452_wdata), .clk(f452_clk), .rst(f452_rst), .rdata(f452_rdata));
  assign f452_clk = clk;
  assign f452_rst = rst;
  // Bindings to f452

  // f454
  logic [0:0] f454_wen;
  logic [31:0] f454_wdata;
  logic [0:0] f454_clk;
  logic [0:0] f454_rst;
  logic [31:0] f454_rdata;
  sr_buffer_32_1 f454(.wen(f454_wen), .wdata(f454_wdata), .clk(f454_clk), .rst(f454_rst), .rdata(f454_rdata));
  assign f454_clk = clk;
  assign f454_rst = rst;
  // Bindings to f454

  // f456
  logic [0:0] f456_wen;
  logic [31:0] f456_wdata;
  logic [0:0] f456_clk;
  logic [0:0] f456_rst;
  logic [31:0] f456_rdata;
  sr_buffer_32_1 f456(.wen(f456_wen), .wdata(f456_wdata), .clk(f456_clk), .rst(f456_rst), .rdata(f456_rdata));
  assign f456_clk = clk;
  assign f456_rst = rst;
  // Bindings to f456

  // f458
  logic [0:0] f458_wen;
  logic [31:0] f458_wdata;
  logic [0:0] f458_clk;
  logic [0:0] f458_rst;
  logic [31:0] f458_rdata;
  sr_buffer_32_1 f458(.wen(f458_wen), .wdata(f458_wdata), .clk(f458_clk), .rst(f458_rst), .rdata(f458_rdata));
  assign f458_clk = clk;
  assign f458_rst = rst;
  // Bindings to f458

  // f460
  logic [0:0] f460_wen;
  logic [31:0] f460_wdata;
  logic [0:0] f460_clk;
  logic [0:0] f460_rst;
  logic [31:0] f460_rdata;
  sr_buffer_32_1 f460(.wen(f460_wen), .wdata(f460_wdata), .clk(f460_clk), .rst(f460_rst), .rdata(f460_rdata));
  assign f460_clk = clk;
  assign f460_rst = rst;
  // Bindings to f460

  // f462
  logic [0:0] f462_wen;
  logic [31:0] f462_wdata;
  logic [0:0] f462_clk;
  logic [0:0] f462_rst;
  logic [31:0] f462_rdata;
  sr_buffer_32_1 f462(.wen(f462_wen), .wdata(f462_wdata), .clk(f462_clk), .rst(f462_rst), .rdata(f462_rdata));
  assign f462_clk = clk;
  assign f462_rst = rst;
  // Bindings to f462

  // f464
  logic [0:0] f464_wen;
  logic [31:0] f464_wdata;
  logic [0:0] f464_clk;
  logic [0:0] f464_rst;
  logic [31:0] f464_rdata;
  sr_buffer_32_1 f464(.wen(f464_wen), .wdata(f464_wdata), .clk(f464_clk), .rst(f464_rst), .rdata(f464_rdata));
  assign f464_clk = clk;
  assign f464_rst = rst;
  // Bindings to f464

  // f466
  logic [0:0] f466_wen;
  logic [31:0] f466_wdata;
  logic [0:0] f466_clk;
  logic [0:0] f466_rst;
  logic [31:0] f466_rdata;
  sr_buffer_32_1 f466(.wen(f466_wen), .wdata(f466_wdata), .clk(f466_clk), .rst(f466_rst), .rdata(f466_rdata));
  assign f466_clk = clk;
  assign f466_rst = rst;
  // Bindings to f466

  // f468
  logic [0:0] f468_wen;
  logic [31:0] f468_wdata;
  logic [0:0] f468_clk;
  logic [0:0] f468_rst;
  logic [31:0] f468_rdata;
  sr_buffer_32_1 f468(.wen(f468_wen), .wdata(f468_wdata), .clk(f468_clk), .rst(f468_rst), .rdata(f468_rdata));
  assign f468_clk = clk;
  assign f468_rst = rst;
  // Bindings to f468

  // f470
  logic [0:0] f470_wen;
  logic [31:0] f470_wdata;
  logic [0:0] f470_clk;
  logic [0:0] f470_rst;
  logic [31:0] f470_rdata;
  sr_buffer_32_1 f470(.wen(f470_wen), .wdata(f470_wdata), .clk(f470_clk), .rst(f470_rst), .rdata(f470_rdata));
  assign f470_clk = clk;
  assign f470_rst = rst;
  // Bindings to f470

  // f472
  logic [0:0] f472_wen;
  logic [31:0] f472_wdata;
  logic [0:0] f472_clk;
  logic [0:0] f472_rst;
  logic [31:0] f472_rdata;
  sr_buffer_32_1 f472(.wen(f472_wen), .wdata(f472_wdata), .clk(f472_clk), .rst(f472_rst), .rdata(f472_rdata));
  assign f472_clk = clk;
  assign f472_rst = rst;
  // Bindings to f472

  // f474
  logic [0:0] f474_wen;
  logic [31:0] f474_wdata;
  logic [0:0] f474_clk;
  logic [0:0] f474_rst;
  logic [31:0] f474_rdata;
  sr_buffer_32_1 f474(.wen(f474_wen), .wdata(f474_wdata), .clk(f474_clk), .rst(f474_rst), .rdata(f474_rdata));
  assign f474_clk = clk;
  assign f474_rst = rst;
  // Bindings to f474

  // f476
  logic [0:0] f476_wen;
  logic [31:0] f476_wdata;
  logic [0:0] f476_clk;
  logic [0:0] f476_rst;
  logic [31:0] f476_rdata;
  sr_buffer_32_1 f476(.wen(f476_wen), .wdata(f476_wdata), .clk(f476_clk), .rst(f476_rst), .rdata(f476_rdata));
  assign f476_clk = clk;
  assign f476_rst = rst;
  // Bindings to f476

  // f478
  logic [0:0] f478_wen;
  logic [31:0] f478_wdata;
  logic [0:0] f478_clk;
  logic [0:0] f478_rst;
  logic [31:0] f478_rdata;
  sr_buffer_32_1 f478(.wen(f478_wen), .wdata(f478_wdata), .clk(f478_clk), .rst(f478_rst), .rdata(f478_rdata));
  assign f478_clk = clk;
  assign f478_rst = rst;
  // Bindings to f478

  // f480
  logic [0:0] f480_wen;
  logic [31:0] f480_wdata;
  logic [0:0] f480_clk;
  logic [0:0] f480_rst;
  logic [31:0] f480_rdata;
  sr_buffer_32_1 f480(.wen(f480_wen), .wdata(f480_wdata), .clk(f480_clk), .rst(f480_rst), .rdata(f480_rdata));
  assign f480_clk = clk;
  assign f480_rst = rst;
  // Bindings to f480

  // f482
  logic [0:0] f482_wen;
  logic [31:0] f482_wdata;
  logic [0:0] f482_clk;
  logic [0:0] f482_rst;
  logic [31:0] f482_rdata;
  sr_buffer_32_1 f482(.wen(f482_wen), .wdata(f482_wdata), .clk(f482_clk), .rst(f482_rst), .rdata(f482_rdata));
  assign f482_clk = clk;
  assign f482_rst = rst;
  // Bindings to f482

  // f484
  logic [0:0] f484_wen;
  logic [31:0] f484_wdata;
  logic [0:0] f484_clk;
  logic [0:0] f484_rst;
  logic [31:0] f484_rdata;
  sr_buffer_32_1 f484(.wen(f484_wen), .wdata(f484_wdata), .clk(f484_clk), .rst(f484_rst), .rdata(f484_rdata));
  assign f484_clk = clk;
  assign f484_rst = rst;
  // Bindings to f484

  // f486
  logic [0:0] f486_wen;
  logic [31:0] f486_wdata;
  logic [0:0] f486_clk;
  logic [0:0] f486_rst;
  logic [31:0] f486_rdata;
  sr_buffer_32_1 f486(.wen(f486_wen), .wdata(f486_wdata), .clk(f486_clk), .rst(f486_rst), .rdata(f486_rdata));
  assign f486_clk = clk;
  assign f486_rst = rst;
  // Bindings to f486

  // f488
  logic [0:0] f488_wen;
  logic [31:0] f488_wdata;
  logic [0:0] f488_clk;
  logic [0:0] f488_rst;
  logic [31:0] f488_rdata;
  sr_buffer_32_1 f488(.wen(f488_wen), .wdata(f488_wdata), .clk(f488_clk), .rst(f488_rst), .rdata(f488_rdata));
  assign f488_clk = clk;
  assign f488_rst = rst;
  // Bindings to f488

  // f490
  logic [0:0] f490_wen;
  logic [31:0] f490_wdata;
  logic [0:0] f490_clk;
  logic [0:0] f490_rst;
  logic [31:0] f490_rdata;
  sr_buffer_32_1 f490(.wen(f490_wen), .wdata(f490_wdata), .clk(f490_clk), .rst(f490_rst), .rdata(f490_rdata));
  assign f490_clk = clk;
  assign f490_rst = rst;
  // Bindings to f490

  // f492
  logic [0:0] f492_wen;
  logic [31:0] f492_wdata;
  logic [0:0] f492_clk;
  logic [0:0] f492_rst;
  logic [31:0] f492_rdata;
  sr_buffer_32_1 f492(.wen(f492_wen), .wdata(f492_wdata), .clk(f492_clk), .rst(f492_rst), .rdata(f492_rdata));
  assign f492_clk = clk;
  assign f492_rst = rst;
  // Bindings to f492

  // f494
  logic [0:0] f494_wen;
  logic [31:0] f494_wdata;
  logic [0:0] f494_clk;
  logic [0:0] f494_rst;
  logic [31:0] f494_rdata;
  sr_buffer_32_1 f494(.wen(f494_wen), .wdata(f494_wdata), .clk(f494_clk), .rst(f494_rst), .rdata(f494_rdata));
  assign f494_clk = clk;
  assign f494_rst = rst;
  // Bindings to f494

  // f496
  logic [0:0] f496_wen;
  logic [31:0] f496_wdata;
  logic [0:0] f496_clk;
  logic [0:0] f496_rst;
  logic [31:0] f496_rdata;
  sr_buffer_32_1 f496(.wen(f496_wen), .wdata(f496_wdata), .clk(f496_clk), .rst(f496_rst), .rdata(f496_rdata));
  assign f496_clk = clk;
  assign f496_rst = rst;
  // Bindings to f496

  // f498
  logic [0:0] f498_wen;
  logic [31:0] f498_wdata;
  logic [0:0] f498_clk;
  logic [0:0] f498_rst;
  logic [31:0] f498_rdata;
  sr_buffer_32_1 f498(.wen(f498_wen), .wdata(f498_wdata), .clk(f498_clk), .rst(f498_rst), .rdata(f498_rdata));
  assign f498_clk = clk;
  assign f498_rst = rst;
  // Bindings to f498

  // f500
  logic [0:0] f500_wen;
  logic [31:0] f500_wdata;
  logic [0:0] f500_clk;
  logic [0:0] f500_rst;
  logic [31:0] f500_rdata;
  sr_buffer_32_1 f500(.wen(f500_wen), .wdata(f500_wdata), .clk(f500_clk), .rst(f500_rst), .rdata(f500_rdata));
  assign f500_clk = clk;
  assign f500_rst = rst;
  // Bindings to f500

  // f502
  logic [0:0] f502_wen;
  logic [31:0] f502_wdata;
  logic [0:0] f502_clk;
  logic [0:0] f502_rst;
  logic [31:0] f502_rdata;
  sr_buffer_32_1 f502(.wen(f502_wen), .wdata(f502_wdata), .clk(f502_clk), .rst(f502_rst), .rdata(f502_rdata));
  assign f502_clk = clk;
  assign f502_rst = rst;
  // Bindings to f502

  // f504
  logic [0:0] f504_wen;
  logic [31:0] f504_wdata;
  logic [0:0] f504_clk;
  logic [0:0] f504_rst;
  logic [31:0] f504_rdata;
  sr_buffer_32_1 f504(.wen(f504_wen), .wdata(f504_wdata), .clk(f504_clk), .rst(f504_rst), .rdata(f504_rdata));
  assign f504_clk = clk;
  assign f504_rst = rst;
  // Bindings to f504

  // f506
  logic [0:0] f506_wen;
  logic [31:0] f506_wdata;
  logic [0:0] f506_clk;
  logic [0:0] f506_rst;
  logic [31:0] f506_rdata;
  sr_buffer_32_1 f506(.wen(f506_wen), .wdata(f506_wdata), .clk(f506_clk), .rst(f506_rst), .rdata(f506_rdata));
  assign f506_clk = clk;
  assign f506_rst = rst;
  // Bindings to f506

  // f508
  logic [0:0] f508_wen;
  logic [31:0] f508_wdata;
  logic [0:0] f508_clk;
  logic [0:0] f508_rst;
  logic [31:0] f508_rdata;
  sr_buffer_32_1 f508(.wen(f508_wen), .wdata(f508_wdata), .clk(f508_clk), .rst(f508_rst), .rdata(f508_rdata));
  assign f508_clk = clk;
  assign f508_rst = rst;
  // Bindings to f508

  // f510
  logic [0:0] f510_wen;
  logic [31:0] f510_wdata;
  logic [0:0] f510_clk;
  logic [0:0] f510_rst;
  logic [31:0] f510_rdata;
  sr_buffer_32_1 f510(.wen(f510_wen), .wdata(f510_wdata), .clk(f510_clk), .rst(f510_rst), .rdata(f510_rdata));
  assign f510_clk = clk;
  assign f510_rst = rst;
  // Bindings to f510

  // f512
  logic [0:0] f512_wen;
  logic [31:0] f512_wdata;
  logic [0:0] f512_clk;
  logic [0:0] f512_rst;
  logic [31:0] f512_rdata;
  sr_buffer_32_1 f512(.wen(f512_wen), .wdata(f512_wdata), .clk(f512_clk), .rst(f512_rst), .rdata(f512_rdata));
  assign f512_clk = clk;
  assign f512_rst = rst;
  // Bindings to f512

  // f514
  logic [0:0] f514_wen;
  logic [31:0] f514_wdata;
  logic [0:0] f514_clk;
  logic [0:0] f514_rst;
  logic [31:0] f514_rdata;
  sr_buffer_32_1 f514(.wen(f514_wen), .wdata(f514_wdata), .clk(f514_clk), .rst(f514_rst), .rdata(f514_rdata));
  assign f514_clk = clk;
  assign f514_rst = rst;
  // Bindings to f514

  // f516
  logic [0:0] f516_wen;
  logic [31:0] f516_wdata;
  logic [0:0] f516_clk;
  logic [0:0] f516_rst;
  logic [31:0] f516_rdata;
  sr_buffer_32_1 f516(.wen(f516_wen), .wdata(f516_wdata), .clk(f516_clk), .rst(f516_rst), .rdata(f516_rdata));
  assign f516_clk = clk;
  assign f516_rst = rst;
  // Bindings to f516

  // f518
  logic [0:0] f518_wen;
  logic [31:0] f518_wdata;
  logic [0:0] f518_clk;
  logic [0:0] f518_rst;
  logic [31:0] f518_rdata;
  sr_buffer_32_1 f518(.wen(f518_wen), .wdata(f518_wdata), .clk(f518_clk), .rst(f518_rst), .rdata(f518_rdata));
  assign f518_clk = clk;
  assign f518_rst = rst;
  // Bindings to f518

  // f520
  logic [0:0] f520_wen;
  logic [31:0] f520_wdata;
  logic [0:0] f520_clk;
  logic [0:0] f520_rst;
  logic [31:0] f520_rdata;
  sr_buffer_32_1 f520(.wen(f520_wen), .wdata(f520_wdata), .clk(f520_clk), .rst(f520_rst), .rdata(f520_rdata));
  assign f520_clk = clk;
  assign f520_rst = rst;
  // Bindings to f520

  // f522
  logic [0:0] f522_wen;
  logic [31:0] f522_wdata;
  logic [0:0] f522_clk;
  logic [0:0] f522_rst;
  logic [31:0] f522_rdata;
  sr_buffer_32_1 f522(.wen(f522_wen), .wdata(f522_wdata), .clk(f522_clk), .rst(f522_rst), .rdata(f522_rdata));
  assign f522_clk = clk;
  assign f522_rst = rst;
  // Bindings to f522

  // f524
  logic [0:0] f524_wen;
  logic [31:0] f524_wdata;
  logic [0:0] f524_clk;
  logic [0:0] f524_rst;
  logic [31:0] f524_rdata;
  sr_buffer_32_1 f524(.wen(f524_wen), .wdata(f524_wdata), .clk(f524_clk), .rst(f524_rst), .rdata(f524_rdata));
  assign f524_clk = clk;
  assign f524_rst = rst;
  // Bindings to f524

  // f526
  logic [0:0] f526_wen;
  logic [31:0] f526_wdata;
  logic [0:0] f526_clk;
  logic [0:0] f526_rst;
  logic [31:0] f526_rdata;
  sr_buffer_32_1 f526(.wen(f526_wen), .wdata(f526_wdata), .clk(f526_clk), .rst(f526_rst), .rdata(f526_rdata));
  assign f526_clk = clk;
  assign f526_rst = rst;
  // Bindings to f526

  // f528
  logic [0:0] f528_wen;
  logic [31:0] f528_wdata;
  logic [0:0] f528_clk;
  logic [0:0] f528_rst;
  logic [31:0] f528_rdata;
  sr_buffer_32_1 f528(.wen(f528_wen), .wdata(f528_wdata), .clk(f528_clk), .rst(f528_rst), .rdata(f528_rdata));
  assign f528_clk = clk;
  assign f528_rst = rst;
  // Bindings to f528

  // f530
  logic [0:0] f530_wen;
  logic [31:0] f530_wdata;
  logic [0:0] f530_clk;
  logic [0:0] f530_rst;
  logic [31:0] f530_rdata;
  sr_buffer_32_1 f530(.wen(f530_wen), .wdata(f530_wdata), .clk(f530_clk), .rst(f530_rst), .rdata(f530_rdata));
  assign f530_clk = clk;
  assign f530_rst = rst;
  // Bindings to f530

  // f532
  logic [0:0] f532_wen;
  logic [31:0] f532_wdata;
  logic [0:0] f532_clk;
  logic [0:0] f532_rst;
  logic [31:0] f532_rdata;
  sr_buffer_32_1 f532(.wen(f532_wen), .wdata(f532_wdata), .clk(f532_clk), .rst(f532_rst), .rdata(f532_rdata));
  assign f532_clk = clk;
  assign f532_rst = rst;
  // Bindings to f532

  // f534
  logic [0:0] f534_wen;
  logic [31:0] f534_wdata;
  logic [0:0] f534_clk;
  logic [0:0] f534_rst;
  logic [31:0] f534_rdata;
  sr_buffer_32_1 f534(.wen(f534_wen), .wdata(f534_wdata), .clk(f534_clk), .rst(f534_rst), .rdata(f534_rdata));
  assign f534_clk = clk;
  assign f534_rst = rst;
  // Bindings to f534

  // f536
  logic [0:0] f536_wen;
  logic [31:0] f536_wdata;
  logic [0:0] f536_clk;
  logic [0:0] f536_rst;
  logic [31:0] f536_rdata;
  sr_buffer_32_1 f536(.wen(f536_wen), .wdata(f536_wdata), .clk(f536_clk), .rst(f536_rst), .rdata(f536_rdata));
  assign f536_clk = clk;
  assign f536_rst = rst;
  // Bindings to f536

  // f538
  logic [0:0] f538_wen;
  logic [31:0] f538_wdata;
  logic [0:0] f538_clk;
  logic [0:0] f538_rst;
  logic [31:0] f538_rdata;
  sr_buffer_32_1 f538(.wen(f538_wen), .wdata(f538_wdata), .clk(f538_clk), .rst(f538_rst), .rdata(f538_rdata));
  assign f538_clk = clk;
  assign f538_rst = rst;
  // Bindings to f538

  // f540
  logic [0:0] f540_wen;
  logic [31:0] f540_wdata;
  logic [0:0] f540_clk;
  logic [0:0] f540_rst;
  logic [31:0] f540_rdata;
  sr_buffer_32_1 f540(.wen(f540_wen), .wdata(f540_wdata), .clk(f540_clk), .rst(f540_rst), .rdata(f540_rdata));
  assign f540_clk = clk;
  assign f540_rst = rst;
  // Bindings to f540

  // f542
  logic [0:0] f542_wen;
  logic [31:0] f542_wdata;
  logic [0:0] f542_clk;
  logic [0:0] f542_rst;
  logic [31:0] f542_rdata;
  sr_buffer_32_1 f542(.wen(f542_wen), .wdata(f542_wdata), .clk(f542_clk), .rst(f542_rst), .rdata(f542_rdata));
  assign f542_clk = clk;
  assign f542_rst = rst;
  // Bindings to f542

  // f544
  logic [0:0] f544_wen;
  logic [31:0] f544_wdata;
  logic [0:0] f544_clk;
  logic [0:0] f544_rst;
  logic [31:0] f544_rdata;
  sr_buffer_32_1 f544(.wen(f544_wen), .wdata(f544_wdata), .clk(f544_clk), .rst(f544_rst), .rdata(f544_rdata));
  assign f544_clk = clk;
  assign f544_rst = rst;
  // Bindings to f544

  // f546
  logic [0:0] f546_wen;
  logic [31:0] f546_wdata;
  logic [0:0] f546_clk;
  logic [0:0] f546_rst;
  logic [31:0] f546_rdata;
  sr_buffer_32_1 f546(.wen(f546_wen), .wdata(f546_wdata), .clk(f546_clk), .rst(f546_rst), .rdata(f546_rdata));
  assign f546_clk = clk;
  assign f546_rst = rst;
  // Bindings to f546

  // f548
  logic [0:0] f548_wen;
  logic [31:0] f548_wdata;
  logic [0:0] f548_clk;
  logic [0:0] f548_rst;
  logic [31:0] f548_rdata;
  sr_buffer_32_1 f548(.wen(f548_wen), .wdata(f548_wdata), .clk(f548_clk), .rst(f548_rst), .rdata(f548_rdata));
  assign f548_clk = clk;
  assign f548_rst = rst;
  // Bindings to f548

  // f550
  logic [0:0] f550_wen;
  logic [31:0] f550_wdata;
  logic [0:0] f550_clk;
  logic [0:0] f550_rst;
  logic [31:0] f550_rdata;
  sr_buffer_32_1 f550(.wen(f550_wen), .wdata(f550_wdata), .clk(f550_clk), .rst(f550_rst), .rdata(f550_rdata));
  assign f550_clk = clk;
  assign f550_rst = rst;
  // Bindings to f550

  // f552
  logic [0:0] f552_wen;
  logic [31:0] f552_wdata;
  logic [0:0] f552_clk;
  logic [0:0] f552_rst;
  logic [31:0] f552_rdata;
  sr_buffer_32_1 f552(.wen(f552_wen), .wdata(f552_wdata), .clk(f552_clk), .rst(f552_rst), .rdata(f552_rdata));
  assign f552_clk = clk;
  assign f552_rst = rst;
  // Bindings to f552

  // f554
  logic [0:0] f554_wen;
  logic [31:0] f554_wdata;
  logic [0:0] f554_clk;
  logic [0:0] f554_rst;
  logic [31:0] f554_rdata;
  sr_buffer_32_1 f554(.wen(f554_wen), .wdata(f554_wdata), .clk(f554_clk), .rst(f554_rst), .rdata(f554_rdata));
  assign f554_clk = clk;
  assign f554_rst = rst;
  // Bindings to f554

  // f556
  logic [0:0] f556_wen;
  logic [31:0] f556_wdata;
  logic [0:0] f556_clk;
  logic [0:0] f556_rst;
  logic [31:0] f556_rdata;
  sr_buffer_32_1 f556(.wen(f556_wen), .wdata(f556_wdata), .clk(f556_clk), .rst(f556_rst), .rdata(f556_rdata));
  assign f556_clk = clk;
  assign f556_rst = rst;
  // Bindings to f556

  // f558
  logic [0:0] f558_wen;
  logic [31:0] f558_wdata;
  logic [0:0] f558_clk;
  logic [0:0] f558_rst;
  logic [31:0] f558_rdata;
  sr_buffer_32_1 f558(.wen(f558_wen), .wdata(f558_wdata), .clk(f558_clk), .rst(f558_rst), .rdata(f558_rdata));
  assign f558_clk = clk;
  assign f558_rst = rst;
  // Bindings to f558

  // f560
  logic [0:0] f560_wen;
  logic [31:0] f560_wdata;
  logic [0:0] f560_clk;
  logic [0:0] f560_rst;
  logic [31:0] f560_rdata;
  sr_buffer_32_1 f560(.wen(f560_wen), .wdata(f560_wdata), .clk(f560_clk), .rst(f560_rst), .rdata(f560_rdata));
  assign f560_clk = clk;
  assign f560_rst = rst;
  // Bindings to f560

  // f562
  logic [0:0] f562_wen;
  logic [31:0] f562_wdata;
  logic [0:0] f562_clk;
  logic [0:0] f562_rst;
  logic [31:0] f562_rdata;
  sr_buffer_32_1 f562(.wen(f562_wen), .wdata(f562_wdata), .clk(f562_clk), .rst(f562_rst), .rdata(f562_rdata));
  assign f562_clk = clk;
  assign f562_rst = rst;
  // Bindings to f562

  // f564
  logic [0:0] f564_wen;
  logic [31:0] f564_wdata;
  logic [0:0] f564_clk;
  logic [0:0] f564_rst;
  logic [31:0] f564_rdata;
  sr_buffer_32_1 f564(.wen(f564_wen), .wdata(f564_wdata), .clk(f564_clk), .rst(f564_rst), .rdata(f564_rdata));
  assign f564_clk = clk;
  assign f564_rst = rst;
  // Bindings to f564

  // f566
  logic [0:0] f566_wen;
  logic [31:0] f566_wdata;
  logic [0:0] f566_clk;
  logic [0:0] f566_rst;
  logic [31:0] f566_rdata;
  sr_buffer_32_1 f566(.wen(f566_wen), .wdata(f566_wdata), .clk(f566_clk), .rst(f566_rst), .rdata(f566_rdata));
  assign f566_clk = clk;
  assign f566_rst = rst;
  // Bindings to f566

  // f568
  logic [0:0] f568_wen;
  logic [31:0] f568_wdata;
  logic [0:0] f568_clk;
  logic [0:0] f568_rst;
  logic [31:0] f568_rdata;
  sr_buffer_32_1 f568(.wen(f568_wen), .wdata(f568_wdata), .clk(f568_clk), .rst(f568_rst), .rdata(f568_rdata));
  assign f568_clk = clk;
  assign f568_rst = rst;
  // Bindings to f568

  // f570
  logic [0:0] f570_wen;
  logic [31:0] f570_wdata;
  logic [0:0] f570_clk;
  logic [0:0] f570_rst;
  logic [31:0] f570_rdata;
  sr_buffer_32_1 f570(.wen(f570_wen), .wdata(f570_wdata), .clk(f570_clk), .rst(f570_rst), .rdata(f570_rdata));
  assign f570_clk = clk;
  assign f570_rst = rst;
  // Bindings to f570

  // f572
  logic [0:0] f572_wen;
  logic [31:0] f572_wdata;
  logic [0:0] f572_clk;
  logic [0:0] f572_rst;
  logic [31:0] f572_rdata;
  sr_buffer_32_1 f572(.wen(f572_wen), .wdata(f572_wdata), .clk(f572_clk), .rst(f572_rst), .rdata(f572_rdata));
  assign f572_clk = clk;
  assign f572_rst = rst;
  // Bindings to f572

  // f574
  logic [0:0] f574_wen;
  logic [31:0] f574_wdata;
  logic [0:0] f574_clk;
  logic [0:0] f574_rst;
  logic [31:0] f574_rdata;
  sr_buffer_32_1 f574(.wen(f574_wen), .wdata(f574_wdata), .clk(f574_clk), .rst(f574_rst), .rdata(f574_rdata));
  assign f574_clk = clk;
  assign f574_rst = rst;
  // Bindings to f574

  // f576
  logic [0:0] f576_wen;
  logic [31:0] f576_wdata;
  logic [0:0] f576_clk;
  logic [0:0] f576_rst;
  logic [31:0] f576_rdata;
  sr_buffer_32_1 f576(.wen(f576_wen), .wdata(f576_wdata), .clk(f576_clk), .rst(f576_rst), .rdata(f576_rdata));
  assign f576_clk = clk;
  assign f576_rst = rst;
  // Bindings to f576

  // f578
  logic [0:0] f578_wen;
  logic [31:0] f578_wdata;
  logic [0:0] f578_clk;
  logic [0:0] f578_rst;
  logic [31:0] f578_rdata;
  sr_buffer_32_1 f578(.wen(f578_wen), .wdata(f578_wdata), .clk(f578_clk), .rst(f578_rst), .rdata(f578_rdata));
  assign f578_clk = clk;
  assign f578_rst = rst;
  // Bindings to f578

  // f580
  logic [0:0] f580_wen;
  logic [31:0] f580_wdata;
  logic [0:0] f580_clk;
  logic [0:0] f580_rst;
  logic [31:0] f580_rdata;
  sr_buffer_32_1 f580(.wen(f580_wen), .wdata(f580_wdata), .clk(f580_clk), .rst(f580_rst), .rdata(f580_rdata));
  assign f580_clk = clk;
  assign f580_rst = rst;
  // Bindings to f580

  // f582
  logic [0:0] f582_wen;
  logic [31:0] f582_wdata;
  logic [0:0] f582_clk;
  logic [0:0] f582_rst;
  logic [31:0] f582_rdata;
  sr_buffer_32_1 f582(.wen(f582_wen), .wdata(f582_wdata), .clk(f582_clk), .rst(f582_rst), .rdata(f582_rdata));
  assign f582_clk = clk;
  assign f582_rst = rst;
  // Bindings to f582

  // f584
  logic [0:0] f584_wen;
  logic [31:0] f584_wdata;
  logic [0:0] f584_clk;
  logic [0:0] f584_rst;
  logic [31:0] f584_rdata;
  sr_buffer_32_1 f584(.wen(f584_wen), .wdata(f584_wdata), .clk(f584_clk), .rst(f584_rst), .rdata(f584_rdata));
  assign f584_clk = clk;
  assign f584_rst = rst;
  // Bindings to f584

  // f586
  logic [0:0] f586_wen;
  logic [31:0] f586_wdata;
  logic [0:0] f586_clk;
  logic [0:0] f586_rst;
  logic [31:0] f586_rdata;
  sr_buffer_32_1 f586(.wen(f586_wen), .wdata(f586_wdata), .clk(f586_clk), .rst(f586_rst), .rdata(f586_rdata));
  assign f586_clk = clk;
  assign f586_rst = rst;
  // Bindings to f586

  // f588
  logic [0:0] f588_wen;
  logic [31:0] f588_wdata;
  logic [0:0] f588_clk;
  logic [0:0] f588_rst;
  logic [31:0] f588_rdata;
  sr_buffer_32_1 f588(.wen(f588_wen), .wdata(f588_wdata), .clk(f588_clk), .rst(f588_rst), .rdata(f588_rdata));
  assign f588_clk = clk;
  assign f588_rst = rst;
  // Bindings to f588

  // f590
  logic [0:0] f590_wen;
  logic [31:0] f590_wdata;
  logic [0:0] f590_clk;
  logic [0:0] f590_rst;
  logic [31:0] f590_rdata;
  sr_buffer_32_1 f590(.wen(f590_wen), .wdata(f590_wdata), .clk(f590_clk), .rst(f590_rst), .rdata(f590_rdata));
  assign f590_clk = clk;
  assign f590_rst = rst;
  // Bindings to f590

  // f592
  logic [0:0] f592_wen;
  logic [31:0] f592_wdata;
  logic [0:0] f592_clk;
  logic [0:0] f592_rst;
  logic [31:0] f592_rdata;
  sr_buffer_32_1 f592(.wen(f592_wen), .wdata(f592_wdata), .clk(f592_clk), .rst(f592_rst), .rdata(f592_rdata));
  assign f592_clk = clk;
  assign f592_rst = rst;
  // Bindings to f592

  // f594
  logic [0:0] f594_wen;
  logic [31:0] f594_wdata;
  logic [0:0] f594_clk;
  logic [0:0] f594_rst;
  logic [31:0] f594_rdata;
  sr_buffer_32_1 f594(.wen(f594_wen), .wdata(f594_wdata), .clk(f594_clk), .rst(f594_rst), .rdata(f594_rdata));
  assign f594_clk = clk;
  assign f594_rst = rst;
  // Bindings to f594

  // f596
  logic [0:0] f596_wen;
  logic [31:0] f596_wdata;
  logic [0:0] f596_clk;
  logic [0:0] f596_rst;
  logic [31:0] f596_rdata;
  sr_buffer_32_1 f596(.wen(f596_wen), .wdata(f596_wdata), .clk(f596_clk), .rst(f596_rst), .rdata(f596_rdata));
  assign f596_clk = clk;
  assign f596_rst = rst;
  // Bindings to f596

  // f598
  logic [0:0] f598_wen;
  logic [31:0] f598_wdata;
  logic [0:0] f598_clk;
  logic [0:0] f598_rst;
  logic [31:0] f598_rdata;
  sr_buffer_32_1 f598(.wen(f598_wen), .wdata(f598_wdata), .clk(f598_clk), .rst(f598_rst), .rdata(f598_rdata));
  assign f598_clk = clk;
  assign f598_rst = rst;
  // Bindings to f598

  // f600
  logic [0:0] f600_wen;
  logic [31:0] f600_wdata;
  logic [0:0] f600_clk;
  logic [0:0] f600_rst;
  logic [31:0] f600_rdata;
  sr_buffer_32_1 f600(.wen(f600_wen), .wdata(f600_wdata), .clk(f600_clk), .rst(f600_rst), .rdata(f600_rdata));
  assign f600_clk = clk;
  assign f600_rst = rst;
  // Bindings to f600

  // f602
  logic [0:0] f602_wen;
  logic [31:0] f602_wdata;
  logic [0:0] f602_clk;
  logic [0:0] f602_rst;
  logic [31:0] f602_rdata;
  sr_buffer_32_1 f602(.wen(f602_wen), .wdata(f602_wdata), .clk(f602_clk), .rst(f602_rst), .rdata(f602_rdata));
  assign f602_clk = clk;
  assign f602_rst = rst;
  // Bindings to f602

  // f604
  logic [0:0] f604_wen;
  logic [31:0] f604_wdata;
  logic [0:0] f604_clk;
  logic [0:0] f604_rst;
  logic [31:0] f604_rdata;
  sr_buffer_32_1 f604(.wen(f604_wen), .wdata(f604_wdata), .clk(f604_clk), .rst(f604_rst), .rdata(f604_rdata));
  assign f604_clk = clk;
  assign f604_rst = rst;
  // Bindings to f604

  // f606
  logic [0:0] f606_wen;
  logic [31:0] f606_wdata;
  logic [0:0] f606_clk;
  logic [0:0] f606_rst;
  logic [31:0] f606_rdata;
  sr_buffer_32_1 f606(.wen(f606_wen), .wdata(f606_wdata), .clk(f606_clk), .rst(f606_rst), .rdata(f606_rdata));
  assign f606_clk = clk;
  assign f606_rst = rst;
  // Bindings to f606

  // f608
  logic [0:0] f608_wen;
  logic [31:0] f608_wdata;
  logic [0:0] f608_clk;
  logic [0:0] f608_rst;
  logic [31:0] f608_rdata;
  sr_buffer_32_1 f608(.wen(f608_wen), .wdata(f608_wdata), .clk(f608_clk), .rst(f608_rst), .rdata(f608_rdata));
  assign f608_clk = clk;
  assign f608_rst = rst;
  // Bindings to f608

  // f610
  logic [0:0] f610_wen;
  logic [31:0] f610_wdata;
  logic [0:0] f610_clk;
  logic [0:0] f610_rst;
  logic [31:0] f610_rdata;
  sr_buffer_32_1 f610(.wen(f610_wen), .wdata(f610_wdata), .clk(f610_clk), .rst(f610_rst), .rdata(f610_rdata));
  assign f610_clk = clk;
  assign f610_rst = rst;
  // Bindings to f610

  // f612
  logic [0:0] f612_wen;
  logic [31:0] f612_wdata;
  logic [0:0] f612_clk;
  logic [0:0] f612_rst;
  logic [31:0] f612_rdata;
  sr_buffer_32_1 f612(.wen(f612_wen), .wdata(f612_wdata), .clk(f612_clk), .rst(f612_rst), .rdata(f612_rdata));
  assign f612_clk = clk;
  assign f612_rst = rst;
  // Bindings to f612

  // f614
  logic [0:0] f614_wen;
  logic [31:0] f614_wdata;
  logic [0:0] f614_clk;
  logic [0:0] f614_rst;
  logic [31:0] f614_rdata;
  sr_buffer_32_1 f614(.wen(f614_wen), .wdata(f614_wdata), .clk(f614_clk), .rst(f614_rst), .rdata(f614_rdata));
  assign f614_clk = clk;
  assign f614_rst = rst;
  // Bindings to f614

  // f616
  logic [0:0] f616_wen;
  logic [31:0] f616_wdata;
  logic [0:0] f616_clk;
  logic [0:0] f616_rst;
  logic [31:0] f616_rdata;
  sr_buffer_32_1 f616(.wen(f616_wen), .wdata(f616_wdata), .clk(f616_clk), .rst(f616_rst), .rdata(f616_rdata));
  assign f616_clk = clk;
  assign f616_rst = rst;
  // Bindings to f616

  // f618
  logic [0:0] f618_wen;
  logic [31:0] f618_wdata;
  logic [0:0] f618_clk;
  logic [0:0] f618_rst;
  logic [31:0] f618_rdata;
  sr_buffer_32_1 f618(.wen(f618_wen), .wdata(f618_wdata), .clk(f618_clk), .rst(f618_rst), .rdata(f618_rdata));
  assign f618_clk = clk;
  assign f618_rst = rst;
  // Bindings to f618

  // f620
  logic [0:0] f620_wen;
  logic [31:0] f620_wdata;
  logic [0:0] f620_clk;
  logic [0:0] f620_rst;
  logic [31:0] f620_rdata;
  sr_buffer_32_1 f620(.wen(f620_wen), .wdata(f620_wdata), .clk(f620_clk), .rst(f620_rst), .rdata(f620_rdata));
  assign f620_clk = clk;
  assign f620_rst = rst;
  // Bindings to f620

  // f622
  logic [0:0] f622_wen;
  logic [31:0] f622_wdata;
  logic [0:0] f622_clk;
  logic [0:0] f622_rst;
  logic [31:0] f622_rdata;
  sr_buffer_32_1 f622(.wen(f622_wen), .wdata(f622_wdata), .clk(f622_clk), .rst(f622_rst), .rdata(f622_rdata));
  assign f622_clk = clk;
  assign f622_rst = rst;
  // Bindings to f622

  // f624
  logic [0:0] f624_wen;
  logic [31:0] f624_wdata;
  logic [0:0] f624_clk;
  logic [0:0] f624_rst;
  logic [31:0] f624_rdata;
  sr_buffer_32_1 f624(.wen(f624_wen), .wdata(f624_wdata), .clk(f624_clk), .rst(f624_rst), .rdata(f624_rdata));
  assign f624_clk = clk;
  assign f624_rst = rst;
  // Bindings to f624



endmodule


module in_wire_final_merged_2_update_0_write_wen(output [0:0] final_merged_2_update_0_write_wen);

endmodule


module in_wire_final_merged_2_update_0_write_wdata(output [31:0] final_merged_2_update_0_write_wdata);

endmodule


module in_wire_in_update_0_write_wen(output [0:0] in_update_0_write_wen);

endmodule


module dark_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module bright_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_in_update_0_write_wdata(output [31:0] in_update_0_write_wdata);

endmodule


module in_wire_bright_update_0_read_dummy(output [31:0] bright_update_0_read_dummy);

endmodule


module out_wire_bright_update_0_read_rdata(input [31:0] bright_update_0_read_rdata);

endmodule


module in_wire_dark_update_0_read_dummy(output [31:0] dark_update_0_read_dummy);

endmodule


module out_wire_dark_update_0_read_rdata(input [31:0] dark_update_0_read_rdata);

endmodule


module in_wire_pyramid_synthetic_exposure_fusion_update_0_write_wen(output [0:0] pyramid_synthetic_exposure_fusion_update_0_write_wen);

endmodule


module in_off_chip(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] in_update_0_read_dummy, output [31:0] in_update_0_read_rdata, input [0:0] in_off_chip_update_0_write_wen, input [31:0] in_off_chip_update_0_write_wdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to in_update_0_read_dummy
    // rd_2
  assign rd_2 = in_update_0_read_dummy;

  // Bindings to in_update_0_read_rdata
    // wr_3
  assign in_update_0_read_rdata = rd_2;

  // Bindings to in_off_chip_update_0_write_wen
    // rd_0
  assign rd_0 = in_off_chip_update_0_write_wen;

  // Bindings to in_off_chip_update_0_write_wdata
    // rd_1
  assign rd_1 = in_off_chip_update_0_write_wdata;



endmodule


module in_wire_pyramid_synthetic_exposure_fusion_update_0_write_wdata(output [31:0] pyramid_synthetic_exposure_fusion_update_0_write_wdata);

endmodule


module bright_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_gauss_blur_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_weights_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_gauss_blur_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module dark_gauss_ds_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module dark_gauss_blur_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_gauss_ds_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module weight_sums_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_gauss_blur_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module final_merged_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module fused_level_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module final_merged_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module final_merged_0_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module pyramid_synthetic_exposure_fusion_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module dark_gauss_blur_2_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (627 - d0 >= 0) ? (1262) : (-628 + d0 == 0) ? (1262) : 0;
    end
  end

endmodule


module dark_laplace_us_0_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (-1 + d1 == 0) ? ((4416 - floord(d0, 2))) : (d1 == 0) ? (3792) : ((-1 - d1) % 2 == 0 && -3 + d1 >= 0) ? ((4416 - floord(d0, 2))) : ((-d1) % 2 == 0 && -2 + d1 >= 0) ? (3792) : 0;
    end
  end

endmodule


module dark_gauss_blur_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1264;
    end
  end

endmodule


module dark_gauss_blur_2_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module dark_gauss_blur_2_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 633;
    end
  end

endmodule


module dark_gauss_blur_2_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1263;
    end
  end

endmodule


module dark_gauss_blur_2_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 632;
    end
  end

endmodule


module dark_gauss_blur_2_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module dark_gauss_blur_2_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_gauss_ds_1_update_0_write_wen(output [0:0] dark_gauss_ds_1_update_0_write_wen);

endmodule


module in_wire_dark_gauss_ds_1_update_0_write_wdata(output [31:0] dark_gauss_ds_1_update_0_write_wdata);

endmodule


module dark_gauss_blur_2_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (627 - d0 >= 0) ? (631) : (-628 + d0 == 0) ? (631) : 0;
    end
  end

endmodule


module dark_gauss_ds_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_gauss_ds_2_update_0_write_wen, output [31:0] dark_laplace_us_1_update_0_read_rdata, input [31:0] dark_laplace_us_1_update_0_read_dummy, output [31:0] dark_laplace_diff_2_update_0_read_rdata, input [31:0] dark_laplace_diff_2_update_0_read_dummy, output [287:0] dark_gauss_blur_3_update_0_read_rdata, input [287:0] dark_gauss_blur_3_update_0_read_dummy, input [31:0] dark_gauss_ds_2_update_0_write_wdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;
  logic [31:0] rd_4;
  logic [31:0] rd_6;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;
  reg [31:0] rd_6_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;
      rd_6_stage_1 <= rd_6;


    end

  end


  // Data processing units...
  // selector_dark_laplace_us_1_rd0_select
  logic [0:0] selector_dark_laplace_us_1_rd0_select_clk;
  logic [0:0] selector_dark_laplace_us_1_rd0_select_rst;
  logic [31:0] selector_dark_laplace_us_1_rd0_select_d0;
  logic [31:0] selector_dark_laplace_us_1_rd0_select_d1;
  logic [31:0] selector_dark_laplace_us_1_rd0_select_out;
  dark_laplace_us_1_rd0_select selector_dark_laplace_us_1_rd0_select(.clk(selector_dark_laplace_us_1_rd0_select_clk), .rst(selector_dark_laplace_us_1_rd0_select_rst), .d0(selector_dark_laplace_us_1_rd0_select_d0), .d1(selector_dark_laplace_us_1_rd0_select_d1), .out(selector_dark_laplace_us_1_rd0_select_out));
  assign selector_dark_laplace_us_1_rd0_select_clk = clk;
  assign selector_dark_laplace_us_1_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_us_1_rd0_select

  // selector_dark_gauss_blur_3_rd8_select
  logic [0:0] selector_dark_gauss_blur_3_rd8_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd8_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd8_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd8_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd8_select_out;
  dark_gauss_blur_3_rd8_select selector_dark_gauss_blur_3_rd8_select(.clk(selector_dark_gauss_blur_3_rd8_select_clk), .rst(selector_dark_gauss_blur_3_rd8_select_rst), .d0(selector_dark_gauss_blur_3_rd8_select_d0), .d1(selector_dark_gauss_blur_3_rd8_select_d1), .out(selector_dark_gauss_blur_3_rd8_select_out));
  assign selector_dark_gauss_blur_3_rd8_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd8_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd8_select

  // selector_dark_gauss_blur_3_rd3_select
  logic [0:0] selector_dark_gauss_blur_3_rd3_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd3_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd3_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd3_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd3_select_out;
  dark_gauss_blur_3_rd3_select selector_dark_gauss_blur_3_rd3_select(.clk(selector_dark_gauss_blur_3_rd3_select_clk), .rst(selector_dark_gauss_blur_3_rd3_select_rst), .d0(selector_dark_gauss_blur_3_rd3_select_d0), .d1(selector_dark_gauss_blur_3_rd3_select_d1), .out(selector_dark_gauss_blur_3_rd3_select_out));
  assign selector_dark_gauss_blur_3_rd3_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd3_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd3_select

  // selector_dark_gauss_blur_3_rd0_select
  logic [0:0] selector_dark_gauss_blur_3_rd0_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd0_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd0_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd0_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd0_select_out;
  dark_gauss_blur_3_rd0_select selector_dark_gauss_blur_3_rd0_select(.clk(selector_dark_gauss_blur_3_rd0_select_clk), .rst(selector_dark_gauss_blur_3_rd0_select_rst), .d0(selector_dark_gauss_blur_3_rd0_select_d0), .d1(selector_dark_gauss_blur_3_rd0_select_d1), .out(selector_dark_gauss_blur_3_rd0_select_out));
  assign selector_dark_gauss_blur_3_rd0_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd0_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd0_select

  // selector_dark_gauss_blur_3_rd1_select
  logic [0:0] selector_dark_gauss_blur_3_rd1_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd1_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd1_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd1_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd1_select_out;
  dark_gauss_blur_3_rd1_select selector_dark_gauss_blur_3_rd1_select(.clk(selector_dark_gauss_blur_3_rd1_select_clk), .rst(selector_dark_gauss_blur_3_rd1_select_rst), .d0(selector_dark_gauss_blur_3_rd1_select_d0), .d1(selector_dark_gauss_blur_3_rd1_select_d1), .out(selector_dark_gauss_blur_3_rd1_select_out));
  assign selector_dark_gauss_blur_3_rd1_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd1_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd1_select

  // dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_clk;
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_rst;
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_start;
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_done;
  dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10 dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10(.clk(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_clk), .rst(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_rst), .start(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_start), .done(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_done));
  assign dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_clk = clk;
  assign dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10

  // Bindings to dark_gauss_ds_2_update_0_write_wen
    // rd_0
  assign rd_0 = dark_gauss_ds_2_update_0_write_wen;

  // selector_dark_gauss_blur_3_rd2_select
  logic [0:0] selector_dark_gauss_blur_3_rd2_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd2_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd2_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd2_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd2_select_out;
  dark_gauss_blur_3_rd2_select selector_dark_gauss_blur_3_rd2_select(.clk(selector_dark_gauss_blur_3_rd2_select_clk), .rst(selector_dark_gauss_blur_3_rd2_select_rst), .d0(selector_dark_gauss_blur_3_rd2_select_d0), .d1(selector_dark_gauss_blur_3_rd2_select_d1), .out(selector_dark_gauss_blur_3_rd2_select_out));
  assign selector_dark_gauss_blur_3_rd2_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd2_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd2_select

  // selector_dark_laplace_diff_2_rd0_select
  logic [0:0] selector_dark_laplace_diff_2_rd0_select_clk;
  logic [0:0] selector_dark_laplace_diff_2_rd0_select_rst;
  logic [31:0] selector_dark_laplace_diff_2_rd0_select_d0;
  logic [31:0] selector_dark_laplace_diff_2_rd0_select_d1;
  logic [31:0] selector_dark_laplace_diff_2_rd0_select_out;
  dark_laplace_diff_2_rd0_select selector_dark_laplace_diff_2_rd0_select(.clk(selector_dark_laplace_diff_2_rd0_select_clk), .rst(selector_dark_laplace_diff_2_rd0_select_rst), .d0(selector_dark_laplace_diff_2_rd0_select_d0), .d1(selector_dark_laplace_diff_2_rd0_select_d1), .out(selector_dark_laplace_diff_2_rd0_select_out));
  assign selector_dark_laplace_diff_2_rd0_select_clk = clk;
  assign selector_dark_laplace_diff_2_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_diff_2_rd0_select

  // selector_dark_gauss_blur_3_rd7_select
  logic [0:0] selector_dark_gauss_blur_3_rd7_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd7_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd7_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd7_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd7_select_out;
  dark_gauss_blur_3_rd7_select selector_dark_gauss_blur_3_rd7_select(.clk(selector_dark_gauss_blur_3_rd7_select_clk), .rst(selector_dark_gauss_blur_3_rd7_select_rst), .d0(selector_dark_gauss_blur_3_rd7_select_d0), .d1(selector_dark_gauss_blur_3_rd7_select_d1), .out(selector_dark_gauss_blur_3_rd7_select_out));
  assign selector_dark_gauss_blur_3_rd7_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd7_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd7_select

  // selector_dark_gauss_blur_3_rd6_select
  logic [0:0] selector_dark_gauss_blur_3_rd6_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd6_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd6_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd6_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd6_select_out;
  dark_gauss_blur_3_rd6_select selector_dark_gauss_blur_3_rd6_select(.clk(selector_dark_gauss_blur_3_rd6_select_clk), .rst(selector_dark_gauss_blur_3_rd6_select_rst), .d0(selector_dark_gauss_blur_3_rd6_select_d0), .d1(selector_dark_gauss_blur_3_rd6_select_d1), .out(selector_dark_gauss_blur_3_rd6_select_out));
  assign selector_dark_gauss_blur_3_rd6_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd6_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd6_select

  // selector_dark_gauss_blur_3_rd5_select
  logic [0:0] selector_dark_gauss_blur_3_rd5_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd5_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd5_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd5_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd5_select_out;
  dark_gauss_blur_3_rd5_select selector_dark_gauss_blur_3_rd5_select(.clk(selector_dark_gauss_blur_3_rd5_select_clk), .rst(selector_dark_gauss_blur_3_rd5_select_rst), .d0(selector_dark_gauss_blur_3_rd5_select_d0), .d1(selector_dark_gauss_blur_3_rd5_select_d1), .out(selector_dark_gauss_blur_3_rd5_select_out));
  assign selector_dark_gauss_blur_3_rd5_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd5_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd5_select

  // selector_dark_gauss_blur_3_rd4_select
  logic [0:0] selector_dark_gauss_blur_3_rd4_select_clk;
  logic [0:0] selector_dark_gauss_blur_3_rd4_select_rst;
  logic [31:0] selector_dark_gauss_blur_3_rd4_select_d0;
  logic [31:0] selector_dark_gauss_blur_3_rd4_select_d1;
  logic [31:0] selector_dark_gauss_blur_3_rd4_select_out;
  dark_gauss_blur_3_rd4_select selector_dark_gauss_blur_3_rd4_select(.clk(selector_dark_gauss_blur_3_rd4_select_clk), .rst(selector_dark_gauss_blur_3_rd4_select_rst), .d0(selector_dark_gauss_blur_3_rd4_select_d0), .d1(selector_dark_gauss_blur_3_rd4_select_d1), .out(selector_dark_gauss_blur_3_rd4_select_out));
  assign selector_dark_gauss_blur_3_rd4_select_clk = clk;
  assign selector_dark_gauss_blur_3_rd4_select_rst = rst;
  // Bindings to selector_dark_gauss_blur_3_rd4_select

  // dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_clk;
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_rst;
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_start;
  logic [0:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_done;
  dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0 dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0(.clk(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_clk), .rst(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_rst), .start(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_start), .done(dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_done));
  assign dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_clk = clk;
  assign dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0_rst = rst;
  // Bindings to dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_to_dark_laplace_us_1_rd0

  // Bindings to dark_laplace_us_1_update_0_read_rdata
    // wr_7
  assign dark_laplace_us_1_update_0_read_rdata = rd_6;

  // Bindings to dark_laplace_us_1_update_0_read_dummy
    // rd_6
  assign rd_6 = dark_laplace_us_1_update_0_read_dummy;

  // Bindings to dark_laplace_diff_2_update_0_read_rdata
    // wr_5
  assign dark_laplace_diff_2_update_0_read_rdata = rd_4;

  // Bindings to dark_laplace_diff_2_update_0_read_dummy
    // rd_4
  assign rd_4 = dark_laplace_diff_2_update_0_read_dummy;

  // Bindings to dark_gauss_blur_3_update_0_read_rdata
    // wr_3
  assign dark_gauss_blur_3_update_0_read_rdata = rd_2;

  // Bindings to dark_gauss_blur_3_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_gauss_blur_3_update_0_read_dummy;

  // Bindings to dark_gauss_ds_2_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_gauss_ds_2_update_0_write_wdata;



endmodule


module in_wire_dark_gauss_blur_2_update_0_read_dummy(output [287:0] dark_gauss_blur_2_update_0_read_dummy);

endmodule


module out_wire_dark_gauss_blur_2_update_0_read_rdata(input [287:0] dark_gauss_blur_2_update_0_read_rdata);

endmodule


module in_wire_dark_laplace_diff_1_update_0_read_dummy(output [31:0] dark_laplace_diff_1_update_0_read_dummy);

endmodule


module out_wire_dark_laplace_diff_1_update_0_read_rdata(input [31:0] dark_laplace_diff_1_update_0_read_rdata);

endmodule


module in_wire_dark_laplace_us_0_update_0_read_dummy(output [31:0] dark_laplace_us_0_update_0_read_dummy);

endmodule


module out_wire_dark_laplace_us_0_update_0_read_rdata(input [31:0] dark_laplace_us_0_update_0_read_rdata);

endmodule


module dark_gauss_ds_2_dark_gauss_ds_2_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_312 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_312 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16



endmodule


module dark_gauss_blur_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 632;
    end
  end

endmodule


module dark_gauss_blur_3_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (311 - d0 >= 0) ? (630) : (-312 + d0 == 0) ? (630) : 0;
    end
  end

endmodule


module dark_gauss_blur_3_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 317;
    end
  end

endmodule


module dark_gauss_blur_3_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module dark_gauss_blur_3_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 631;
    end
  end

endmodule


module dark_gauss_blur_3_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 316;
    end
  end

endmodule


module dark_gauss_blur_3_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module dark_gauss_blur_3_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_laplace_us_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (-1 + d1 == 0) ? ((944 - floord(d0, 2))) : (d1 == 0) ? (632) : ((-1 - d1) % 2 == 0 && -3 + d1 >= 0) ? ((944 - floord(d0, 2))) : ((-d1) % 2 == 0 && -2 + d1 >= 0) ? (632) : 0;
    end
  end

endmodule


module dark_gauss_blur_3_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (311 - d0 >= 0) ? (315) : (-312 + d0 == 0) ? (315) : 0;
    end
  end

endmodule


module in_wire_dark_laplace_diff_0_update_0_write_wdata(output [31:0] dark_laplace_diff_0_update_0_write_wdata);

endmodule


module in_wire_dark_laplace_diff_0_update_0_write_wen(output [0:0] dark_laplace_diff_0_update_0_write_wen);

endmodule


module dark_weights_normed_gauss_blur_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] dark_weights_normed_gauss_ds_1_update_0_read_rdata, input [31:0] dark_weights_normed_gauss_ds_1_update_0_read_dummy, input [31:0] dark_weights_normed_gauss_blur_1_update_0_write_wdata, input [0:0] dark_weights_normed_gauss_blur_1_update_0_write_wen);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_weights_normed_gauss_ds_1_update_0_read_rdata
    // wr_3
  assign dark_weights_normed_gauss_ds_1_update_0_read_rdata = rd_2;

  // Bindings to dark_weights_normed_gauss_ds_1_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_weights_normed_gauss_ds_1_update_0_read_dummy;

  // Bindings to dark_weights_normed_gauss_blur_1_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_normed_gauss_blur_1_update_0_write_wdata;

  // selector_dark_weights_normed_gauss_ds_1_rd0_select
  logic [0:0] selector_dark_weights_normed_gauss_ds_1_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_ds_1_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_ds_1_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_ds_1_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_ds_1_rd0_select_out;
  dark_weights_normed_gauss_ds_1_rd0_select selector_dark_weights_normed_gauss_ds_1_rd0_select(.clk(selector_dark_weights_normed_gauss_ds_1_rd0_select_clk), .rst(selector_dark_weights_normed_gauss_ds_1_rd0_select_rst), .d0(selector_dark_weights_normed_gauss_ds_1_rd0_select_d0), .d1(selector_dark_weights_normed_gauss_ds_1_rd0_select_d1), .out(selector_dark_weights_normed_gauss_ds_1_rd0_select_out));
  assign selector_dark_weights_normed_gauss_ds_1_rd0_select_clk = clk;
  assign selector_dark_weights_normed_gauss_ds_1_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_ds_1_rd0_select

  // Bindings to dark_weights_normed_gauss_blur_1_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_normed_gauss_blur_1_update_0_write_wen;

  // dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1
  logic [0:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_done;
  dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1 dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1(.clk(dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_clk), .rst(dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_rst), .start(dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_start), .done(dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_done));
  assign dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_clk = clk;
  assign dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write0_merged_banks_1



endmodule


module in_wire_dark_weights_normed_gauss_blur_2_update_0_write_wen(output [0:0] dark_weights_normed_gauss_blur_2_update_0_write_wen);

endmodule


module dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module dark_weights_normed_gauss_ds_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_gauss_blur_2_update_0_write_wdata(output [31:0] dark_weights_normed_gauss_blur_2_update_0_write_wdata);

endmodule


module dark_weights_normed_gauss_blur_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_weights_normed_gauss_blur_2_update_0_write_wen, input [31:0] dark_weights_normed_gauss_blur_2_update_0_write_wdata, input [31:0] dark_weights_normed_gauss_ds_2_update_0_read_dummy, output [31:0] dark_weights_normed_gauss_ds_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_weights_normed_gauss_blur_2_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_normed_gauss_blur_2_update_0_write_wen;

  // dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1
  logic [0:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_done;
  dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1 dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1(.clk(dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_clk), .rst(dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_rst), .start(dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_start), .done(dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_done));
  assign dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_clk = clk;
  assign dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write0_merged_banks_1

  // selector_dark_weights_normed_gauss_ds_2_rd0_select
  logic [0:0] selector_dark_weights_normed_gauss_ds_2_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_ds_2_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_ds_2_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_ds_2_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_ds_2_rd0_select_out;
  dark_weights_normed_gauss_ds_2_rd0_select selector_dark_weights_normed_gauss_ds_2_rd0_select(.clk(selector_dark_weights_normed_gauss_ds_2_rd0_select_clk), .rst(selector_dark_weights_normed_gauss_ds_2_rd0_select_rst), .d0(selector_dark_weights_normed_gauss_ds_2_rd0_select_d0), .d1(selector_dark_weights_normed_gauss_ds_2_rd0_select_d1), .out(selector_dark_weights_normed_gauss_ds_2_rd0_select_out));
  assign selector_dark_weights_normed_gauss_ds_2_rd0_select_clk = clk;
  assign selector_dark_weights_normed_gauss_ds_2_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_ds_2_rd0_select

  // Bindings to dark_weights_normed_gauss_blur_2_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_normed_gauss_blur_2_update_0_write_wdata;

  // Bindings to dark_weights_normed_gauss_ds_2_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_weights_normed_gauss_ds_2_update_0_read_dummy;

  // Bindings to dark_weights_normed_gauss_ds_2_update_0_read_rdata
    // wr_3
  assign dark_weights_normed_gauss_ds_2_update_0_read_rdata = rd_2;



endmodule


module in_wire_dark_weights_normed_gauss_ds_2_update_0_read_dummy(output [31:0] dark_weights_normed_gauss_ds_2_update_0_read_dummy);

endmodule


module out_wire_dark_weights_normed_gauss_ds_2_update_0_read_rdata(input [31:0] dark_weights_normed_gauss_ds_2_update_0_read_rdata);

endmodule


module in_wire_dark_weights_normed_gauss_blur_3_update_0_write_wen(output [0:0] dark_weights_normed_gauss_blur_3_update_0_write_wen);

endmodule


module dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module dark_weights_normed_gauss_ds_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_gauss_blur_3_update_0_write_wdata(output [31:0] dark_weights_normed_gauss_blur_3_update_0_write_wdata);

endmodule


module in_wire_dark_weights_normed_gauss_ds_3_update_0_read_dummy(output [31:0] dark_weights_normed_gauss_ds_3_update_0_read_dummy);

endmodule


module out_wire_dark_weights_normed_gauss_ds_3_update_0_read_rdata(input [31:0] dark_weights_normed_gauss_ds_3_update_0_read_rdata);

endmodule


module dark_weights_normed_gauss_blur_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_weights_normed_gauss_blur_3_update_0_write_wen, input [31:0] dark_weights_normed_gauss_blur_3_update_0_write_wdata, input [31:0] dark_weights_normed_gauss_ds_3_update_0_read_dummy, output [31:0] dark_weights_normed_gauss_ds_3_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_weights_normed_gauss_blur_3_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_normed_gauss_blur_3_update_0_write_wen;

  // dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1
  logic [0:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_done;
  dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1 dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1(.clk(dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_clk), .rst(dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_rst), .start(dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_start), .done(dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_done));
  assign dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_clk = clk;
  assign dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write0_merged_banks_1

  // selector_dark_weights_normed_gauss_ds_3_rd0_select
  logic [0:0] selector_dark_weights_normed_gauss_ds_3_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_ds_3_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_ds_3_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_ds_3_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_ds_3_rd0_select_out;
  dark_weights_normed_gauss_ds_3_rd0_select selector_dark_weights_normed_gauss_ds_3_rd0_select(.clk(selector_dark_weights_normed_gauss_ds_3_rd0_select_clk), .rst(selector_dark_weights_normed_gauss_ds_3_rd0_select_rst), .d0(selector_dark_weights_normed_gauss_ds_3_rd0_select_d0), .d1(selector_dark_weights_normed_gauss_ds_3_rd0_select_d1), .out(selector_dark_weights_normed_gauss_ds_3_rd0_select_out));
  assign selector_dark_weights_normed_gauss_ds_3_rd0_select_clk = clk;
  assign selector_dark_weights_normed_gauss_ds_3_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_ds_3_rd0_select

  // Bindings to dark_weights_normed_gauss_blur_3_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_normed_gauss_blur_3_update_0_write_wdata;

  // Bindings to dark_weights_normed_gauss_ds_3_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_weights_normed_gauss_ds_3_update_0_read_dummy;

  // Bindings to dark_weights_normed_gauss_ds_3_update_0_read_rdata
    // wr_3
  assign dark_weights_normed_gauss_ds_3_update_0_read_rdata = rd_2;



endmodule


module dark_weights_normed_gauss_blur_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1264;
    end
  end

endmodule


module dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_628 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_628 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f17
  logic [0:0] f17_wen;
  logic [31:0] f17_wdata;
  logic [0:0] f17_clk;
  logic [0:0] f17_rst;
  logic [31:0] f17_rdata;
  sr_buffer_32_2527 f17(.wen(f17_wen), .wdata(f17_wdata), .clk(f17_clk), .rst(f17_rst), .rdata(f17_rdata));
  assign f17_clk = clk;
  assign f17_rst = rst;
  // Bindings to f17

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18



endmodule


module dark_weights_normed_gauss_blur_2_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 633;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_2_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1263;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_2_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_2_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 632;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_2_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_312 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_312 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0



endmodule


module dark_weights_normed_gauss_blur_3_rd1_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 317;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_3_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 632;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_3_rd2_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 2;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_3_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (311 - d0 >= 0) ? (630) : (-312 + d0 == 0) ? (630) : 0;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_3_rd3_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 631;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_3_rd4_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 316;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_3_rd5_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 1;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_3_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_final_merged_1_update_0_read_dummy(output [31:0] final_merged_1_update_0_read_dummy);

endmodule


module dark_weights_normed_gauss_blur_3_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (311 - d0 >= 0) ? (315) : (-312 + d0 == 0) ? (315) : 0;
    end
  end

endmodule


module out_wire_final_merged_1_update_0_read_rdata(input [31:0] final_merged_1_update_0_read_rdata);

endmodule


module in_wire_fused_level_0_update_0_write_wen(output [0:0] fused_level_0_update_0_write_wen);

endmodule


module final_merged_0_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_fused_level_0_update_0_write_wdata(output [31:0] fused_level_0_update_0_write_wdata);

endmodule


module in_wire_fused_level_1_update_0_write_wen(output [0:0] fused_level_1_update_0_write_wen);

endmodule


module final_merged_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_fused_level_1_update_0_write_wdata(output [31:0] fused_level_1_update_0_write_wdata);

endmodule


module in_wire_fused_level_2_update_0_write_wen(output [0:0] fused_level_2_update_0_write_wen);

endmodule


module in_wire_fused_level_2_update_0_write_wdata(output [31:0] fused_level_2_update_0_write_wdata);

endmodule


module in_wire_final_merged_2_update_0_read_dummy(output [31:0] final_merged_2_update_0_read_dummy);

endmodule


module out_wire_final_merged_2_update_0_read_rdata(input [31:0] final_merged_2_update_0_read_rdata);

endmodule


module dark_laplace_us_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module dark_weights_normed_gauss_blur_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_weights_normed_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module fused_level_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module in_wire_dark_gauss_ds_2_update_0_write_wdata(output [31:0] dark_gauss_ds_2_update_0_write_wdata);

endmodule


module dark_laplace_diff_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] dark_laplace_diff_0_update_0_write_wdata, output [31:0] fused_level_0_update_0_read_rdata, input [31:0] fused_level_0_update_0_read_dummy, input [0:0] dark_laplace_diff_0_update_0_write_wen);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1
  logic [0:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_done;
  dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1 dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1(.clk(dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_clk), .rst(dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_rst), .start(dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_start), .done(dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_done));
  assign dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_clk = clk;
  assign dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_laplace_diff_0_dark_laplace_diff_0_update_0_write0_merged_banks_1

  // selector_fused_level_0_rd0_select
  logic [0:0] selector_fused_level_0_rd0_select_clk;
  logic [0:0] selector_fused_level_0_rd0_select_rst;
  logic [31:0] selector_fused_level_0_rd0_select_d0;
  logic [31:0] selector_fused_level_0_rd0_select_d1;
  logic [31:0] selector_fused_level_0_rd0_select_out;
  fused_level_0_rd0_select selector_fused_level_0_rd0_select(.clk(selector_fused_level_0_rd0_select_clk), .rst(selector_fused_level_0_rd0_select_rst), .d0(selector_fused_level_0_rd0_select_d0), .d1(selector_fused_level_0_rd0_select_d1), .out(selector_fused_level_0_rd0_select_out));
  assign selector_fused_level_0_rd0_select_clk = clk;
  assign selector_fused_level_0_rd0_select_rst = rst;
  // Bindings to selector_fused_level_0_rd0_select

  // Bindings to dark_laplace_diff_0_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_laplace_diff_0_update_0_write_wdata;

  // Bindings to fused_level_0_update_0_read_rdata
    // wr_3
  assign fused_level_0_update_0_read_rdata = rd_2;

  // Bindings to fused_level_0_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_0_update_0_read_dummy;

  // Bindings to dark_laplace_diff_0_update_0_write_wen
    // rd_0
  assign rd_0 = dark_laplace_diff_0_update_0_write_wen;



endmodule


module in_wire_dark_gauss_blur_3_update_0_read_dummy(output [287:0] dark_gauss_blur_3_update_0_read_dummy);

endmodule


module out_wire_dark_gauss_blur_3_update_0_read_rdata(input [287:0] dark_gauss_blur_3_update_0_read_rdata);

endmodule


module in_wire_dark_laplace_diff_2_update_0_read_dummy(output [31:0] dark_laplace_diff_2_update_0_read_dummy);

endmodule


module out_wire_dark_laplace_diff_2_update_0_read_rdata(input [31:0] dark_laplace_diff_2_update_0_read_rdata);

endmodule


module in_wire_dark_laplace_us_1_update_0_read_dummy(output [31:0] dark_laplace_us_1_update_0_read_dummy);

endmodule


module out_wire_dark_laplace_us_1_update_0_read_rdata(input [31:0] dark_laplace_us_1_update_0_read_rdata);

endmodule


module dark_laplace_diff_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] dark_laplace_diff_1_update_0_write_wdata, output [31:0] fused_level_1_update_0_read_rdata, input [0:0] dark_laplace_diff_1_update_0_write_wen, input [31:0] fused_level_1_update_0_read_dummy);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_laplace_diff_1_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_laplace_diff_1_update_0_write_wdata;

  // Bindings to fused_level_1_update_0_read_rdata
    // wr_3
  assign fused_level_1_update_0_read_rdata = rd_2;

  // Bindings to dark_laplace_diff_1_update_0_write_wen
    // rd_0
  assign rd_0 = dark_laplace_diff_1_update_0_write_wen;

  // Bindings to fused_level_1_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_1_update_0_read_dummy;

  // selector_fused_level_1_rd0_select
  logic [0:0] selector_fused_level_1_rd0_select_clk;
  logic [0:0] selector_fused_level_1_rd0_select_rst;
  logic [31:0] selector_fused_level_1_rd0_select_d0;
  logic [31:0] selector_fused_level_1_rd0_select_d1;
  logic [31:0] selector_fused_level_1_rd0_select_out;
  fused_level_1_rd0_select selector_fused_level_1_rd0_select(.clk(selector_fused_level_1_rd0_select_clk), .rst(selector_fused_level_1_rd0_select_rst), .d0(selector_fused_level_1_rd0_select_d0), .d1(selector_fused_level_1_rd0_select_d1), .out(selector_fused_level_1_rd0_select_out));
  assign selector_fused_level_1_rd0_select_clk = clk;
  assign selector_fused_level_1_rd0_select_rst = rst;
  // Bindings to selector_fused_level_1_rd0_select

  // dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1
  logic [0:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_done;
  dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1 dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1(.clk(dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_clk), .rst(dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_rst), .start(dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_start), .done(dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_done));
  assign dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_clk = clk;
  assign dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1



endmodule


module dark_laplace_diff_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_laplace_diff_2_update_0_write_wen, input [31:0] fused_level_2_update_0_read_dummy, input [31:0] dark_laplace_diff_2_update_0_write_wdata, output [31:0] fused_level_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_laplace_diff_2_update_0_write_wen
    // rd_0
  assign rd_0 = dark_laplace_diff_2_update_0_write_wen;

  // Bindings to fused_level_2_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_2_update_0_read_dummy;

  // selector_fused_level_2_rd0_select
  logic [0:0] selector_fused_level_2_rd0_select_clk;
  logic [0:0] selector_fused_level_2_rd0_select_rst;
  logic [31:0] selector_fused_level_2_rd0_select_d0;
  logic [31:0] selector_fused_level_2_rd0_select_d1;
  logic [31:0] selector_fused_level_2_rd0_select_out;
  fused_level_2_rd0_select selector_fused_level_2_rd0_select(.clk(selector_fused_level_2_rd0_select_clk), .rst(selector_fused_level_2_rd0_select_rst), .d0(selector_fused_level_2_rd0_select_d0), .d1(selector_fused_level_2_rd0_select_d1), .out(selector_fused_level_2_rd0_select_out));
  assign selector_fused_level_2_rd0_select_clk = clk;
  assign selector_fused_level_2_rd0_select_rst = rst;
  // Bindings to selector_fused_level_2_rd0_select

  // Bindings to dark_laplace_diff_2_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_laplace_diff_2_update_0_write_wdata;

  // Bindings to fused_level_2_update_0_read_rdata
    // wr_3
  assign fused_level_2_update_0_read_rdata = rd_2;

  // dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1
  logic [0:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_done;
  dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1 dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1(.clk(dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_clk), .rst(dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_rst), .start(dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_start), .done(dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_done));
  assign dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_clk = clk;
  assign dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1



endmodule


module dark_laplace_diff_1_dark_laplace_diff_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module dark_laplace_us_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_laplace_us_0_update_0_write_wen, input [31:0] dark_laplace_us_0_update_0_write_wdata, input [31:0] dark_laplace_diff_0_update_0_read_dummy, output [31:0] dark_laplace_diff_0_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to dark_laplace_us_0_update_0_write_wen
    // rd_0
  assign rd_0 = dark_laplace_us_0_update_0_write_wen;

  // selector_dark_laplace_diff_0_rd0_select
  logic [0:0] selector_dark_laplace_diff_0_rd0_select_clk;
  logic [0:0] selector_dark_laplace_diff_0_rd0_select_rst;
  logic [31:0] selector_dark_laplace_diff_0_rd0_select_d0;
  logic [31:0] selector_dark_laplace_diff_0_rd0_select_d1;
  logic [31:0] selector_dark_laplace_diff_0_rd0_select_out;
  dark_laplace_diff_0_rd0_select selector_dark_laplace_diff_0_rd0_select(.clk(selector_dark_laplace_diff_0_rd0_select_clk), .rst(selector_dark_laplace_diff_0_rd0_select_rst), .d0(selector_dark_laplace_diff_0_rd0_select_d0), .d1(selector_dark_laplace_diff_0_rd0_select_d1), .out(selector_dark_laplace_diff_0_rd0_select_out));
  assign selector_dark_laplace_diff_0_rd0_select_clk = clk;
  assign selector_dark_laplace_diff_0_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_diff_0_rd0_select

  // Bindings to dark_laplace_us_0_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_laplace_us_0_update_0_write_wdata;

  // Bindings to dark_laplace_diff_0_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_laplace_diff_0_update_0_read_dummy;

  // Bindings to dark_laplace_diff_0_update_0_read_rdata
    // wr_3
  assign dark_laplace_diff_0_update_0_read_rdata = rd_2;

  // dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1
  logic [0:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_done;
  dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1 dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1(.clk(dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_clk), .rst(dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_rst), .start(dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_start), .done(dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_done));
  assign dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_clk = clk;
  assign dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1



endmodule


module dark_laplace_diff_2_dark_laplace_diff_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_laplace_us_1_update_0_write_wen(output [0:0] dark_laplace_us_1_update_0_write_wen);

endmodule


module dark_laplace_us_0_dark_laplace_us_0_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module dark_laplace_diff_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_laplace_us_1_update_0_write_wdata(output [31:0] dark_laplace_us_1_update_0_write_wdata);

endmodule


module dark_laplace_us_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] dark_laplace_diff_1_update_0_read_dummy, output [31:0] dark_laplace_diff_1_update_0_read_rdata, input [31:0] dark_laplace_us_1_update_0_write_wdata, input [0:0] dark_laplace_us_1_update_0_write_wen);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // selector_dark_laplace_diff_1_rd0_select
  logic [0:0] selector_dark_laplace_diff_1_rd0_select_clk;
  logic [0:0] selector_dark_laplace_diff_1_rd0_select_rst;
  logic [31:0] selector_dark_laplace_diff_1_rd0_select_d0;
  logic [31:0] selector_dark_laplace_diff_1_rd0_select_d1;
  logic [31:0] selector_dark_laplace_diff_1_rd0_select_out;
  dark_laplace_diff_1_rd0_select selector_dark_laplace_diff_1_rd0_select(.clk(selector_dark_laplace_diff_1_rd0_select_clk), .rst(selector_dark_laplace_diff_1_rd0_select_rst), .d0(selector_dark_laplace_diff_1_rd0_select_d0), .d1(selector_dark_laplace_diff_1_rd0_select_d1), .out(selector_dark_laplace_diff_1_rd0_select_out));
  assign selector_dark_laplace_diff_1_rd0_select_clk = clk;
  assign selector_dark_laplace_diff_1_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_diff_1_rd0_select

  // Bindings to dark_laplace_diff_1_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_laplace_diff_1_update_0_read_dummy;

  // Bindings to dark_laplace_diff_1_update_0_read_rdata
    // wr_3
  assign dark_laplace_diff_1_update_0_read_rdata = rd_2;

  // Bindings to dark_laplace_us_1_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_laplace_us_1_update_0_write_wdata;

  // Bindings to dark_laplace_us_1_update_0_write_wen
    // rd_0
  assign rd_0 = dark_laplace_us_1_update_0_write_wen;

  // dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1
  logic [0:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_done;
  dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1 dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1(.clk(dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_clk), .rst(dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_rst), .start(dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_start), .done(dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_done));
  assign dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_clk = clk;
  assign dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_laplace_us_1_dark_laplace_us_1_update_0_write0_merged_banks_1



endmodule


module in_wire_dark_laplace_us_2_update_0_write_wen(output [0:0] dark_laplace_us_2_update_0_write_wen);

endmodule


module dark_laplace_diff_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_laplace_us_2_update_0_write_wdata(output [31:0] dark_laplace_us_2_update_0_write_wdata);

endmodule


module dark_laplace_us_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] dark_laplace_diff_2_update_0_read_rdata, input [31:0] dark_laplace_diff_2_update_0_read_dummy, input [31:0] dark_laplace_us_2_update_0_write_wdata, input [0:0] dark_laplace_us_2_update_0_write_wen);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1
  logic [0:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_done;
  dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1 dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1(.clk(dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_clk), .rst(dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_rst), .start(dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_start), .done(dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_done));
  assign dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_clk = clk;
  assign dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_laplace_us_2_dark_laplace_us_2_update_0_write0_merged_banks_1

  // Bindings to dark_laplace_diff_2_update_0_read_rdata
    // wr_3
  assign dark_laplace_diff_2_update_0_read_rdata = rd_2;

  // Bindings to dark_laplace_diff_2_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_laplace_diff_2_update_0_read_dummy;

  // Bindings to dark_laplace_us_2_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_laplace_us_2_update_0_write_wdata;

  // Bindings to dark_laplace_us_2_update_0_write_wen
    // rd_0
  assign rd_0 = dark_laplace_us_2_update_0_write_wen;

  // selector_dark_laplace_diff_2_rd0_select
  logic [0:0] selector_dark_laplace_diff_2_rd0_select_clk;
  logic [0:0] selector_dark_laplace_diff_2_rd0_select_rst;
  logic [31:0] selector_dark_laplace_diff_2_rd0_select_d0;
  logic [31:0] selector_dark_laplace_diff_2_rd0_select_d1;
  logic [31:0] selector_dark_laplace_diff_2_rd0_select_out;
  dark_laplace_diff_2_rd0_select selector_dark_laplace_diff_2_rd0_select(.clk(selector_dark_laplace_diff_2_rd0_select_clk), .rst(selector_dark_laplace_diff_2_rd0_select_rst), .d0(selector_dark_laplace_diff_2_rd0_select_d0), .d1(selector_dark_laplace_diff_2_rd0_select_d1), .out(selector_dark_laplace_diff_2_rd0_select_out));
  assign selector_dark_laplace_diff_2_rd0_select_clk = clk;
  assign selector_dark_laplace_diff_2_rd0_select_rst = rst;
  // Bindings to selector_dark_laplace_diff_2_rd0_select



endmodule


module in_wire_dark_weights_update_0_write_wen(output [0:0] dark_weights_update_0_write_wen);

endmodule


module dark_weights_dark_weights_update_0_write0_merged_banks_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in_wire_dark_weights_update_0_write_wdata(output [31:0] dark_weights_update_0_write_wdata);

endmodule


module weight_sums_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_dark_weights_normed_update_0_read_dummy(output [31:0] dark_weights_normed_update_0_read_dummy);

endmodule


module out_wire_dark_weights_normed_update_0_read_rdata(input [31:0] dark_weights_normed_update_0_read_rdata);

endmodule


module dark_weights(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] dark_weights_update_0_write_wen, input [31:0] dark_weights_normed_update_0_read_dummy, input [31:0] dark_weights_update_0_write_wdata, output [31:0] weight_sums_update_0_read_rdata, input [31:0] weight_sums_update_0_read_dummy, output [31:0] dark_weights_normed_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // Bindings to dark_weights_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_update_0_write_wen;

  // Bindings to dark_weights_normed_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_weights_normed_update_0_read_dummy;

  // Bindings to dark_weights_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_update_0_write_wdata;

  // selector_dark_weights_normed_rd0_select
  logic [0:0] selector_dark_weights_normed_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_rd0_select_out;
  dark_weights_normed_rd0_select selector_dark_weights_normed_rd0_select(.clk(selector_dark_weights_normed_rd0_select_clk), .rst(selector_dark_weights_normed_rd0_select_rst), .d0(selector_dark_weights_normed_rd0_select_d0), .d1(selector_dark_weights_normed_rd0_select_d1), .out(selector_dark_weights_normed_rd0_select_out));
  assign selector_dark_weights_normed_rd0_select_clk = clk;
  assign selector_dark_weights_normed_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_rd0_select

  // selector_weight_sums_rd0_select
  logic [0:0] selector_weight_sums_rd0_select_clk;
  logic [0:0] selector_weight_sums_rd0_select_rst;
  logic [31:0] selector_weight_sums_rd0_select_d0;
  logic [31:0] selector_weight_sums_rd0_select_d1;
  logic [31:0] selector_weight_sums_rd0_select_out;
  weight_sums_rd0_select selector_weight_sums_rd0_select(.clk(selector_weight_sums_rd0_select_clk), .rst(selector_weight_sums_rd0_select_rst), .d0(selector_weight_sums_rd0_select_d0), .d1(selector_weight_sums_rd0_select_d1), .out(selector_weight_sums_rd0_select_out));
  assign selector_weight_sums_rd0_select_clk = clk;
  assign selector_weight_sums_rd0_select_rst = rst;
  // Bindings to selector_weight_sums_rd0_select

  // dark_weights_dark_weights_update_0_write0_merged_banks_2
  logic [0:0] dark_weights_dark_weights_update_0_write0_merged_banks_2_clk;
  logic [0:0] dark_weights_dark_weights_update_0_write0_merged_banks_2_rst;
  logic [0:0] dark_weights_dark_weights_update_0_write0_merged_banks_2_start;
  logic [0:0] dark_weights_dark_weights_update_0_write0_merged_banks_2_done;
  dark_weights_dark_weights_update_0_write0_merged_banks_2 dark_weights_dark_weights_update_0_write0_merged_banks_2(.clk(dark_weights_dark_weights_update_0_write0_merged_banks_2_clk), .rst(dark_weights_dark_weights_update_0_write0_merged_banks_2_rst), .start(dark_weights_dark_weights_update_0_write0_merged_banks_2_start), .done(dark_weights_dark_weights_update_0_write0_merged_banks_2_done));
  assign dark_weights_dark_weights_update_0_write0_merged_banks_2_clk = clk;
  assign dark_weights_dark_weights_update_0_write0_merged_banks_2_rst = rst;
  // Bindings to dark_weights_dark_weights_update_0_write0_merged_banks_2

  // Bindings to weight_sums_update_0_read_rdata
    // wr_5
  assign weight_sums_update_0_read_rdata = rd_4;

  // Bindings to weight_sums_update_0_read_dummy
    // rd_4
  assign rd_4 = weight_sums_update_0_read_dummy;

  // Bindings to dark_weights_normed_update_0_read_rdata
    // wr_3
  assign dark_weights_normed_update_0_read_rdata = rd_2;



endmodule


module dark_weights_normed_gauss_blur_2_rd6_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (627 - d0 >= 0) ? (1262) : (-628 + d0 == 0) ? (1262) : 0;
    end
  end

endmodule


module dark_weights_normed_gauss_blur_2_rd7_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = (627 - d0 >= 0) ? (631) : (-628 + d0 == 0) ? (631) : 0;
    end
  end

endmodule


module dark_weights_normed_dark_weights_normed_update_0_write0_merged_banks_9(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f11
  logic [0:0] f11_wen;
  logic [31:0] f11_wdata;
  logic [0:0] f11_clk;
  logic [0:0] f11_rst;
  logic [31:0] f11_rdata;
  sr_buffer_32_1260 f11(.wen(f11_wen), .wdata(f11_wdata), .clk(f11_clk), .rst(f11_rst), .rdata(f11_rdata));
  assign f11_clk = clk;
  assign f11_rst = rst;
  // Bindings to f11

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f5
  logic [0:0] f5_wen;
  logic [31:0] f5_wdata;
  logic [0:0] f5_clk;
  logic [0:0] f5_rst;
  logic [31:0] f5_rdata;
  sr_buffer_32_1260 f5(.wen(f5_wen), .wdata(f5_wdata), .clk(f5_clk), .rst(f5_rst), .rdata(f5_rdata));
  assign f5_clk = clk;
  assign f5_rst = rst;
  // Bindings to f5

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0



endmodule


module dark_weights_normed_gauss_blur_2_rd8_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module fused_level_1_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 3792;
    end
  end

endmodule


module in_wire_dark_weights_normed_gauss_ds_1_update_0_write_wen(output [0:0] dark_weights_normed_gauss_ds_1_update_0_write_wen);

endmodule


module in_wire_dark_weights_normed_gauss_ds_1_update_0_write_wdata(output [31:0] dark_weights_normed_gauss_ds_1_update_0_write_wdata);

endmodule


module in_wire_dark_weights_normed_gauss_blur_2_update_0_read_dummy(output [287:0] dark_weights_normed_gauss_blur_2_update_0_read_dummy);

endmodule


module out_wire_dark_weights_normed_gauss_blur_2_update_0_read_rdata(input [287:0] dark_weights_normed_gauss_blur_2_update_0_read_rdata);

endmodule


module dark_weights_normed_gauss_ds_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] dark_weights_normed_gauss_ds_1_update_0_write_wdata, output [31:0] fused_level_1_update_0_read_rdata, output [287:0] dark_weights_normed_gauss_blur_2_update_0_read_rdata, input [287:0] dark_weights_normed_gauss_blur_2_update_0_read_dummy, input [31:0] fused_level_1_update_0_read_dummy, input [0:0] dark_weights_normed_gauss_ds_1_update_0_write_wen);

  logic [31:0] rd_4;
  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_4_stage_1;
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_4_stage_1 <= rd_4;
      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10
  logic [0:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_clk;
  logic [0:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_rst;
  logic [0:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_start;
  logic [0:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_done;
  dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10 dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10(.clk(dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_clk), .rst(dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_rst), .start(dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_start), .done(dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_done));
  assign dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_clk = clk;
  assign dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write0_merged_banks_10

  // selector_dark_weights_normed_gauss_blur_2_rd0_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd0_select_out;
  dark_weights_normed_gauss_blur_2_rd0_select selector_dark_weights_normed_gauss_blur_2_rd0_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd0_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd0_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd0_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd0_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd0_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd0_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd0_select

  // selector_dark_weights_normed_gauss_blur_2_rd1_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd1_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd1_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd1_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd1_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd1_select_out;
  dark_weights_normed_gauss_blur_2_rd1_select selector_dark_weights_normed_gauss_blur_2_rd1_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd1_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd1_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd1_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd1_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd1_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd1_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd1_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd1_select

  // selector_dark_weights_normed_gauss_blur_2_rd2_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd2_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd2_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd2_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd2_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd2_select_out;
  dark_weights_normed_gauss_blur_2_rd2_select selector_dark_weights_normed_gauss_blur_2_rd2_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd2_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd2_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd2_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd2_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd2_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd2_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd2_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd2_select

  // selector_dark_weights_normed_gauss_blur_2_rd3_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd3_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd3_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd3_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd3_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd3_select_out;
  dark_weights_normed_gauss_blur_2_rd3_select selector_dark_weights_normed_gauss_blur_2_rd3_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd3_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd3_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd3_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd3_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd3_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd3_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd3_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd3_select

  // selector_dark_weights_normed_gauss_blur_2_rd4_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd4_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd4_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd4_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd4_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd4_select_out;
  dark_weights_normed_gauss_blur_2_rd4_select selector_dark_weights_normed_gauss_blur_2_rd4_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd4_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd4_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd4_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd4_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd4_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd4_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd4_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd4_select

  // selector_dark_weights_normed_gauss_blur_2_rd5_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd5_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd5_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd5_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd5_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd5_select_out;
  dark_weights_normed_gauss_blur_2_rd5_select selector_dark_weights_normed_gauss_blur_2_rd5_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd5_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd5_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd5_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd5_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd5_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd5_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd5_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd5_select

  // Bindings to dark_weights_normed_gauss_ds_1_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_normed_gauss_ds_1_update_0_write_wdata;

  // selector_dark_weights_normed_gauss_blur_2_rd7_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd7_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd7_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd7_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd7_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd7_select_out;
  dark_weights_normed_gauss_blur_2_rd7_select selector_dark_weights_normed_gauss_blur_2_rd7_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd7_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd7_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd7_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd7_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd7_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd7_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd7_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd7_select

  // Bindings to fused_level_1_update_0_read_rdata
    // wr_5
  assign fused_level_1_update_0_read_rdata = rd_4;

  // selector_dark_weights_normed_gauss_blur_2_rd6_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd6_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd6_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd6_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd6_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd6_select_out;
  dark_weights_normed_gauss_blur_2_rd6_select selector_dark_weights_normed_gauss_blur_2_rd6_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd6_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd6_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd6_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd6_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd6_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd6_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd6_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd6_select

  // Bindings to dark_weights_normed_gauss_blur_2_update_0_read_rdata
    // wr_3
  assign dark_weights_normed_gauss_blur_2_update_0_read_rdata = rd_2;

  // Bindings to dark_weights_normed_gauss_blur_2_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_weights_normed_gauss_blur_2_update_0_read_dummy;

  // Bindings to fused_level_1_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_1_update_0_read_dummy;

  // selector_dark_weights_normed_gauss_blur_2_rd8_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd8_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_2_rd8_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd8_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd8_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_2_rd8_select_out;
  dark_weights_normed_gauss_blur_2_rd8_select selector_dark_weights_normed_gauss_blur_2_rd8_select(.clk(selector_dark_weights_normed_gauss_blur_2_rd8_select_clk), .rst(selector_dark_weights_normed_gauss_blur_2_rd8_select_rst), .d0(selector_dark_weights_normed_gauss_blur_2_rd8_select_d0), .d1(selector_dark_weights_normed_gauss_blur_2_rd8_select_d1), .out(selector_dark_weights_normed_gauss_blur_2_rd8_select_out));
  assign selector_dark_weights_normed_gauss_blur_2_rd8_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_2_rd8_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_2_rd8_select

  // Bindings to dark_weights_normed_gauss_ds_1_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_normed_gauss_ds_1_update_0_write_wen;

  // selector_fused_level_1_rd0_select
  logic [0:0] selector_fused_level_1_rd0_select_clk;
  logic [0:0] selector_fused_level_1_rd0_select_rst;
  logic [31:0] selector_fused_level_1_rd0_select_d0;
  logic [31:0] selector_fused_level_1_rd0_select_d1;
  logic [31:0] selector_fused_level_1_rd0_select_out;
  fused_level_1_rd0_select selector_fused_level_1_rd0_select(.clk(selector_fused_level_1_rd0_select_clk), .rst(selector_fused_level_1_rd0_select_rst), .d0(selector_fused_level_1_rd0_select_d0), .d1(selector_fused_level_1_rd0_select_d1), .out(selector_fused_level_1_rd0_select_out));
  assign selector_fused_level_1_rd0_select_clk = clk;
  assign selector_fused_level_1_rd0_select_rst = rst;
  // Bindings to selector_fused_level_1_rd0_select



endmodule


module dark_weights_normed_gauss_ds_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] fused_level_2_update_0_read_rdata, output [287:0] dark_weights_normed_gauss_blur_3_update_0_read_rdata, input [287:0] dark_weights_normed_gauss_blur_3_update_0_read_dummy, input [31:0] fused_level_2_update_0_read_dummy, input [31:0] dark_weights_normed_gauss_ds_2_update_0_write_wdata, input [0:0] dark_weights_normed_gauss_ds_2_update_0_write_wen);

  logic [31:0] rd_4;
  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [287:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_4_stage_1;
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [287:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_4_stage_1 <= rd_4;
      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to fused_level_2_update_0_read_rdata
    // wr_5
  assign fused_level_2_update_0_read_rdata = rd_4;

  // Bindings to dark_weights_normed_gauss_blur_3_update_0_read_rdata
    // wr_3
  assign dark_weights_normed_gauss_blur_3_update_0_read_rdata = rd_2;

  // Bindings to dark_weights_normed_gauss_blur_3_update_0_read_dummy
    // rd_2
  assign rd_2 = dark_weights_normed_gauss_blur_3_update_0_read_dummy;

  // Bindings to fused_level_2_update_0_read_dummy
    // rd_4
  assign rd_4 = fused_level_2_update_0_read_dummy;

  // Bindings to dark_weights_normed_gauss_ds_2_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_normed_gauss_ds_2_update_0_write_wdata;

  // Bindings to dark_weights_normed_gauss_ds_2_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_normed_gauss_ds_2_update_0_write_wen;

  // selector_fused_level_2_rd0_select
  logic [0:0] selector_fused_level_2_rd0_select_clk;
  logic [0:0] selector_fused_level_2_rd0_select_rst;
  logic [31:0] selector_fused_level_2_rd0_select_d0;
  logic [31:0] selector_fused_level_2_rd0_select_d1;
  logic [31:0] selector_fused_level_2_rd0_select_out;
  fused_level_2_rd0_select selector_fused_level_2_rd0_select(.clk(selector_fused_level_2_rd0_select_clk), .rst(selector_fused_level_2_rd0_select_rst), .d0(selector_fused_level_2_rd0_select_d0), .d1(selector_fused_level_2_rd0_select_d1), .out(selector_fused_level_2_rd0_select_out));
  assign selector_fused_level_2_rd0_select_clk = clk;
  assign selector_fused_level_2_rd0_select_rst = rst;
  // Bindings to selector_fused_level_2_rd0_select

  // selector_dark_weights_normed_gauss_blur_3_rd8_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd8_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd8_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd8_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd8_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd8_select_out;
  dark_weights_normed_gauss_blur_3_rd8_select selector_dark_weights_normed_gauss_blur_3_rd8_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd8_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd8_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd8_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd8_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd8_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd8_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd8_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd8_select

  // dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10
  logic [0:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_clk;
  logic [0:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_rst;
  logic [0:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_start;
  logic [0:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_done;
  dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10 dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10(.clk(dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_clk), .rst(dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_rst), .start(dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_start), .done(dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_done));
  assign dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_clk = clk;
  assign dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10_rst = rst;
  // Bindings to dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write0_merged_banks_10

  // selector_dark_weights_normed_gauss_blur_3_rd0_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd0_select_out;
  dark_weights_normed_gauss_blur_3_rd0_select selector_dark_weights_normed_gauss_blur_3_rd0_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd0_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd0_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd0_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd0_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd0_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd0_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd0_select

  // selector_dark_weights_normed_gauss_blur_3_rd2_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd2_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd2_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd2_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd2_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd2_select_out;
  dark_weights_normed_gauss_blur_3_rd2_select selector_dark_weights_normed_gauss_blur_3_rd2_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd2_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd2_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd2_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd2_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd2_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd2_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd2_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd2_select

  // selector_dark_weights_normed_gauss_blur_3_rd1_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd1_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd1_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd1_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd1_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd1_select_out;
  dark_weights_normed_gauss_blur_3_rd1_select selector_dark_weights_normed_gauss_blur_3_rd1_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd1_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd1_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd1_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd1_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd1_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd1_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd1_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd1_select

  // selector_dark_weights_normed_gauss_blur_3_rd3_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd3_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd3_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd3_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd3_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd3_select_out;
  dark_weights_normed_gauss_blur_3_rd3_select selector_dark_weights_normed_gauss_blur_3_rd3_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd3_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd3_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd3_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd3_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd3_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd3_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd3_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd3_select

  // selector_dark_weights_normed_gauss_blur_3_rd4_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd4_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd4_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd4_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd4_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd4_select_out;
  dark_weights_normed_gauss_blur_3_rd4_select selector_dark_weights_normed_gauss_blur_3_rd4_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd4_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd4_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd4_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd4_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd4_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd4_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd4_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd4_select

  // selector_dark_weights_normed_gauss_blur_3_rd6_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd6_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd6_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd6_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd6_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd6_select_out;
  dark_weights_normed_gauss_blur_3_rd6_select selector_dark_weights_normed_gauss_blur_3_rd6_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd6_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd6_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd6_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd6_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd6_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd6_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd6_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd6_select

  // selector_dark_weights_normed_gauss_blur_3_rd5_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd5_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd5_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd5_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd5_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd5_select_out;
  dark_weights_normed_gauss_blur_3_rd5_select selector_dark_weights_normed_gauss_blur_3_rd5_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd5_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd5_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd5_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd5_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd5_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd5_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd5_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd5_select

  // selector_dark_weights_normed_gauss_blur_3_rd7_select
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd7_select_clk;
  logic [0:0] selector_dark_weights_normed_gauss_blur_3_rd7_select_rst;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd7_select_d0;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd7_select_d1;
  logic [31:0] selector_dark_weights_normed_gauss_blur_3_rd7_select_out;
  dark_weights_normed_gauss_blur_3_rd7_select selector_dark_weights_normed_gauss_blur_3_rd7_select(.clk(selector_dark_weights_normed_gauss_blur_3_rd7_select_clk), .rst(selector_dark_weights_normed_gauss_blur_3_rd7_select_rst), .d0(selector_dark_weights_normed_gauss_blur_3_rd7_select_d0), .d1(selector_dark_weights_normed_gauss_blur_3_rd7_select_d1), .out(selector_dark_weights_normed_gauss_blur_3_rd7_select_out));
  assign selector_dark_weights_normed_gauss_blur_3_rd7_select_clk = clk;
  assign selector_dark_weights_normed_gauss_blur_3_rd7_select_rst = rst;
  // Bindings to selector_dark_weights_normed_gauss_blur_3_rd7_select



endmodule


module dark_weights_normed_gauss_ds_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] dark_weights_normed_gauss_ds_3_update_0_write_wdata, input [0:0] dark_weights_normed_gauss_ds_3_update_0_write_wen, input [31:0] fused_level_3_update_0_read_dummy, output [31:0] fused_level_3_update_0_read_rdata);

  logic [31:0] rd_2;
  logic [0:0] rd_0;
  logic [31:0] rd_1;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_2_stage_1;
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_2_stage_1 <= rd_2;
      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;


    end

  end


  // Data processing units...
  // Bindings to dark_weights_normed_gauss_ds_3_update_0_write_wdata
    // rd_1
  assign rd_1 = dark_weights_normed_gauss_ds_3_update_0_write_wdata;

  // dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1
  logic [0:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_clk;
  logic [0:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_rst;
  logic [0:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_start;
  logic [0:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_done;
  dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1 dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1(.clk(dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_clk), .rst(dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_rst), .start(dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_start), .done(dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_done));
  assign dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_clk = clk;
  assign dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1_rst = rst;
  // Bindings to dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1

  // Bindings to dark_weights_normed_gauss_ds_3_update_0_write_wen
    // rd_0
  assign rd_0 = dark_weights_normed_gauss_ds_3_update_0_write_wen;

  // selector_fused_level_3_rd0_select
  logic [0:0] selector_fused_level_3_rd0_select_clk;
  logic [0:0] selector_fused_level_3_rd0_select_rst;
  logic [31:0] selector_fused_level_3_rd0_select_d0;
  logic [31:0] selector_fused_level_3_rd0_select_d1;
  logic [31:0] selector_fused_level_3_rd0_select_out;
  fused_level_3_rd0_select selector_fused_level_3_rd0_select(.clk(selector_fused_level_3_rd0_select_clk), .rst(selector_fused_level_3_rd0_select_rst), .d0(selector_fused_level_3_rd0_select_d0), .d1(selector_fused_level_3_rd0_select_d1), .out(selector_fused_level_3_rd0_select_out));
  assign selector_fused_level_3_rd0_select_clk = clk;
  assign selector_fused_level_3_rd0_select_rst = rst;
  // Bindings to selector_fused_level_3_rd0_select

  // Bindings to fused_level_3_update_0_read_dummy
    // rd_2
  assign rd_2 = fused_level_3_update_0_read_dummy;

  // Bindings to fused_level_3_update_0_read_rdata
    // wr_3
  assign fused_level_3_update_0_read_rdata = rd_2;



endmodule


module dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write0_merged_banks_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module final_merged_1(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] final_merged_0_update_0_read_dummy, input [31:0] final_merged_1_update_0_write_wdata, input [0:0] final_merged_1_update_0_write_wen, output [31:0] final_merged_0_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // Bindings to final_merged_0_update_0_read_dummy
    // rd_2
  assign rd_2 = final_merged_0_update_0_read_dummy;

  // Bindings to final_merged_1_update_0_write_wdata
    // rd_1
  assign rd_1 = final_merged_1_update_0_write_wdata;

  // selector_final_merged_0_rd0_select
  logic [0:0] selector_final_merged_0_rd0_select_clk;
  logic [0:0] selector_final_merged_0_rd0_select_rst;
  logic [31:0] selector_final_merged_0_rd0_select_d0;
  logic [31:0] selector_final_merged_0_rd0_select_d1;
  logic [31:0] selector_final_merged_0_rd0_select_out;
  final_merged_0_rd0_select selector_final_merged_0_rd0_select(.clk(selector_final_merged_0_rd0_select_clk), .rst(selector_final_merged_0_rd0_select_rst), .d0(selector_final_merged_0_rd0_select_d0), .d1(selector_final_merged_0_rd0_select_d1), .out(selector_final_merged_0_rd0_select_out));
  assign selector_final_merged_0_rd0_select_clk = clk;
  assign selector_final_merged_0_rd0_select_rst = rst;
  // Bindings to selector_final_merged_0_rd0_select

  // Bindings to final_merged_1_update_0_write_wen
    // rd_0
  assign rd_0 = final_merged_1_update_0_write_wen;

  // Bindings to final_merged_0_update_0_read_rdata
    // wr_3
  assign final_merged_0_update_0_read_rdata = rd_2;

  // final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0
  logic [0:0] final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_clk;
  logic [0:0] final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_rst;
  logic [0:0] final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_start;
  logic [0:0] final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_done;
  final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0 final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0(.clk(final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_clk), .rst(final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_rst), .start(final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_start), .done(final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_done));
  assign final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_clk = clk;
  assign final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0_rst = rst;
  // Bindings to final_merged_1_final_merged_1_update_0_write0_to_final_merged_0_rd0



endmodule


module fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f106
  logic [0:0] f106_wen;
  logic [31:0] f106_wdata;
  logic [0:0] f106_clk;
  logic [0:0] f106_rst;
  logic [31:0] f106_rdata;
  sr_buffer_32_1 f106(.wen(f106_wen), .wdata(f106_wdata), .clk(f106_clk), .rst(f106_rst), .rdata(f106_rdata));
  assign f106_clk = clk;
  assign f106_rst = rst;
  // Bindings to f106

  // f110
  logic [0:0] f110_wen;
  logic [31:0] f110_wdata;
  logic [0:0] f110_clk;
  logic [0:0] f110_rst;
  logic [31:0] f110_rdata;
  sr_buffer_32_1 f110(.wen(f110_wen), .wdata(f110_wdata), .clk(f110_clk), .rst(f110_rst), .rdata(f110_rdata));
  assign f110_clk = clk;
  assign f110_rst = rst;
  // Bindings to f110

  // f112
  logic [0:0] f112_wen;
  logic [31:0] f112_wdata;
  logic [0:0] f112_clk;
  logic [0:0] f112_rst;
  logic [31:0] f112_rdata;
  sr_buffer_32_1 f112(.wen(f112_wen), .wdata(f112_wdata), .clk(f112_clk), .rst(f112_rst), .rdata(f112_rdata));
  assign f112_clk = clk;
  assign f112_rst = rst;
  // Bindings to f112

  // f108
  logic [0:0] f108_wen;
  logic [31:0] f108_wdata;
  logic [0:0] f108_clk;
  logic [0:0] f108_rst;
  logic [31:0] f108_rdata;
  sr_buffer_32_1 f108(.wen(f108_wen), .wdata(f108_wdata), .clk(f108_clk), .rst(f108_rst), .rdata(f108_rdata));
  assign f108_clk = clk;
  assign f108_rst = rst;
  // Bindings to f108

  // f114
  logic [0:0] f114_wen;
  logic [31:0] f114_wdata;
  logic [0:0] f114_clk;
  logic [0:0] f114_rst;
  logic [31:0] f114_rdata;
  sr_buffer_32_1 f114(.wen(f114_wen), .wdata(f114_wdata), .clk(f114_clk), .rst(f114_rst), .rdata(f114_rdata));
  assign f114_clk = clk;
  assign f114_rst = rst;
  // Bindings to f114

  // f116
  logic [0:0] f116_wen;
  logic [31:0] f116_wdata;
  logic [0:0] f116_clk;
  logic [0:0] f116_rst;
  logic [31:0] f116_rdata;
  sr_buffer_32_1 f116(.wen(f116_wen), .wdata(f116_wdata), .clk(f116_clk), .rst(f116_rst), .rdata(f116_rdata));
  assign f116_clk = clk;
  assign f116_rst = rst;
  // Bindings to f116

  // f122
  logic [0:0] f122_wen;
  logic [31:0] f122_wdata;
  logic [0:0] f122_clk;
  logic [0:0] f122_rst;
  logic [31:0] f122_rdata;
  sr_buffer_32_1 f122(.wen(f122_wen), .wdata(f122_wdata), .clk(f122_clk), .rst(f122_rst), .rdata(f122_rdata));
  assign f122_clk = clk;
  assign f122_rst = rst;
  // Bindings to f122

  // f124
  logic [0:0] f124_wen;
  logic [31:0] f124_wdata;
  logic [0:0] f124_clk;
  logic [0:0] f124_rst;
  logic [31:0] f124_rdata;
  sr_buffer_32_1 f124(.wen(f124_wen), .wdata(f124_wdata), .clk(f124_clk), .rst(f124_rst), .rdata(f124_rdata));
  assign f124_clk = clk;
  assign f124_rst = rst;
  // Bindings to f124

  // f126
  logic [0:0] f126_wen;
  logic [31:0] f126_wdata;
  logic [0:0] f126_clk;
  logic [0:0] f126_rst;
  logic [31:0] f126_rdata;
  sr_buffer_32_1 f126(.wen(f126_wen), .wdata(f126_wdata), .clk(f126_clk), .rst(f126_rst), .rdata(f126_rdata));
  assign f126_clk = clk;
  assign f126_rst = rst;
  // Bindings to f126

  // f120
  logic [0:0] f120_wen;
  logic [31:0] f120_wdata;
  logic [0:0] f120_clk;
  logic [0:0] f120_rst;
  logic [31:0] f120_rdata;
  sr_buffer_32_1 f120(.wen(f120_wen), .wdata(f120_wdata), .clk(f120_clk), .rst(f120_rst), .rdata(f120_rdata));
  assign f120_clk = clk;
  assign f120_rst = rst;
  // Bindings to f120

  // f130
  logic [0:0] f130_wen;
  logic [31:0] f130_wdata;
  logic [0:0] f130_clk;
  logic [0:0] f130_rst;
  logic [31:0] f130_rdata;
  sr_buffer_32_1 f130(.wen(f130_wen), .wdata(f130_wdata), .clk(f130_clk), .rst(f130_rst), .rdata(f130_rdata));
  assign f130_clk = clk;
  assign f130_rst = rst;
  // Bindings to f130

  // f128
  logic [0:0] f128_wen;
  logic [31:0] f128_wdata;
  logic [0:0] f128_clk;
  logic [0:0] f128_rst;
  logic [31:0] f128_rdata;
  sr_buffer_32_1 f128(.wen(f128_wen), .wdata(f128_wdata), .clk(f128_clk), .rst(f128_rst), .rdata(f128_rdata));
  assign f128_clk = clk;
  assign f128_rst = rst;
  // Bindings to f128

  // f132
  logic [0:0] f132_wen;
  logic [31:0] f132_wdata;
  logic [0:0] f132_clk;
  logic [0:0] f132_rst;
  logic [31:0] f132_rdata;
  sr_buffer_32_1 f132(.wen(f132_wen), .wdata(f132_wdata), .clk(f132_clk), .rst(f132_rst), .rdata(f132_rdata));
  assign f132_clk = clk;
  assign f132_rst = rst;
  // Bindings to f132

  // f134
  logic [0:0] f134_wen;
  logic [31:0] f134_wdata;
  logic [0:0] f134_clk;
  logic [0:0] f134_rst;
  logic [31:0] f134_rdata;
  sr_buffer_32_1 f134(.wen(f134_wen), .wdata(f134_wdata), .clk(f134_clk), .rst(f134_rst), .rdata(f134_rdata));
  assign f134_clk = clk;
  assign f134_rst = rst;
  // Bindings to f134

  // f136
  logic [0:0] f136_wen;
  logic [31:0] f136_wdata;
  logic [0:0] f136_clk;
  logic [0:0] f136_rst;
  logic [31:0] f136_rdata;
  sr_buffer_32_1 f136(.wen(f136_wen), .wdata(f136_wdata), .clk(f136_clk), .rst(f136_rst), .rdata(f136_rdata));
  assign f136_clk = clk;
  assign f136_rst = rst;
  // Bindings to f136

  // f140
  logic [0:0] f140_wen;
  logic [31:0] f140_wdata;
  logic [0:0] f140_clk;
  logic [0:0] f140_rst;
  logic [31:0] f140_rdata;
  sr_buffer_32_1 f140(.wen(f140_wen), .wdata(f140_wdata), .clk(f140_clk), .rst(f140_rst), .rdata(f140_rdata));
  assign f140_clk = clk;
  assign f140_rst = rst;
  // Bindings to f140

  // f138
  logic [0:0] f138_wen;
  logic [31:0] f138_wdata;
  logic [0:0] f138_clk;
  logic [0:0] f138_rst;
  logic [31:0] f138_rdata;
  sr_buffer_32_1 f138(.wen(f138_wen), .wdata(f138_wdata), .clk(f138_clk), .rst(f138_rst), .rdata(f138_rdata));
  assign f138_clk = clk;
  assign f138_rst = rst;
  // Bindings to f138

  // f142
  logic [0:0] f142_wen;
  logic [31:0] f142_wdata;
  logic [0:0] f142_clk;
  logic [0:0] f142_rst;
  logic [31:0] f142_rdata;
  sr_buffer_32_1 f142(.wen(f142_wen), .wdata(f142_wdata), .clk(f142_clk), .rst(f142_rst), .rdata(f142_rdata));
  assign f142_clk = clk;
  assign f142_rst = rst;
  // Bindings to f142

  // f144
  logic [0:0] f144_wen;
  logic [31:0] f144_wdata;
  logic [0:0] f144_clk;
  logic [0:0] f144_rst;
  logic [31:0] f144_rdata;
  sr_buffer_32_1 f144(.wen(f144_wen), .wdata(f144_wdata), .clk(f144_clk), .rst(f144_rst), .rdata(f144_rdata));
  assign f144_clk = clk;
  assign f144_rst = rst;
  // Bindings to f144

  // f146
  logic [0:0] f146_wen;
  logic [31:0] f146_wdata;
  logic [0:0] f146_clk;
  logic [0:0] f146_rst;
  logic [31:0] f146_rdata;
  sr_buffer_32_1 f146(.wen(f146_wen), .wdata(f146_wdata), .clk(f146_clk), .rst(f146_rst), .rdata(f146_rdata));
  assign f146_clk = clk;
  assign f146_rst = rst;
  // Bindings to f146

  // f148
  logic [0:0] f148_wen;
  logic [31:0] f148_wdata;
  logic [0:0] f148_clk;
  logic [0:0] f148_rst;
  logic [31:0] f148_rdata;
  sr_buffer_32_1 f148(.wen(f148_wen), .wdata(f148_wdata), .clk(f148_clk), .rst(f148_rst), .rdata(f148_rdata));
  assign f148_clk = clk;
  assign f148_rst = rst;
  // Bindings to f148

  // f118
  logic [0:0] f118_wen;
  logic [31:0] f118_wdata;
  logic [0:0] f118_clk;
  logic [0:0] f118_rst;
  logic [31:0] f118_rdata;
  sr_buffer_32_1 f118(.wen(f118_wen), .wdata(f118_wdata), .clk(f118_clk), .rst(f118_rst), .rdata(f118_rdata));
  assign f118_clk = clk;
  assign f118_rst = rst;
  // Bindings to f118

  // f150
  logic [0:0] f150_wen;
  logic [31:0] f150_wdata;
  logic [0:0] f150_clk;
  logic [0:0] f150_rst;
  logic [31:0] f150_rdata;
  sr_buffer_32_1 f150(.wen(f150_wen), .wdata(f150_wdata), .clk(f150_clk), .rst(f150_rst), .rdata(f150_rdata));
  assign f150_clk = clk;
  assign f150_rst = rst;
  // Bindings to f150

  // f104
  logic [0:0] f104_wen;
  logic [31:0] f104_wdata;
  logic [0:0] f104_clk;
  logic [0:0] f104_rst;
  logic [31:0] f104_rdata;
  sr_buffer_32_1 f104(.wen(f104_wen), .wdata(f104_wdata), .clk(f104_clk), .rst(f104_rst), .rdata(f104_rdata));
  assign f104_clk = clk;
  assign f104_rst = rst;
  // Bindings to f104

  // f100
  logic [0:0] f100_wen;
  logic [31:0] f100_wdata;
  logic [0:0] f100_clk;
  logic [0:0] f100_rst;
  logic [31:0] f100_rdata;
  sr_buffer_32_1 f100(.wen(f100_wen), .wdata(f100_wdata), .clk(f100_clk), .rst(f100_rst), .rdata(f100_rdata));
  assign f100_clk = clk;
  assign f100_rst = rst;
  // Bindings to f100

  // f102
  logic [0:0] f102_wen;
  logic [31:0] f102_wdata;
  logic [0:0] f102_clk;
  logic [0:0] f102_rst;
  logic [31:0] f102_rdata;
  sr_buffer_32_1 f102(.wen(f102_wen), .wdata(f102_wdata), .clk(f102_clk), .rst(f102_rst), .rdata(f102_rdata));
  assign f102_clk = clk;
  assign f102_rst = rst;
  // Bindings to f102

  // f98
  logic [0:0] f98_wen;
  logic [31:0] f98_wdata;
  logic [0:0] f98_clk;
  logic [0:0] f98_rst;
  logic [31:0] f98_rdata;
  sr_buffer_32_1 f98(.wen(f98_wen), .wdata(f98_wdata), .clk(f98_clk), .rst(f98_rst), .rdata(f98_rdata));
  assign f98_clk = clk;
  assign f98_rst = rst;
  // Bindings to f98

  // f96
  logic [0:0] f96_wen;
  logic [31:0] f96_wdata;
  logic [0:0] f96_clk;
  logic [0:0] f96_rst;
  logic [31:0] f96_rdata;
  sr_buffer_32_1 f96(.wen(f96_wen), .wdata(f96_wdata), .clk(f96_clk), .rst(f96_rst), .rdata(f96_rdata));
  assign f96_clk = clk;
  assign f96_rst = rst;
  // Bindings to f96

  // f94
  logic [0:0] f94_wen;
  logic [31:0] f94_wdata;
  logic [0:0] f94_clk;
  logic [0:0] f94_rst;
  logic [31:0] f94_rdata;
  sr_buffer_32_1 f94(.wen(f94_wen), .wdata(f94_wdata), .clk(f94_clk), .rst(f94_rst), .rdata(f94_rdata));
  assign f94_clk = clk;
  assign f94_rst = rst;
  // Bindings to f94

  // f92
  logic [0:0] f92_wen;
  logic [31:0] f92_wdata;
  logic [0:0] f92_clk;
  logic [0:0] f92_rst;
  logic [31:0] f92_rdata;
  sr_buffer_32_1 f92(.wen(f92_wen), .wdata(f92_wdata), .clk(f92_clk), .rst(f92_rst), .rdata(f92_rdata));
  assign f92_clk = clk;
  assign f92_rst = rst;
  // Bindings to f92

  // f90
  logic [0:0] f90_wen;
  logic [31:0] f90_wdata;
  logic [0:0] f90_clk;
  logic [0:0] f90_rst;
  logic [31:0] f90_rdata;
  sr_buffer_32_1 f90(.wen(f90_wen), .wdata(f90_wdata), .clk(f90_clk), .rst(f90_rst), .rdata(f90_rdata));
  assign f90_clk = clk;
  assign f90_rst = rst;
  // Bindings to f90

  // f88
  logic [0:0] f88_wen;
  logic [31:0] f88_wdata;
  logic [0:0] f88_clk;
  logic [0:0] f88_rst;
  logic [31:0] f88_rdata;
  sr_buffer_32_1 f88(.wen(f88_wen), .wdata(f88_wdata), .clk(f88_clk), .rst(f88_rst), .rdata(f88_rdata));
  assign f88_clk = clk;
  assign f88_rst = rst;
  // Bindings to f88

  // f86
  logic [0:0] f86_wen;
  logic [31:0] f86_wdata;
  logic [0:0] f86_clk;
  logic [0:0] f86_rst;
  logic [31:0] f86_rdata;
  sr_buffer_32_1 f86(.wen(f86_wen), .wdata(f86_wdata), .clk(f86_clk), .rst(f86_rst), .rdata(f86_rdata));
  assign f86_clk = clk;
  assign f86_rst = rst;
  // Bindings to f86

  // f82
  logic [0:0] f82_wen;
  logic [31:0] f82_wdata;
  logic [0:0] f82_clk;
  logic [0:0] f82_rst;
  logic [31:0] f82_rdata;
  sr_buffer_32_1 f82(.wen(f82_wen), .wdata(f82_wdata), .clk(f82_clk), .rst(f82_rst), .rdata(f82_rdata));
  assign f82_clk = clk;
  assign f82_rst = rst;
  // Bindings to f82

  // f84
  logic [0:0] f84_wen;
  logic [31:0] f84_wdata;
  logic [0:0] f84_clk;
  logic [0:0] f84_rst;
  logic [31:0] f84_rdata;
  sr_buffer_32_1 f84(.wen(f84_wen), .wdata(f84_wdata), .clk(f84_clk), .rst(f84_rst), .rdata(f84_rdata));
  assign f84_clk = clk;
  assign f84_rst = rst;
  // Bindings to f84

  // f74
  logic [0:0] f74_wen;
  logic [31:0] f74_wdata;
  logic [0:0] f74_clk;
  logic [0:0] f74_rst;
  logic [31:0] f74_rdata;
  sr_buffer_32_1 f74(.wen(f74_wen), .wdata(f74_wdata), .clk(f74_clk), .rst(f74_rst), .rdata(f74_rdata));
  assign f74_clk = clk;
  assign f74_rst = rst;
  // Bindings to f74

  // f80
  logic [0:0] f80_wen;
  logic [31:0] f80_wdata;
  logic [0:0] f80_clk;
  logic [0:0] f80_rst;
  logic [31:0] f80_rdata;
  sr_buffer_32_1 f80(.wen(f80_wen), .wdata(f80_wdata), .clk(f80_clk), .rst(f80_rst), .rdata(f80_rdata));
  assign f80_clk = clk;
  assign f80_rst = rst;
  // Bindings to f80

  // f78
  logic [0:0] f78_wen;
  logic [31:0] f78_wdata;
  logic [0:0] f78_clk;
  logic [0:0] f78_rst;
  logic [31:0] f78_rdata;
  sr_buffer_32_1 f78(.wen(f78_wen), .wdata(f78_wdata), .clk(f78_clk), .rst(f78_rst), .rdata(f78_rdata));
  assign f78_clk = clk;
  assign f78_rst = rst;
  // Bindings to f78

  // f76
  logic [0:0] f76_wen;
  logic [31:0] f76_wdata;
  logic [0:0] f76_clk;
  logic [0:0] f76_rst;
  logic [31:0] f76_rdata;
  sr_buffer_32_1 f76(.wen(f76_wen), .wdata(f76_wdata), .clk(f76_clk), .rst(f76_rst), .rdata(f76_rdata));
  assign f76_clk = clk;
  assign f76_rst = rst;
  // Bindings to f76

  // f72
  logic [0:0] f72_wen;
  logic [31:0] f72_wdata;
  logic [0:0] f72_clk;
  logic [0:0] f72_rst;
  logic [31:0] f72_rdata;
  sr_buffer_32_1 f72(.wen(f72_wen), .wdata(f72_wdata), .clk(f72_clk), .rst(f72_rst), .rdata(f72_rdata));
  assign f72_clk = clk;
  assign f72_rst = rst;
  // Bindings to f72

  // f68
  logic [0:0] f68_wen;
  logic [31:0] f68_wdata;
  logic [0:0] f68_clk;
  logic [0:0] f68_rst;
  logic [31:0] f68_rdata;
  sr_buffer_32_1 f68(.wen(f68_wen), .wdata(f68_wdata), .clk(f68_clk), .rst(f68_rst), .rdata(f68_rdata));
  assign f68_clk = clk;
  assign f68_rst = rst;
  // Bindings to f68

  // f70
  logic [0:0] f70_wen;
  logic [31:0] f70_wdata;
  logic [0:0] f70_clk;
  logic [0:0] f70_rst;
  logic [31:0] f70_rdata;
  sr_buffer_32_1 f70(.wen(f70_wen), .wdata(f70_wdata), .clk(f70_clk), .rst(f70_rst), .rdata(f70_rdata));
  assign f70_clk = clk;
  assign f70_rst = rst;
  // Bindings to f70

  // f60
  logic [0:0] f60_wen;
  logic [31:0] f60_wdata;
  logic [0:0] f60_clk;
  logic [0:0] f60_rst;
  logic [31:0] f60_rdata;
  sr_buffer_32_1 f60(.wen(f60_wen), .wdata(f60_wdata), .clk(f60_clk), .rst(f60_rst), .rdata(f60_rdata));
  assign f60_clk = clk;
  assign f60_rst = rst;
  // Bindings to f60

  // f66
  logic [0:0] f66_wen;
  logic [31:0] f66_wdata;
  logic [0:0] f66_clk;
  logic [0:0] f66_rst;
  logic [31:0] f66_rdata;
  sr_buffer_32_1 f66(.wen(f66_wen), .wdata(f66_wdata), .clk(f66_clk), .rst(f66_rst), .rdata(f66_rdata));
  assign f66_clk = clk;
  assign f66_rst = rst;
  // Bindings to f66

  // f64
  logic [0:0] f64_wen;
  logic [31:0] f64_wdata;
  logic [0:0] f64_clk;
  logic [0:0] f64_rst;
  logic [31:0] f64_rdata;
  sr_buffer_32_1 f64(.wen(f64_wen), .wdata(f64_wdata), .clk(f64_clk), .rst(f64_rst), .rdata(f64_rdata));
  assign f64_clk = clk;
  assign f64_rst = rst;
  // Bindings to f64

  // f62
  logic [0:0] f62_wen;
  logic [31:0] f62_wdata;
  logic [0:0] f62_clk;
  logic [0:0] f62_rst;
  logic [31:0] f62_rdata;
  sr_buffer_32_1 f62(.wen(f62_wen), .wdata(f62_wdata), .clk(f62_clk), .rst(f62_rst), .rdata(f62_rdata));
  assign f62_clk = clk;
  assign f62_rst = rst;
  // Bindings to f62

  // f58
  logic [0:0] f58_wen;
  logic [31:0] f58_wdata;
  logic [0:0] f58_clk;
  logic [0:0] f58_rst;
  logic [31:0] f58_rdata;
  sr_buffer_32_1 f58(.wen(f58_wen), .wdata(f58_wdata), .clk(f58_clk), .rst(f58_rst), .rdata(f58_rdata));
  assign f58_clk = clk;
  assign f58_rst = rst;
  // Bindings to f58

  // f56
  logic [0:0] f56_wen;
  logic [31:0] f56_wdata;
  logic [0:0] f56_clk;
  logic [0:0] f56_rst;
  logic [31:0] f56_rdata;
  sr_buffer_32_1 f56(.wen(f56_wen), .wdata(f56_wdata), .clk(f56_clk), .rst(f56_rst), .rdata(f56_rdata));
  assign f56_clk = clk;
  assign f56_rst = rst;
  // Bindings to f56

  // f54
  logic [0:0] f54_wen;
  logic [31:0] f54_wdata;
  logic [0:0] f54_clk;
  logic [0:0] f54_rst;
  logic [31:0] f54_rdata;
  sr_buffer_32_1 f54(.wen(f54_wen), .wdata(f54_wdata), .clk(f54_clk), .rst(f54_rst), .rdata(f54_rdata));
  assign f54_clk = clk;
  assign f54_rst = rst;
  // Bindings to f54

  // f52
  logic [0:0] f52_wen;
  logic [31:0] f52_wdata;
  logic [0:0] f52_clk;
  logic [0:0] f52_rst;
  logic [31:0] f52_rdata;
  sr_buffer_32_1 f52(.wen(f52_wen), .wdata(f52_wdata), .clk(f52_clk), .rst(f52_rst), .rdata(f52_rdata));
  assign f52_clk = clk;
  assign f52_rst = rst;
  // Bindings to f52

  // f50
  logic [0:0] f50_wen;
  logic [31:0] f50_wdata;
  logic [0:0] f50_clk;
  logic [0:0] f50_rst;
  logic [31:0] f50_rdata;
  sr_buffer_32_1 f50(.wen(f50_wen), .wdata(f50_wdata), .clk(f50_clk), .rst(f50_rst), .rdata(f50_rdata));
  assign f50_clk = clk;
  assign f50_rst = rst;
  // Bindings to f50

  // f48
  logic [0:0] f48_wen;
  logic [31:0] f48_wdata;
  logic [0:0] f48_clk;
  logic [0:0] f48_rst;
  logic [31:0] f48_rdata;
  sr_buffer_32_1 f48(.wen(f48_wen), .wdata(f48_wdata), .clk(f48_clk), .rst(f48_rst), .rdata(f48_rdata));
  assign f48_clk = clk;
  assign f48_rst = rst;
  // Bindings to f48

  // f46
  logic [0:0] f46_wen;
  logic [31:0] f46_wdata;
  logic [0:0] f46_clk;
  logic [0:0] f46_rst;
  logic [31:0] f46_rdata;
  sr_buffer_32_1 f46(.wen(f46_wen), .wdata(f46_wdata), .clk(f46_clk), .rst(f46_rst), .rdata(f46_rdata));
  assign f46_clk = clk;
  assign f46_rst = rst;
  // Bindings to f46

  // f44
  logic [0:0] f44_wen;
  logic [31:0] f44_wdata;
  logic [0:0] f44_clk;
  logic [0:0] f44_rst;
  logic [31:0] f44_rdata;
  sr_buffer_32_1 f44(.wen(f44_wen), .wdata(f44_wdata), .clk(f44_clk), .rst(f44_rst), .rdata(f44_rdata));
  assign f44_clk = clk;
  assign f44_rst = rst;
  // Bindings to f44

  // f42
  logic [0:0] f42_wen;
  logic [31:0] f42_wdata;
  logic [0:0] f42_clk;
  logic [0:0] f42_rst;
  logic [31:0] f42_rdata;
  sr_buffer_32_1 f42(.wen(f42_wen), .wdata(f42_wdata), .clk(f42_clk), .rst(f42_rst), .rdata(f42_rdata));
  assign f42_clk = clk;
  assign f42_rst = rst;
  // Bindings to f42

  // f40
  logic [0:0] f40_wen;
  logic [31:0] f40_wdata;
  logic [0:0] f40_clk;
  logic [0:0] f40_rst;
  logic [31:0] f40_rdata;
  sr_buffer_32_1 f40(.wen(f40_wen), .wdata(f40_wdata), .clk(f40_clk), .rst(f40_rst), .rdata(f40_rdata));
  assign f40_clk = clk;
  assign f40_rst = rst;
  // Bindings to f40

  // f34
  logic [0:0] f34_wen;
  logic [31:0] f34_wdata;
  logic [0:0] f34_clk;
  logic [0:0] f34_rst;
  logic [31:0] f34_rdata;
  sr_buffer_32_1 f34(.wen(f34_wen), .wdata(f34_wdata), .clk(f34_clk), .rst(f34_rst), .rdata(f34_rdata));
  assign f34_clk = clk;
  assign f34_rst = rst;
  // Bindings to f34

  // f38
  logic [0:0] f38_wen;
  logic [31:0] f38_wdata;
  logic [0:0] f38_clk;
  logic [0:0] f38_rst;
  logic [31:0] f38_rdata;
  sr_buffer_32_1 f38(.wen(f38_wen), .wdata(f38_wdata), .clk(f38_clk), .rst(f38_rst), .rdata(f38_rdata));
  assign f38_clk = clk;
  assign f38_rst = rst;
  // Bindings to f38

  // f36
  logic [0:0] f36_wen;
  logic [31:0] f36_wdata;
  logic [0:0] f36_clk;
  logic [0:0] f36_rst;
  logic [31:0] f36_rdata;
  sr_buffer_32_1 f36(.wen(f36_wen), .wdata(f36_wdata), .clk(f36_clk), .rst(f36_rst), .rdata(f36_rdata));
  assign f36_clk = clk;
  assign f36_rst = rst;
  // Bindings to f36

  // f32
  logic [0:0] f32_wen;
  logic [31:0] f32_wdata;
  logic [0:0] f32_clk;
  logic [0:0] f32_rst;
  logic [31:0] f32_rdata;
  sr_buffer_32_1 f32(.wen(f32_wen), .wdata(f32_wdata), .clk(f32_clk), .rst(f32_rst), .rdata(f32_rdata));
  assign f32_clk = clk;
  assign f32_rst = rst;
  // Bindings to f32

  // f30
  logic [0:0] f30_wen;
  logic [31:0] f30_wdata;
  logic [0:0] f30_clk;
  logic [0:0] f30_rst;
  logic [31:0] f30_rdata;
  sr_buffer_32_1 f30(.wen(f30_wen), .wdata(f30_wdata), .clk(f30_clk), .rst(f30_rst), .rdata(f30_rdata));
  assign f30_clk = clk;
  assign f30_rst = rst;
  // Bindings to f30

  // f28
  logic [0:0] f28_wen;
  logic [31:0] f28_wdata;
  logic [0:0] f28_clk;
  logic [0:0] f28_rst;
  logic [31:0] f28_rdata;
  sr_buffer_32_1 f28(.wen(f28_wen), .wdata(f28_wdata), .clk(f28_clk), .rst(f28_rst), .rdata(f28_rdata));
  assign f28_clk = clk;
  assign f28_rst = rst;
  // Bindings to f28

  // f26
  logic [0:0] f26_wen;
  logic [31:0] f26_wdata;
  logic [0:0] f26_clk;
  logic [0:0] f26_rst;
  logic [31:0] f26_rdata;
  sr_buffer_32_1 f26(.wen(f26_wen), .wdata(f26_wdata), .clk(f26_clk), .rst(f26_rst), .rdata(f26_rdata));
  assign f26_clk = clk;
  assign f26_rst = rst;
  // Bindings to f26

  // f22
  logic [0:0] f22_wen;
  logic [31:0] f22_wdata;
  logic [0:0] f22_clk;
  logic [0:0] f22_rst;
  logic [31:0] f22_rdata;
  sr_buffer_32_1 f22(.wen(f22_wen), .wdata(f22_wdata), .clk(f22_clk), .rst(f22_rst), .rdata(f22_rdata));
  assign f22_clk = clk;
  assign f22_rst = rst;
  // Bindings to f22

  // f24
  logic [0:0] f24_wen;
  logic [31:0] f24_wdata;
  logic [0:0] f24_clk;
  logic [0:0] f24_rst;
  logic [31:0] f24_rdata;
  sr_buffer_32_1 f24(.wen(f24_wen), .wdata(f24_wdata), .clk(f24_clk), .rst(f24_rst), .rdata(f24_rdata));
  assign f24_clk = clk;
  assign f24_rst = rst;
  // Bindings to f24

  // f14
  logic [0:0] f14_wen;
  logic [31:0] f14_wdata;
  logic [0:0] f14_clk;
  logic [0:0] f14_rst;
  logic [31:0] f14_rdata;
  sr_buffer_32_1 f14(.wen(f14_wen), .wdata(f14_wdata), .clk(f14_clk), .rst(f14_rst), .rdata(f14_rdata));
  assign f14_clk = clk;
  assign f14_rst = rst;
  // Bindings to f14

  // f20
  logic [0:0] f20_wen;
  logic [31:0] f20_wdata;
  logic [0:0] f20_clk;
  logic [0:0] f20_rst;
  logic [31:0] f20_rdata;
  sr_buffer_32_1 f20(.wen(f20_wen), .wdata(f20_wdata), .clk(f20_clk), .rst(f20_rst), .rdata(f20_rdata));
  assign f20_clk = clk;
  assign f20_rst = rst;
  // Bindings to f20

  // f18
  logic [0:0] f18_wen;
  logic [31:0] f18_wdata;
  logic [0:0] f18_clk;
  logic [0:0] f18_rst;
  logic [31:0] f18_rdata;
  sr_buffer_32_1 f18(.wen(f18_wen), .wdata(f18_wdata), .clk(f18_clk), .rst(f18_rst), .rdata(f18_rdata));
  assign f18_clk = clk;
  assign f18_rst = rst;
  // Bindings to f18

  // f16
  logic [0:0] f16_wen;
  logic [31:0] f16_wdata;
  logic [0:0] f16_clk;
  logic [0:0] f16_rst;
  logic [31:0] f16_rdata;
  sr_buffer_32_1 f16(.wen(f16_wen), .wdata(f16_wdata), .clk(f16_clk), .rst(f16_rst), .rdata(f16_rdata));
  assign f16_clk = clk;
  assign f16_rst = rst;
  // Bindings to f16

  // f12
  logic [0:0] f12_wen;
  logic [31:0] f12_wdata;
  logic [0:0] f12_clk;
  logic [0:0] f12_rst;
  logic [31:0] f12_rdata;
  sr_buffer_32_1 f12(.wen(f12_wen), .wdata(f12_wdata), .clk(f12_clk), .rst(f12_rst), .rdata(f12_rdata));
  assign f12_clk = clk;
  assign f12_rst = rst;
  // Bindings to f12

  // f10
  logic [0:0] f10_wen;
  logic [31:0] f10_wdata;
  logic [0:0] f10_clk;
  logic [0:0] f10_rst;
  logic [31:0] f10_rdata;
  sr_buffer_32_1 f10(.wen(f10_wen), .wdata(f10_wdata), .clk(f10_clk), .rst(f10_rst), .rdata(f10_rdata));
  assign f10_clk = clk;
  assign f10_rst = rst;
  // Bindings to f10

  // f4
  logic [0:0] f4_wen;
  logic [31:0] f4_wdata;
  logic [0:0] f4_clk;
  logic [0:0] f4_rst;
  logic [31:0] f4_rdata;
  sr_buffer_32_1 f4(.wen(f4_wen), .wdata(f4_wdata), .clk(f4_clk), .rst(f4_rst), .rdata(f4_rdata));
  assign f4_clk = clk;
  assign f4_rst = rst;
  // Bindings to f4

  // f8
  logic [0:0] f8_wen;
  logic [31:0] f8_wdata;
  logic [0:0] f8_clk;
  logic [0:0] f8_rst;
  logic [31:0] f8_rdata;
  sr_buffer_32_1 f8(.wen(f8_wen), .wdata(f8_wdata), .clk(f8_clk), .rst(f8_rst), .rdata(f8_rdata));
  assign f8_clk = clk;
  assign f8_rst = rst;
  // Bindings to f8

  // f6
  logic [0:0] f6_wen;
  logic [31:0] f6_wdata;
  logic [0:0] f6_clk;
  logic [0:0] f6_rst;
  logic [31:0] f6_rdata;
  sr_buffer_32_1 f6(.wen(f6_wen), .wdata(f6_wdata), .clk(f6_clk), .rst(f6_rst), .rdata(f6_rdata));
  assign f6_clk = clk;
  assign f6_rst = rst;
  // Bindings to f6

  // f2
  logic [0:0] f2_wen;
  logic [31:0] f2_wdata;
  logic [0:0] f2_clk;
  logic [0:0] f2_rst;
  logic [31:0] f2_rdata;
  sr_buffer_32_1 f2(.wen(f2_wen), .wdata(f2_wdata), .clk(f2_clk), .rst(f2_rst), .rdata(f2_rdata));
  assign f2_clk = clk;
  assign f2_rst = rst;
  // Bindings to f2

  // f0
  logic [0:0] f0_wen;
  logic [31:0] f0_wdata;
  logic [0:0] f0_clk;
  logic [0:0] f0_rst;
  logic [31:0] f0_rdata;
  sr_buffer_32_1 f0(.wen(f0_wen), .wdata(f0_wdata), .clk(f0_clk), .rst(f0_rst), .rdata(f0_rdata));
  assign f0_clk = clk;
  assign f0_rst = rst;
  // Bindings to f0

  // f162
  logic [0:0] f162_wen;
  logic [31:0] f162_wdata;
  logic [0:0] f162_clk;
  logic [0:0] f162_rst;
  logic [31:0] f162_rdata;
  sr_buffer_32_1 f162(.wen(f162_wen), .wdata(f162_wdata), .clk(f162_clk), .rst(f162_rst), .rdata(f162_rdata));
  assign f162_clk = clk;
  assign f162_rst = rst;
  // Bindings to f162

  // f166
  logic [0:0] f166_wen;
  logic [31:0] f166_wdata;
  logic [0:0] f166_clk;
  logic [0:0] f166_rst;
  logic [31:0] f166_rdata;
  sr_buffer_32_1 f166(.wen(f166_wen), .wdata(f166_wdata), .clk(f166_clk), .rst(f166_rst), .rdata(f166_rdata));
  assign f166_clk = clk;
  assign f166_rst = rst;
  // Bindings to f166

  // f164
  logic [0:0] f164_wen;
  logic [31:0] f164_wdata;
  logic [0:0] f164_clk;
  logic [0:0] f164_rst;
  logic [31:0] f164_rdata;
  sr_buffer_32_1 f164(.wen(f164_wen), .wdata(f164_wdata), .clk(f164_clk), .rst(f164_rst), .rdata(f164_rdata));
  assign f164_clk = clk;
  assign f164_rst = rst;
  // Bindings to f164

  // f152
  logic [0:0] f152_wen;
  logic [31:0] f152_wdata;
  logic [0:0] f152_clk;
  logic [0:0] f152_rst;
  logic [31:0] f152_rdata;
  sr_buffer_32_1 f152(.wen(f152_wen), .wdata(f152_wdata), .clk(f152_clk), .rst(f152_rst), .rdata(f152_rdata));
  assign f152_clk = clk;
  assign f152_rst = rst;
  // Bindings to f152

  // f160
  logic [0:0] f160_wen;
  logic [31:0] f160_wdata;
  logic [0:0] f160_clk;
  logic [0:0] f160_rst;
  logic [31:0] f160_rdata;
  sr_buffer_32_1 f160(.wen(f160_wen), .wdata(f160_wdata), .clk(f160_clk), .rst(f160_rst), .rdata(f160_rdata));
  assign f160_clk = clk;
  assign f160_rst = rst;
  // Bindings to f160

  // f158
  logic [0:0] f158_wen;
  logic [31:0] f158_wdata;
  logic [0:0] f158_clk;
  logic [0:0] f158_rst;
  logic [31:0] f158_rdata;
  sr_buffer_32_1 f158(.wen(f158_wen), .wdata(f158_wdata), .clk(f158_clk), .rst(f158_rst), .rdata(f158_rdata));
  assign f158_clk = clk;
  assign f158_rst = rst;
  // Bindings to f158

  // f156
  logic [0:0] f156_wen;
  logic [31:0] f156_wdata;
  logic [0:0] f156_clk;
  logic [0:0] f156_rst;
  logic [31:0] f156_rdata;
  sr_buffer_32_1 f156(.wen(f156_wen), .wdata(f156_wdata), .clk(f156_clk), .rst(f156_rst), .rdata(f156_rdata));
  assign f156_clk = clk;
  assign f156_rst = rst;
  // Bindings to f156

  // f154
  logic [0:0] f154_wen;
  logic [31:0] f154_wdata;
  logic [0:0] f154_clk;
  logic [0:0] f154_rst;
  logic [31:0] f154_rdata;
  sr_buffer_32_1 f154(.wen(f154_wen), .wdata(f154_wdata), .clk(f154_clk), .rst(f154_rst), .rdata(f154_rdata));
  assign f154_clk = clk;
  assign f154_rst = rst;
  // Bindings to f154

  // f210
  logic [0:0] f210_wen;
  logic [31:0] f210_wdata;
  logic [0:0] f210_clk;
  logic [0:0] f210_rst;
  logic [31:0] f210_rdata;
  sr_buffer_32_1 f210(.wen(f210_wen), .wdata(f210_wdata), .clk(f210_clk), .rst(f210_rst), .rdata(f210_rdata));
  assign f210_clk = clk;
  assign f210_rst = rst;
  // Bindings to f210

  // f214
  logic [0:0] f214_wen;
  logic [31:0] f214_wdata;
  logic [0:0] f214_clk;
  logic [0:0] f214_rst;
  logic [31:0] f214_rdata;
  sr_buffer_32_1 f214(.wen(f214_wen), .wdata(f214_wdata), .clk(f214_clk), .rst(f214_rst), .rdata(f214_rdata));
  assign f214_clk = clk;
  assign f214_rst = rst;
  // Bindings to f214

  // f216
  logic [0:0] f216_wen;
  logic [31:0] f216_wdata;
  logic [0:0] f216_clk;
  logic [0:0] f216_rst;
  logic [31:0] f216_rdata;
  sr_buffer_32_1 f216(.wen(f216_wen), .wdata(f216_wdata), .clk(f216_clk), .rst(f216_rst), .rdata(f216_rdata));
  assign f216_clk = clk;
  assign f216_rst = rst;
  // Bindings to f216

  // f208
  logic [0:0] f208_wen;
  logic [31:0] f208_wdata;
  logic [0:0] f208_clk;
  logic [0:0] f208_rst;
  logic [31:0] f208_rdata;
  sr_buffer_32_1 f208(.wen(f208_wen), .wdata(f208_wdata), .clk(f208_clk), .rst(f208_rst), .rdata(f208_rdata));
  assign f208_clk = clk;
  assign f208_rst = rst;
  // Bindings to f208

  // f224
  logic [0:0] f224_wen;
  logic [31:0] f224_wdata;
  logic [0:0] f224_clk;
  logic [0:0] f224_rst;
  logic [31:0] f224_rdata;
  sr_buffer_32_1 f224(.wen(f224_wen), .wdata(f224_wdata), .clk(f224_clk), .rst(f224_rst), .rdata(f224_rdata));
  assign f224_clk = clk;
  assign f224_rst = rst;
  // Bindings to f224

  // f186
  logic [0:0] f186_wen;
  logic [31:0] f186_wdata;
  logic [0:0] f186_clk;
  logic [0:0] f186_rst;
  logic [31:0] f186_rdata;
  sr_buffer_32_1 f186(.wen(f186_wen), .wdata(f186_wdata), .clk(f186_clk), .rst(f186_rst), .rdata(f186_rdata));
  assign f186_clk = clk;
  assign f186_rst = rst;
  // Bindings to f186

  // f188
  logic [0:0] f188_wen;
  logic [31:0] f188_wdata;
  logic [0:0] f188_clk;
  logic [0:0] f188_rst;
  logic [31:0] f188_rdata;
  sr_buffer_32_1 f188(.wen(f188_wen), .wdata(f188_wdata), .clk(f188_clk), .rst(f188_rst), .rdata(f188_rdata));
  assign f188_clk = clk;
  assign f188_rst = rst;
  // Bindings to f188

  // f200
  logic [0:0] f200_wen;
  logic [31:0] f200_wdata;
  logic [0:0] f200_clk;
  logic [0:0] f200_rst;
  logic [31:0] f200_rdata;
  sr_buffer_32_1 f200(.wen(f200_wen), .wdata(f200_wdata), .clk(f200_clk), .rst(f200_rst), .rdata(f200_rdata));
  assign f200_clk = clk;
  assign f200_rst = rst;
  // Bindings to f200

  // f192
  logic [0:0] f192_wen;
  logic [31:0] f192_wdata;
  logic [0:0] f192_clk;
  logic [0:0] f192_rst;
  logic [31:0] f192_rdata;
  sr_buffer_32_1 f192(.wen(f192_wen), .wdata(f192_wdata), .clk(f192_clk), .rst(f192_rst), .rdata(f192_rdata));
  assign f192_clk = clk;
  assign f192_rst = rst;
  // Bindings to f192

  // f194
  logic [0:0] f194_wen;
  logic [31:0] f194_wdata;
  logic [0:0] f194_clk;
  logic [0:0] f194_rst;
  logic [31:0] f194_rdata;
  sr_buffer_32_1 f194(.wen(f194_wen), .wdata(f194_wdata), .clk(f194_clk), .rst(f194_rst), .rdata(f194_rdata));
  assign f194_clk = clk;
  assign f194_rst = rst;
  // Bindings to f194

  // f228
  logic [0:0] f228_wen;
  logic [31:0] f228_wdata;
  logic [0:0] f228_clk;
  logic [0:0] f228_rst;
  logic [31:0] f228_rdata;
  sr_buffer_32_1 f228(.wen(f228_wen), .wdata(f228_wdata), .clk(f228_clk), .rst(f228_rst), .rdata(f228_rdata));
  assign f228_clk = clk;
  assign f228_rst = rst;
  // Bindings to f228

  // f196
  logic [0:0] f196_wen;
  logic [31:0] f196_wdata;
  logic [0:0] f196_clk;
  logic [0:0] f196_rst;
  logic [31:0] f196_rdata;
  sr_buffer_32_1 f196(.wen(f196_wen), .wdata(f196_wdata), .clk(f196_clk), .rst(f196_rst), .rdata(f196_rdata));
  assign f196_clk = clk;
  assign f196_rst = rst;
  // Bindings to f196

  // f190
  logic [0:0] f190_wen;
  logic [31:0] f190_wdata;
  logic [0:0] f190_clk;
  logic [0:0] f190_rst;
  logic [31:0] f190_rdata;
  sr_buffer_32_1 f190(.wen(f190_wen), .wdata(f190_wdata), .clk(f190_clk), .rst(f190_rst), .rdata(f190_rdata));
  assign f190_clk = clk;
  assign f190_rst = rst;
  // Bindings to f190

  // f202
  logic [0:0] f202_wen;
  logic [31:0] f202_wdata;
  logic [0:0] f202_clk;
  logic [0:0] f202_rst;
  logic [31:0] f202_rdata;
  sr_buffer_32_1 f202(.wen(f202_wen), .wdata(f202_wdata), .clk(f202_clk), .rst(f202_rst), .rdata(f202_rdata));
  assign f202_clk = clk;
  assign f202_rst = rst;
  // Bindings to f202

  // f230
  logic [0:0] f230_wen;
  logic [31:0] f230_wdata;
  logic [0:0] f230_clk;
  logic [0:0] f230_rst;
  logic [31:0] f230_rdata;
  sr_buffer_32_1 f230(.wen(f230_wen), .wdata(f230_wdata), .clk(f230_clk), .rst(f230_rst), .rdata(f230_rdata));
  assign f230_clk = clk;
  assign f230_rst = rst;
  // Bindings to f230

  // f218
  logic [0:0] f218_wen;
  logic [31:0] f218_wdata;
  logic [0:0] f218_clk;
  logic [0:0] f218_rst;
  logic [31:0] f218_rdata;
  sr_buffer_32_1 f218(.wen(f218_wen), .wdata(f218_wdata), .clk(f218_clk), .rst(f218_rst), .rdata(f218_rdata));
  assign f218_clk = clk;
  assign f218_rst = rst;
  // Bindings to f218

  // f178
  logic [0:0] f178_wen;
  logic [31:0] f178_wdata;
  logic [0:0] f178_clk;
  logic [0:0] f178_rst;
  logic [31:0] f178_rdata;
  sr_buffer_32_1 f178(.wen(f178_wen), .wdata(f178_wdata), .clk(f178_clk), .rst(f178_rst), .rdata(f178_rdata));
  assign f178_clk = clk;
  assign f178_rst = rst;
  // Bindings to f178

  // f234
  logic [0:0] f234_wen;
  logic [31:0] f234_wdata;
  logic [0:0] f234_clk;
  logic [0:0] f234_rst;
  logic [31:0] f234_rdata;
  sr_buffer_32_1 f234(.wen(f234_wen), .wdata(f234_wdata), .clk(f234_clk), .rst(f234_rst), .rdata(f234_rdata));
  assign f234_clk = clk;
  assign f234_rst = rst;
  // Bindings to f234

  // f220
  logic [0:0] f220_wen;
  logic [31:0] f220_wdata;
  logic [0:0] f220_clk;
  logic [0:0] f220_rst;
  logic [31:0] f220_rdata;
  sr_buffer_32_1 f220(.wen(f220_wen), .wdata(f220_wdata), .clk(f220_clk), .rst(f220_rst), .rdata(f220_rdata));
  assign f220_clk = clk;
  assign f220_rst = rst;
  // Bindings to f220

  // f222
  logic [0:0] f222_wen;
  logic [31:0] f222_wdata;
  logic [0:0] f222_clk;
  logic [0:0] f222_rst;
  logic [31:0] f222_rdata;
  sr_buffer_32_1 f222(.wen(f222_wen), .wdata(f222_wdata), .clk(f222_clk), .rst(f222_rst), .rdata(f222_rdata));
  assign f222_clk = clk;
  assign f222_rst = rst;
  // Bindings to f222

  // f212
  logic [0:0] f212_wen;
  logic [31:0] f212_wdata;
  logic [0:0] f212_clk;
  logic [0:0] f212_rst;
  logic [31:0] f212_rdata;
  sr_buffer_32_1 f212(.wen(f212_wen), .wdata(f212_wdata), .clk(f212_clk), .rst(f212_rst), .rdata(f212_rdata));
  assign f212_clk = clk;
  assign f212_rst = rst;
  // Bindings to f212

  // f226
  logic [0:0] f226_wen;
  logic [31:0] f226_wdata;
  logic [0:0] f226_clk;
  logic [0:0] f226_rst;
  logic [31:0] f226_rdata;
  sr_buffer_32_1 f226(.wen(f226_wen), .wdata(f226_wdata), .clk(f226_clk), .rst(f226_rst), .rdata(f226_rdata));
  assign f226_clk = clk;
  assign f226_rst = rst;
  // Bindings to f226

  // f198
  logic [0:0] f198_wen;
  logic [31:0] f198_wdata;
  logic [0:0] f198_clk;
  logic [0:0] f198_rst;
  logic [31:0] f198_rdata;
  sr_buffer_32_1 f198(.wen(f198_wen), .wdata(f198_wdata), .clk(f198_clk), .rst(f198_rst), .rdata(f198_rdata));
  assign f198_clk = clk;
  assign f198_rst = rst;
  // Bindings to f198

  // f232
  logic [0:0] f232_wen;
  logic [31:0] f232_wdata;
  logic [0:0] f232_clk;
  logic [0:0] f232_rst;
  logic [31:0] f232_rdata;
  sr_buffer_32_1 f232(.wen(f232_wen), .wdata(f232_wdata), .clk(f232_clk), .rst(f232_rst), .rdata(f232_rdata));
  assign f232_clk = clk;
  assign f232_rst = rst;
  // Bindings to f232

  // f206
  logic [0:0] f206_wen;
  logic [31:0] f206_wdata;
  logic [0:0] f206_clk;
  logic [0:0] f206_rst;
  logic [31:0] f206_rdata;
  sr_buffer_32_1 f206(.wen(f206_wen), .wdata(f206_wdata), .clk(f206_clk), .rst(f206_rst), .rdata(f206_rdata));
  assign f206_clk = clk;
  assign f206_rst = rst;
  // Bindings to f206

  // f204
  logic [0:0] f204_wen;
  logic [31:0] f204_wdata;
  logic [0:0] f204_clk;
  logic [0:0] f204_rst;
  logic [31:0] f204_rdata;
  sr_buffer_32_1 f204(.wen(f204_wen), .wdata(f204_wdata), .clk(f204_clk), .rst(f204_rst), .rdata(f204_rdata));
  assign f204_clk = clk;
  assign f204_rst = rst;
  // Bindings to f204

  // f170
  logic [0:0] f170_wen;
  logic [31:0] f170_wdata;
  logic [0:0] f170_clk;
  logic [0:0] f170_rst;
  logic [31:0] f170_rdata;
  sr_buffer_32_1 f170(.wen(f170_wen), .wdata(f170_wdata), .clk(f170_clk), .rst(f170_rst), .rdata(f170_rdata));
  assign f170_clk = clk;
  assign f170_rst = rst;
  // Bindings to f170

  // f174
  logic [0:0] f174_wen;
  logic [31:0] f174_wdata;
  logic [0:0] f174_clk;
  logic [0:0] f174_rst;
  logic [31:0] f174_rdata;
  sr_buffer_32_1 f174(.wen(f174_wen), .wdata(f174_wdata), .clk(f174_clk), .rst(f174_rst), .rdata(f174_rdata));
  assign f174_clk = clk;
  assign f174_rst = rst;
  // Bindings to f174

  // f172
  logic [0:0] f172_wen;
  logic [31:0] f172_wdata;
  logic [0:0] f172_clk;
  logic [0:0] f172_rst;
  logic [31:0] f172_rdata;
  sr_buffer_32_1 f172(.wen(f172_wen), .wdata(f172_wdata), .clk(f172_clk), .rst(f172_rst), .rdata(f172_rdata));
  assign f172_clk = clk;
  assign f172_rst = rst;
  // Bindings to f172

  // f168
  logic [0:0] f168_wen;
  logic [31:0] f168_wdata;
  logic [0:0] f168_clk;
  logic [0:0] f168_rst;
  logic [31:0] f168_rdata;
  sr_buffer_32_1 f168(.wen(f168_wen), .wdata(f168_wdata), .clk(f168_clk), .rst(f168_rst), .rdata(f168_rdata));
  assign f168_clk = clk;
  assign f168_rst = rst;
  // Bindings to f168

  // f176
  logic [0:0] f176_wen;
  logic [31:0] f176_wdata;
  logic [0:0] f176_clk;
  logic [0:0] f176_rst;
  logic [31:0] f176_rdata;
  sr_buffer_32_1 f176(.wen(f176_wen), .wdata(f176_wdata), .clk(f176_clk), .rst(f176_rst), .rdata(f176_rdata));
  assign f176_clk = clk;
  assign f176_rst = rst;
  // Bindings to f176

  // f182
  logic [0:0] f182_wen;
  logic [31:0] f182_wdata;
  logic [0:0] f182_clk;
  logic [0:0] f182_rst;
  logic [31:0] f182_rdata;
  sr_buffer_32_1 f182(.wen(f182_wen), .wdata(f182_wdata), .clk(f182_clk), .rst(f182_rst), .rdata(f182_rdata));
  assign f182_clk = clk;
  assign f182_rst = rst;
  // Bindings to f182

  // f180
  logic [0:0] f180_wen;
  logic [31:0] f180_wdata;
  logic [0:0] f180_clk;
  logic [0:0] f180_rst;
  logic [31:0] f180_rdata;
  sr_buffer_32_1 f180(.wen(f180_wen), .wdata(f180_wdata), .clk(f180_clk), .rst(f180_rst), .rdata(f180_rdata));
  assign f180_clk = clk;
  assign f180_rst = rst;
  // Bindings to f180

  // f184
  logic [0:0] f184_wen;
  logic [31:0] f184_wdata;
  logic [0:0] f184_clk;
  logic [0:0] f184_rst;
  logic [31:0] f184_rdata;
  sr_buffer_32_1 f184(.wen(f184_wen), .wdata(f184_wdata), .clk(f184_clk), .rst(f184_rst), .rdata(f184_rdata));
  assign f184_clk = clk;
  assign f184_rst = rst;
  // Bindings to f184

  // f236
  logic [0:0] f236_wen;
  logic [31:0] f236_wdata;
  logic [0:0] f236_clk;
  logic [0:0] f236_rst;
  logic [31:0] f236_rdata;
  sr_buffer_32_1 f236(.wen(f236_wen), .wdata(f236_wdata), .clk(f236_clk), .rst(f236_rst), .rdata(f236_rdata));
  assign f236_clk = clk;
  assign f236_rst = rst;
  // Bindings to f236

  // f238
  logic [0:0] f238_wen;
  logic [31:0] f238_wdata;
  logic [0:0] f238_clk;
  logic [0:0] f238_rst;
  logic [31:0] f238_rdata;
  sr_buffer_32_1 f238(.wen(f238_wen), .wdata(f238_wdata), .clk(f238_clk), .rst(f238_rst), .rdata(f238_rdata));
  assign f238_clk = clk;
  assign f238_rst = rst;
  // Bindings to f238

  // f240
  logic [0:0] f240_wen;
  logic [31:0] f240_wdata;
  logic [0:0] f240_clk;
  logic [0:0] f240_rst;
  logic [31:0] f240_rdata;
  sr_buffer_32_1 f240(.wen(f240_wen), .wdata(f240_wdata), .clk(f240_clk), .rst(f240_rst), .rdata(f240_rdata));
  assign f240_clk = clk;
  assign f240_rst = rst;
  // Bindings to f240

  // f242
  logic [0:0] f242_wen;
  logic [31:0] f242_wdata;
  logic [0:0] f242_clk;
  logic [0:0] f242_rst;
  logic [31:0] f242_rdata;
  sr_buffer_32_1 f242(.wen(f242_wen), .wdata(f242_wdata), .clk(f242_clk), .rst(f242_rst), .rdata(f242_rdata));
  assign f242_clk = clk;
  assign f242_rst = rst;
  // Bindings to f242

  // f244
  logic [0:0] f244_wen;
  logic [31:0] f244_wdata;
  logic [0:0] f244_clk;
  logic [0:0] f244_rst;
  logic [31:0] f244_rdata;
  sr_buffer_32_1 f244(.wen(f244_wen), .wdata(f244_wdata), .clk(f244_clk), .rst(f244_rst), .rdata(f244_rdata));
  assign f244_clk = clk;
  assign f244_rst = rst;
  // Bindings to f244

  // f246
  logic [0:0] f246_wen;
  logic [31:0] f246_wdata;
  logic [0:0] f246_clk;
  logic [0:0] f246_rst;
  logic [31:0] f246_rdata;
  sr_buffer_32_1 f246(.wen(f246_wen), .wdata(f246_wdata), .clk(f246_clk), .rst(f246_rst), .rdata(f246_rdata));
  assign f246_clk = clk;
  assign f246_rst = rst;
  // Bindings to f246

  // f248
  logic [0:0] f248_wen;
  logic [31:0] f248_wdata;
  logic [0:0] f248_clk;
  logic [0:0] f248_rst;
  logic [31:0] f248_rdata;
  sr_buffer_32_1 f248(.wen(f248_wen), .wdata(f248_wdata), .clk(f248_clk), .rst(f248_rst), .rdata(f248_rdata));
  assign f248_clk = clk;
  assign f248_rst = rst;
  // Bindings to f248

  // f250
  logic [0:0] f250_wen;
  logic [31:0] f250_wdata;
  logic [0:0] f250_clk;
  logic [0:0] f250_rst;
  logic [31:0] f250_rdata;
  sr_buffer_32_1 f250(.wen(f250_wen), .wdata(f250_wdata), .clk(f250_clk), .rst(f250_rst), .rdata(f250_rdata));
  assign f250_clk = clk;
  assign f250_rst = rst;
  // Bindings to f250

  // f252
  logic [0:0] f252_wen;
  logic [31:0] f252_wdata;
  logic [0:0] f252_clk;
  logic [0:0] f252_rst;
  logic [31:0] f252_rdata;
  sr_buffer_32_1 f252(.wen(f252_wen), .wdata(f252_wdata), .clk(f252_clk), .rst(f252_rst), .rdata(f252_rdata));
  assign f252_clk = clk;
  assign f252_rst = rst;
  // Bindings to f252

  // f254
  logic [0:0] f254_wen;
  logic [31:0] f254_wdata;
  logic [0:0] f254_clk;
  logic [0:0] f254_rst;
  logic [31:0] f254_rdata;
  sr_buffer_32_1 f254(.wen(f254_wen), .wdata(f254_wdata), .clk(f254_clk), .rst(f254_rst), .rdata(f254_rdata));
  assign f254_clk = clk;
  assign f254_rst = rst;
  // Bindings to f254

  // f256
  logic [0:0] f256_wen;
  logic [31:0] f256_wdata;
  logic [0:0] f256_clk;
  logic [0:0] f256_rst;
  logic [31:0] f256_rdata;
  sr_buffer_32_1 f256(.wen(f256_wen), .wdata(f256_wdata), .clk(f256_clk), .rst(f256_rst), .rdata(f256_rdata));
  assign f256_clk = clk;
  assign f256_rst = rst;
  // Bindings to f256

  // f258
  logic [0:0] f258_wen;
  logic [31:0] f258_wdata;
  logic [0:0] f258_clk;
  logic [0:0] f258_rst;
  logic [31:0] f258_rdata;
  sr_buffer_32_1 f258(.wen(f258_wen), .wdata(f258_wdata), .clk(f258_clk), .rst(f258_rst), .rdata(f258_rdata));
  assign f258_clk = clk;
  assign f258_rst = rst;
  // Bindings to f258

  // f260
  logic [0:0] f260_wen;
  logic [31:0] f260_wdata;
  logic [0:0] f260_clk;
  logic [0:0] f260_rst;
  logic [31:0] f260_rdata;
  sr_buffer_32_1 f260(.wen(f260_wen), .wdata(f260_wdata), .clk(f260_clk), .rst(f260_rst), .rdata(f260_rdata));
  assign f260_clk = clk;
  assign f260_rst = rst;
  // Bindings to f260

  // f262
  logic [0:0] f262_wen;
  logic [31:0] f262_wdata;
  logic [0:0] f262_clk;
  logic [0:0] f262_rst;
  logic [31:0] f262_rdata;
  sr_buffer_32_1 f262(.wen(f262_wen), .wdata(f262_wdata), .clk(f262_clk), .rst(f262_rst), .rdata(f262_rdata));
  assign f262_clk = clk;
  assign f262_rst = rst;
  // Bindings to f262

  // f264
  logic [0:0] f264_wen;
  logic [31:0] f264_wdata;
  logic [0:0] f264_clk;
  logic [0:0] f264_rst;
  logic [31:0] f264_rdata;
  sr_buffer_32_1 f264(.wen(f264_wen), .wdata(f264_wdata), .clk(f264_clk), .rst(f264_rst), .rdata(f264_rdata));
  assign f264_clk = clk;
  assign f264_rst = rst;
  // Bindings to f264

  // f266
  logic [0:0] f266_wen;
  logic [31:0] f266_wdata;
  logic [0:0] f266_clk;
  logic [0:0] f266_rst;
  logic [31:0] f266_rdata;
  sr_buffer_32_1 f266(.wen(f266_wen), .wdata(f266_wdata), .clk(f266_clk), .rst(f266_rst), .rdata(f266_rdata));
  assign f266_clk = clk;
  assign f266_rst = rst;
  // Bindings to f266

  // f268
  logic [0:0] f268_wen;
  logic [31:0] f268_wdata;
  logic [0:0] f268_clk;
  logic [0:0] f268_rst;
  logic [31:0] f268_rdata;
  sr_buffer_32_1 f268(.wen(f268_wen), .wdata(f268_wdata), .clk(f268_clk), .rst(f268_rst), .rdata(f268_rdata));
  assign f268_clk = clk;
  assign f268_rst = rst;
  // Bindings to f268

  // f270
  logic [0:0] f270_wen;
  logic [31:0] f270_wdata;
  logic [0:0] f270_clk;
  logic [0:0] f270_rst;
  logic [31:0] f270_rdata;
  sr_buffer_32_1 f270(.wen(f270_wen), .wdata(f270_wdata), .clk(f270_clk), .rst(f270_rst), .rdata(f270_rdata));
  assign f270_clk = clk;
  assign f270_rst = rst;
  // Bindings to f270

  // f272
  logic [0:0] f272_wen;
  logic [31:0] f272_wdata;
  logic [0:0] f272_clk;
  logic [0:0] f272_rst;
  logic [31:0] f272_rdata;
  sr_buffer_32_1 f272(.wen(f272_wen), .wdata(f272_wdata), .clk(f272_clk), .rst(f272_rst), .rdata(f272_rdata));
  assign f272_clk = clk;
  assign f272_rst = rst;
  // Bindings to f272

  // f274
  logic [0:0] f274_wen;
  logic [31:0] f274_wdata;
  logic [0:0] f274_clk;
  logic [0:0] f274_rst;
  logic [31:0] f274_rdata;
  sr_buffer_32_1 f274(.wen(f274_wen), .wdata(f274_wdata), .clk(f274_clk), .rst(f274_rst), .rdata(f274_rdata));
  assign f274_clk = clk;
  assign f274_rst = rst;
  // Bindings to f274

  // f276
  logic [0:0] f276_wen;
  logic [31:0] f276_wdata;
  logic [0:0] f276_clk;
  logic [0:0] f276_rst;
  logic [31:0] f276_rdata;
  sr_buffer_32_1 f276(.wen(f276_wen), .wdata(f276_wdata), .clk(f276_clk), .rst(f276_rst), .rdata(f276_rdata));
  assign f276_clk = clk;
  assign f276_rst = rst;
  // Bindings to f276

  // f278
  logic [0:0] f278_wen;
  logic [31:0] f278_wdata;
  logic [0:0] f278_clk;
  logic [0:0] f278_rst;
  logic [31:0] f278_rdata;
  sr_buffer_32_1 f278(.wen(f278_wen), .wdata(f278_wdata), .clk(f278_clk), .rst(f278_rst), .rdata(f278_rdata));
  assign f278_clk = clk;
  assign f278_rst = rst;
  // Bindings to f278

  // f280
  logic [0:0] f280_wen;
  logic [31:0] f280_wdata;
  logic [0:0] f280_clk;
  logic [0:0] f280_rst;
  logic [31:0] f280_rdata;
  sr_buffer_32_1 f280(.wen(f280_wen), .wdata(f280_wdata), .clk(f280_clk), .rst(f280_rst), .rdata(f280_rdata));
  assign f280_clk = clk;
  assign f280_rst = rst;
  // Bindings to f280

  // f282
  logic [0:0] f282_wen;
  logic [31:0] f282_wdata;
  logic [0:0] f282_clk;
  logic [0:0] f282_rst;
  logic [31:0] f282_rdata;
  sr_buffer_32_1 f282(.wen(f282_wen), .wdata(f282_wdata), .clk(f282_clk), .rst(f282_rst), .rdata(f282_rdata));
  assign f282_clk = clk;
  assign f282_rst = rst;
  // Bindings to f282

  // f284
  logic [0:0] f284_wen;
  logic [31:0] f284_wdata;
  logic [0:0] f284_clk;
  logic [0:0] f284_rst;
  logic [31:0] f284_rdata;
  sr_buffer_32_1 f284(.wen(f284_wen), .wdata(f284_wdata), .clk(f284_clk), .rst(f284_rst), .rdata(f284_rdata));
  assign f284_clk = clk;
  assign f284_rst = rst;
  // Bindings to f284

  // f286
  logic [0:0] f286_wen;
  logic [31:0] f286_wdata;
  logic [0:0] f286_clk;
  logic [0:0] f286_rst;
  logic [31:0] f286_rdata;
  sr_buffer_32_1 f286(.wen(f286_wen), .wdata(f286_wdata), .clk(f286_clk), .rst(f286_rst), .rdata(f286_rdata));
  assign f286_clk = clk;
  assign f286_rst = rst;
  // Bindings to f286

  // f288
  logic [0:0] f288_wen;
  logic [31:0] f288_wdata;
  logic [0:0] f288_clk;
  logic [0:0] f288_rst;
  logic [31:0] f288_rdata;
  sr_buffer_32_1 f288(.wen(f288_wen), .wdata(f288_wdata), .clk(f288_clk), .rst(f288_rst), .rdata(f288_rdata));
  assign f288_clk = clk;
  assign f288_rst = rst;
  // Bindings to f288

  // f290
  logic [0:0] f290_wen;
  logic [31:0] f290_wdata;
  logic [0:0] f290_clk;
  logic [0:0] f290_rst;
  logic [31:0] f290_rdata;
  sr_buffer_32_1 f290(.wen(f290_wen), .wdata(f290_wdata), .clk(f290_clk), .rst(f290_rst), .rdata(f290_rdata));
  assign f290_clk = clk;
  assign f290_rst = rst;
  // Bindings to f290

  // f292
  logic [0:0] f292_wen;
  logic [31:0] f292_wdata;
  logic [0:0] f292_clk;
  logic [0:0] f292_rst;
  logic [31:0] f292_rdata;
  sr_buffer_32_1 f292(.wen(f292_wen), .wdata(f292_wdata), .clk(f292_clk), .rst(f292_rst), .rdata(f292_rdata));
  assign f292_clk = clk;
  assign f292_rst = rst;
  // Bindings to f292

  // f294
  logic [0:0] f294_wen;
  logic [31:0] f294_wdata;
  logic [0:0] f294_clk;
  logic [0:0] f294_rst;
  logic [31:0] f294_rdata;
  sr_buffer_32_1 f294(.wen(f294_wen), .wdata(f294_wdata), .clk(f294_clk), .rst(f294_rst), .rdata(f294_rdata));
  assign f294_clk = clk;
  assign f294_rst = rst;
  // Bindings to f294

  // f296
  logic [0:0] f296_wen;
  logic [31:0] f296_wdata;
  logic [0:0] f296_clk;
  logic [0:0] f296_rst;
  logic [31:0] f296_rdata;
  sr_buffer_32_1 f296(.wen(f296_wen), .wdata(f296_wdata), .clk(f296_clk), .rst(f296_rst), .rdata(f296_rdata));
  assign f296_clk = clk;
  assign f296_rst = rst;
  // Bindings to f296

  // f298
  logic [0:0] f298_wen;
  logic [31:0] f298_wdata;
  logic [0:0] f298_clk;
  logic [0:0] f298_rst;
  logic [31:0] f298_rdata;
  sr_buffer_32_1 f298(.wen(f298_wen), .wdata(f298_wdata), .clk(f298_clk), .rst(f298_rst), .rdata(f298_rdata));
  assign f298_clk = clk;
  assign f298_rst = rst;
  // Bindings to f298

  // f300
  logic [0:0] f300_wen;
  logic [31:0] f300_wdata;
  logic [0:0] f300_clk;
  logic [0:0] f300_rst;
  logic [31:0] f300_rdata;
  sr_buffer_32_1 f300(.wen(f300_wen), .wdata(f300_wdata), .clk(f300_clk), .rst(f300_rst), .rdata(f300_rdata));
  assign f300_clk = clk;
  assign f300_rst = rst;
  // Bindings to f300

  // f302
  logic [0:0] f302_wen;
  logic [31:0] f302_wdata;
  logic [0:0] f302_clk;
  logic [0:0] f302_rst;
  logic [31:0] f302_rdata;
  sr_buffer_32_1 f302(.wen(f302_wen), .wdata(f302_wdata), .clk(f302_clk), .rst(f302_rst), .rdata(f302_rdata));
  assign f302_clk = clk;
  assign f302_rst = rst;
  // Bindings to f302

  // f304
  logic [0:0] f304_wen;
  logic [31:0] f304_wdata;
  logic [0:0] f304_clk;
  logic [0:0] f304_rst;
  logic [31:0] f304_rdata;
  sr_buffer_32_1 f304(.wen(f304_wen), .wdata(f304_wdata), .clk(f304_clk), .rst(f304_rst), .rdata(f304_rdata));
  assign f304_clk = clk;
  assign f304_rst = rst;
  // Bindings to f304

  // f306
  logic [0:0] f306_wen;
  logic [31:0] f306_wdata;
  logic [0:0] f306_clk;
  logic [0:0] f306_rst;
  logic [31:0] f306_rdata;
  sr_buffer_32_1 f306(.wen(f306_wen), .wdata(f306_wdata), .clk(f306_clk), .rst(f306_rst), .rdata(f306_rdata));
  assign f306_clk = clk;
  assign f306_rst = rst;
  // Bindings to f306

  // f308
  logic [0:0] f308_wen;
  logic [31:0] f308_wdata;
  logic [0:0] f308_clk;
  logic [0:0] f308_rst;
  logic [31:0] f308_rdata;
  sr_buffer_32_1 f308(.wen(f308_wen), .wdata(f308_wdata), .clk(f308_clk), .rst(f308_rst), .rdata(f308_rdata));
  assign f308_clk = clk;
  assign f308_rst = rst;
  // Bindings to f308

  // f310
  logic [0:0] f310_wen;
  logic [31:0] f310_wdata;
  logic [0:0] f310_clk;
  logic [0:0] f310_rst;
  logic [31:0] f310_rdata;
  sr_buffer_32_1 f310(.wen(f310_wen), .wdata(f310_wdata), .clk(f310_clk), .rst(f310_rst), .rdata(f310_rdata));
  assign f310_clk = clk;
  assign f310_rst = rst;
  // Bindings to f310

  // f312
  logic [0:0] f312_wen;
  logic [31:0] f312_wdata;
  logic [0:0] f312_clk;
  logic [0:0] f312_rst;
  logic [31:0] f312_rdata;
  sr_buffer_32_1 f312(.wen(f312_wen), .wdata(f312_wdata), .clk(f312_clk), .rst(f312_rst), .rdata(f312_rdata));
  assign f312_clk = clk;
  assign f312_rst = rst;
  // Bindings to f312



endmodule


module in_wire_fused_level_3_update_0_write_wen(output [0:0] fused_level_3_update_0_write_wen);

endmodule


module final_merged_2_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = ((-1 - d1) % 2 == 0 && 311 - d0 >= 0) ? ((156 - floord(2*d0, 4))) : 0;
    end
  end

endmodule


module in_wire_fused_level_3_update_0_write_wdata(output [31:0] fused_level_3_update_0_write_wdata);

endmodule


module fused_level_3(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] fused_level_3_update_0_write_wdata, input [0:0] fused_level_3_update_0_write_wen, input [31:0] final_merged_2_update_0_read_dummy, output [31:0] final_merged_2_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;


    end

  end


  // Data processing units...
  // selector_final_merged_2_rd0_select
  logic [0:0] selector_final_merged_2_rd0_select_clk;
  logic [0:0] selector_final_merged_2_rd0_select_rst;
  logic [31:0] selector_final_merged_2_rd0_select_d0;
  logic [31:0] selector_final_merged_2_rd0_select_d1;
  logic [31:0] selector_final_merged_2_rd0_select_out;
  final_merged_2_rd0_select selector_final_merged_2_rd0_select(.clk(selector_final_merged_2_rd0_select_clk), .rst(selector_final_merged_2_rd0_select_rst), .d0(selector_final_merged_2_rd0_select_d0), .d1(selector_final_merged_2_rd0_select_d1), .out(selector_final_merged_2_rd0_select_out));
  assign selector_final_merged_2_rd0_select_clk = clk;
  assign selector_final_merged_2_rd0_select_rst = rst;
  // Bindings to selector_final_merged_2_rd0_select

  // fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0
  logic [0:0] fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_clk;
  logic [0:0] fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_rst;
  logic [0:0] fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_start;
  logic [0:0] fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_done;
  fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0 fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0(.clk(fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_clk), .rst(fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_rst), .start(fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_start), .done(fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_done));
  assign fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_clk = clk;
  assign fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0_rst = rst;
  // Bindings to fused_level_3_fused_level_3_update_0_write0_to_final_merged_2_rd0

  // Bindings to fused_level_3_update_0_write_wdata
    // rd_1
  assign rd_1 = fused_level_3_update_0_write_wdata;

  // Bindings to fused_level_3_update_0_write_wen
    // rd_0
  assign rd_0 = fused_level_3_update_0_write_wen;

  // Bindings to final_merged_2_update_0_read_dummy
    // rd_2
  assign rd_2 = final_merged_2_update_0_read_dummy;

  // Bindings to final_merged_2_update_0_read_rdata
    // wr_3
  assign final_merged_2_update_0_read_rdata = rd_2;



endmodule


module in_in_update_0_write0_merged_banks_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module in(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] dark_update_0_read_dummy, output [31:0] bright_update_0_read_rdata, input [31:0] bright_update_0_read_dummy, input [0:0] in_update_0_write_wen, input [31:0] in_update_0_write_wdata, output [31:0] dark_update_0_read_rdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;
  logic [31:0] rd_2;
  logic [31:0] rd_4;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;
  reg [31:0] rd_4_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_4_stage_1 <= rd_4;


    end

  end


  // Data processing units...
  // Bindings to dark_update_0_read_dummy
    // rd_4
  assign rd_4 = dark_update_0_read_dummy;

  // Bindings to bright_update_0_read_rdata
    // wr_3
  assign bright_update_0_read_rdata = rd_2;

  // Bindings to bright_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_update_0_read_dummy;

  // Bindings to in_update_0_write_wen
    // rd_0
  assign rd_0 = in_update_0_write_wen;

  // Bindings to in_update_0_write_wdata
    // rd_1
  assign rd_1 = in_update_0_write_wdata;

  // in_in_update_0_write0_merged_banks_2
  logic [0:0] in_in_update_0_write0_merged_banks_2_clk;
  logic [0:0] in_in_update_0_write0_merged_banks_2_rst;
  logic [0:0] in_in_update_0_write0_merged_banks_2_start;
  logic [0:0] in_in_update_0_write0_merged_banks_2_done;
  in_in_update_0_write0_merged_banks_2 in_in_update_0_write0_merged_banks_2(.clk(in_in_update_0_write0_merged_banks_2_clk), .rst(in_in_update_0_write0_merged_banks_2_rst), .start(in_in_update_0_write0_merged_banks_2_start), .done(in_in_update_0_write0_merged_banks_2_done));
  assign in_in_update_0_write0_merged_banks_2_clk = clk;
  assign in_in_update_0_write0_merged_banks_2_rst = rst;
  // Bindings to in_in_update_0_write0_merged_banks_2

  // selector_bright_rd0_select
  logic [0:0] selector_bright_rd0_select_clk;
  logic [0:0] selector_bright_rd0_select_rst;
  logic [31:0] selector_bright_rd0_select_d0;
  logic [31:0] selector_bright_rd0_select_d1;
  logic [31:0] selector_bright_rd0_select_out;
  bright_rd0_select selector_bright_rd0_select(.clk(selector_bright_rd0_select_clk), .rst(selector_bright_rd0_select_rst), .d0(selector_bright_rd0_select_d0), .d1(selector_bright_rd0_select_d1), .out(selector_bright_rd0_select_out));
  assign selector_bright_rd0_select_clk = clk;
  assign selector_bright_rd0_select_rst = rst;
  // Bindings to selector_bright_rd0_select

  // selector_dark_rd0_select
  logic [0:0] selector_dark_rd0_select_clk;
  logic [0:0] selector_dark_rd0_select_rst;
  logic [31:0] selector_dark_rd0_select_d0;
  logic [31:0] selector_dark_rd0_select_d1;
  logic [31:0] selector_dark_rd0_select_out;
  dark_rd0_select selector_dark_rd0_select(.clk(selector_dark_rd0_select_clk), .rst(selector_dark_rd0_select_rst), .d0(selector_dark_rd0_select_d0), .d1(selector_dark_rd0_select_d1), .out(selector_dark_rd0_select_out));
  assign selector_dark_rd0_select_clk = clk;
  assign selector_dark_rd0_select_rst = rst;
  // Bindings to selector_dark_rd0_select

  // Bindings to dark_update_0_read_rdata
    // wr_5
  assign dark_update_0_read_rdata = rd_4;



endmodule


module in_wire_in_off_chip_update_0_write_wdata(output [31:0] in_off_chip_update_0_write_wdata);

endmodule


module in_wire_in_update_0_read_dummy(output [31:0] in_update_0_read_dummy);

endmodule


module out_wire_in_update_0_read_rdata(input [31:0] in_update_0_read_rdata);

endmodule


module pyramid_synthetic_exposure_fusion(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [0:0] pyramid_synthetic_exposure_fusion_update_0_write_wen, input [31:0] pyramid_synthetic_exposure_fusion_update_0_write_wdata);

  logic [0:0] rd_0;
  logic [31:0] rd_1;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [0:0] rd_0_stage_1;
  reg [31:0] rd_1_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;
      rd_1_stage_1 <= rd_1;


    end

  end


  // Data processing units...
  // Bindings to pyramid_synthetic_exposure_fusion_update_0_write_wen
    // rd_0
  assign rd_0 = pyramid_synthetic_exposure_fusion_update_0_write_wen;

  // Bindings to pyramid_synthetic_exposure_fusion_update_0_write_wdata
    // rd_1
  assign rd_1 = pyramid_synthetic_exposure_fusion_update_0_write_wdata;



endmodule


module in_wire_weight_sums_update_0_write_wen(output [0:0] weight_sums_update_0_write_wen);

endmodule


module in_wire_in_off_chip_update_0_write_wen(output [0:0] in_off_chip_update_0_write_wen);

endmodule


module bright_weights_normed_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_wire_weight_sums_update_0_write_wdata(output [31:0] weight_sums_update_0_write_wdata);

endmodule


module weight_sums_weight_sums_update_0_write0_merged_banks_2(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done);


  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end




    end

  end


  // Data processing units...
  // f1
  logic [0:0] f1_wen;
  logic [31:0] f1_wdata;
  logic [0:0] f1_clk;
  logic [0:0] f1_rst;
  logic [31:0] f1_rdata;
  sr_buffer_32_1 f1(.wen(f1_wen), .wdata(f1_wdata), .clk(f1_clk), .rst(f1_rst), .rdata(f1_rdata));
  assign f1_clk = clk;
  assign f1_rst = rst;
  // Bindings to f1



endmodule


module wire_32(input [31:0] in, output [31:0] out);
  assign out = in;
endmodule


module dark_weights_normed_rd0_select(input [0:0] clk, input [0:0] rst, input [31:0] d0, input [31:0] d1, output [31:0] out);
  always @(*) begin
    if (1) begin
      out = 0;
    end
  end

endmodule


module in_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module weight_sums(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, input [31:0] dark_weights_normed_update_0_read_dummy, input [0:0] weight_sums_update_0_write_wen, output [31:0] bright_weights_normed_update_0_read_rdata, input [31:0] bright_weights_normed_update_0_read_dummy, output [31:0] dark_weights_normed_update_0_read_rdata, input [31:0] weight_sums_update_0_write_wdata);

  logic [31:0] rd_4;
  logic [31:0] rd_1;
  logic [31:0] rd_2;
  logic [0:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_4_stage_1;
  reg [31:0] rd_1_stage_1;
  reg [31:0] rd_2_stage_1;
  reg [0:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_4_stage_1 <= rd_4;
      rd_1_stage_1 <= rd_1;
      rd_2_stage_1 <= rd_2;
      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to dark_weights_normed_update_0_read_dummy
    // rd_4
  assign rd_4 = dark_weights_normed_update_0_read_dummy;

  // selector_bright_weights_normed_rd0_select
  logic [0:0] selector_bright_weights_normed_rd0_select_clk;
  logic [0:0] selector_bright_weights_normed_rd0_select_rst;
  logic [31:0] selector_bright_weights_normed_rd0_select_d0;
  logic [31:0] selector_bright_weights_normed_rd0_select_d1;
  logic [31:0] selector_bright_weights_normed_rd0_select_out;
  bright_weights_normed_rd0_select selector_bright_weights_normed_rd0_select(.clk(selector_bright_weights_normed_rd0_select_clk), .rst(selector_bright_weights_normed_rd0_select_rst), .d0(selector_bright_weights_normed_rd0_select_d0), .d1(selector_bright_weights_normed_rd0_select_d1), .out(selector_bright_weights_normed_rd0_select_out));
  assign selector_bright_weights_normed_rd0_select_clk = clk;
  assign selector_bright_weights_normed_rd0_select_rst = rst;
  // Bindings to selector_bright_weights_normed_rd0_select

  // weight_sums_weight_sums_update_0_write0_merged_banks_2
  logic [0:0] weight_sums_weight_sums_update_0_write0_merged_banks_2_clk;
  logic [0:0] weight_sums_weight_sums_update_0_write0_merged_banks_2_rst;
  logic [0:0] weight_sums_weight_sums_update_0_write0_merged_banks_2_start;
  logic [0:0] weight_sums_weight_sums_update_0_write0_merged_banks_2_done;
  weight_sums_weight_sums_update_0_write0_merged_banks_2 weight_sums_weight_sums_update_0_write0_merged_banks_2(.clk(weight_sums_weight_sums_update_0_write0_merged_banks_2_clk), .rst(weight_sums_weight_sums_update_0_write0_merged_banks_2_rst), .start(weight_sums_weight_sums_update_0_write0_merged_banks_2_start), .done(weight_sums_weight_sums_update_0_write0_merged_banks_2_done));
  assign weight_sums_weight_sums_update_0_write0_merged_banks_2_clk = clk;
  assign weight_sums_weight_sums_update_0_write0_merged_banks_2_rst = rst;
  // Bindings to weight_sums_weight_sums_update_0_write0_merged_banks_2

  // Bindings to weight_sums_update_0_write_wen
    // rd_0
  assign rd_0 = weight_sums_update_0_write_wen;

  // Bindings to bright_weights_normed_update_0_read_rdata
    // wr_3
  assign bright_weights_normed_update_0_read_rdata = rd_2;

  // Bindings to bright_weights_normed_update_0_read_dummy
    // rd_2
  assign rd_2 = bright_weights_normed_update_0_read_dummy;

  // Bindings to dark_weights_normed_update_0_read_rdata
    // wr_5
  assign dark_weights_normed_update_0_read_rdata = rd_4;

  // Bindings to weight_sums_update_0_write_wdata
    // rd_1
  assign rd_1 = weight_sums_update_0_write_wdata;

  // selector_dark_weights_normed_rd0_select
  logic [0:0] selector_dark_weights_normed_rd0_select_clk;
  logic [0:0] selector_dark_weights_normed_rd0_select_rst;
  logic [31:0] selector_dark_weights_normed_rd0_select_d0;
  logic [31:0] selector_dark_weights_normed_rd0_select_d1;
  logic [31:0] selector_dark_weights_normed_rd0_select_out;
  dark_weights_normed_rd0_select selector_dark_weights_normed_rd0_select(.clk(selector_dark_weights_normed_rd0_select_clk), .rst(selector_dark_weights_normed_rd0_select_rst), .d0(selector_dark_weights_normed_rd0_select_d0), .d1(selector_dark_weights_normed_rd0_select_d1), .out(selector_dark_weights_normed_rd0_select_out));
  assign selector_dark_weights_normed_rd0_select_clk = clk;
  assign selector_dark_weights_normed_rd0_select_rst = rst;
  // Bindings to selector_dark_weights_normed_rd0_select



endmodule


module out_wire_out(input [31:0] out);

endmodule


module dark_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_gauss_ds_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_weights_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module dark_weights_normed_gauss_ds_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_laplace_diff_0_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module fused_level_0_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_weights_normed_gauss_ds_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module bright_weights_normed_gauss_blur_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_gauss_blur_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_laplace_us_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_laplace_diff_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module fused_level_1_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] out, output [31:0] src_in, input [31:0] src_out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to out
    // wr_1
  assign out = rd_0;

  // Bindings to src
    // rd_0
  assign rd_0 = src_out;



endmodule


module bright_weights_normed_gauss_ds_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_weights_normed_gauss_blur_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_gauss_ds_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_laplace_us_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_laplace_diff_2_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule


module bright_weights_normed_gauss_ds_3_update_0(input [0:0] clk, input [0:0] rst, input [0:0] start, output [0:0] done, output [31:0] src_in, input [31:0] src_out, output [31:0] out);

  logic [31:0] rd_0;

  logic started;

  logic stage_0_active;

  logic stage_0_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_0_active;

  // Pipeline datapath registers...
  reg [31:0] rd_0_stage_1;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end


      rd_0_stage_1 <= rd_0;


    end

  end


  // Data processing units...
  // Bindings to src
    // rd_0
  assign rd_0 = src_out;

  // Bindings to out
    // wr_1
  assign out = rd_0;



endmodule



