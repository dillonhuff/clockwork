// Module `hw_kernel_global_wrapper_stencil_ub` defined externally
// Module `hw_input_global_wrapper_stencil_ub` defined externally
// Module `conv_stencil_ub` defined externally
module op_hcompute_hw_output_stencil_write_start_pt__U34 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_write_start_control_vars_pt__U36 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_read_start_pt__U23 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_read_start_control_vars_pt__U24 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_exe_start_pt__U25 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U27 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U100 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U101 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U96 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U97 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U98 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U99 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U129 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U130 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U125 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U126 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U127 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U128 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_write_start_pt__U64 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_write_start_control_vars_pt__U65 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_read_start_pt__U60 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_read_start_control_vars_pt__U61 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_exe_start_pt__U62 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_exe_start_control_vars_pt__U63 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_write_start_pt__U323 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_write_start_control_vars_pt__U325 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_read_start_pt__U311 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_read_start_control_vars_pt__U312 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_exe_start_pt__U313 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U315 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_write_start_pt__U271 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_write_start_control_vars_pt__U273 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_read_start_pt__U259 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_read_start_control_vars_pt__U260 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_exe_start_pt__U261 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U263 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_write_start_pt__U219 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_write_start_control_vars_pt__U221 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_read_start_pt__U207 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_read_start_control_vars_pt__U208 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_exe_start_pt__U209 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U211 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_write_start_pt__U175 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_write_start_control_vars_pt__U176 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_read_start_pt__U171 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_read_start_control_vars_pt__U172 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_exe_start_pt__U173 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U174 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_write_start_pt__U152 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_write_start_control_vars_pt__U153 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_read_start_pt__U148 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_read_start_control_vars_pt__U149 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_exe_start_pt__U150 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U151 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module hcompute_hw_output_stencil (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
assign out_hw_output_stencil = in0_conv_stencil[0];
endmodule

module hcompute_hw_kernel_global_wrapper_stencil (
    output [15:0] out_hw_kernel_global_wrapper_stencil,
    input [15:0] in0_hw_kernel_stencil [0:0]
);
assign out_hw_kernel_global_wrapper_stencil = in0_hw_kernel_stencil[0];
endmodule

module hcompute_hw_input_global_wrapper_stencil (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
assign out_hw_input_global_wrapper_stencil = in0_hw_input_stencil[0];
endmodule

module cu_op_hcompute_hw_output_stencil (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0],
    output [15:0] hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
hcompute_hw_output_stencil inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_op_hcompute_hw_output_stencil_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module cu_op_hcompute_hw_kernel_global_wrapper_stencil (
    input clk,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_kernel_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_kernel_stencil [0:0];
assign inner_compute_in0_hw_kernel_stencil[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
hcompute_hw_kernel_global_wrapper_stencil inner_compute (
    .out_hw_kernel_global_wrapper_stencil(inner_compute_out_hw_kernel_global_wrapper_stencil),
    .in0_hw_kernel_stencil(inner_compute_in0_hw_kernel_stencil)
);
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = inner_compute_out_hw_kernel_global_wrapper_stencil;
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil (
    input clk,
    input [15:0] hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0];
hcompute_hw_input_global_wrapper_stencil inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module coreir_reg #(
    parameter width = 1,
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input [width-1:0] in,
    output [width-1:0] out
);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out
);
wire reg0_clk;
wire [15:0] reg0_in;
assign reg0_clk = clk;
assign reg0_in = in;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(reg0_clk),
    .in(reg0_in),
    .out(out)
);
endmodule

module mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out,
    input en
);
wire reg0_clk;
wire [15:0] reg0_in;
assign reg0_clk = clk;
assign reg0_in = en ? in : out;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(reg0_clk),
    .in(reg0_in),
    .out(out)
);
endmodule

module hcompute_conv_stencil_2 (
    output [15:0] out_conv_stencil
);
assign out_conv_stencil = 16'h0000;
endmodule

module cu_op_hcompute_conv_stencil_2 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_2 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_1 (
    output [15:0] out_conv_stencil
);
assign out_conv_stencil = 16'h0000;
endmodule

module cu_op_hcompute_conv_stencil_1 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_1 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil (
    output [15:0] out_conv_stencil
);
assign out_conv_stencil = 16'h0000;
endmodule

module cu_op_hcompute_conv_stencil (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_5 (
    output [15:0] out_conv_stencil,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0]
);
assign out_conv_stencil = 16'((16'(in2_hw_kernel_global_wrapper_stencil[0] * in1_hw_input_global_wrapper_stencil[0])) + (16'(in0_conv_stencil[0] + (16'((16'(in2_hw_kernel_global_wrapper_stencil[1] * in1_hw_input_global_wrapper_stencil[1])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[2] * in1_hw_input_global_wrapper_stencil[2])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[3] * in1_hw_input_global_wrapper_stencil[3])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[4] * in1_hw_input_global_wrapper_stencil[4])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[5] * in1_hw_input_global_wrapper_stencil[5])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[6] * in1_hw_input_global_wrapper_stencil[6])) + (16'(in2_hw_kernel_global_wrapper_stencil[7] * in1_hw_input_global_wrapper_stencil[7])))))))))))))))));
endmodule

module cu_op_hcompute_conv_stencil_5 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_5_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_5_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
hcompute_conv_stencil_5 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_4 (
    output [15:0] out_conv_stencil,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0]
);
assign out_conv_stencil = 16'((16'(in2_hw_kernel_global_wrapper_stencil[7] * in1_hw_input_global_wrapper_stencil[7])) + (16'(in0_conv_stencil[0] + (16'((16'(in2_hw_kernel_global_wrapper_stencil[0] * in1_hw_input_global_wrapper_stencil[0])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[1] * in1_hw_input_global_wrapper_stencil[1])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[2] * in1_hw_input_global_wrapper_stencil[2])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[3] * in1_hw_input_global_wrapper_stencil[3])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[4] * in1_hw_input_global_wrapper_stencil[4])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[5] * in1_hw_input_global_wrapper_stencil[5])) + (16'(in2_hw_kernel_global_wrapper_stencil[6] * in1_hw_input_global_wrapper_stencil[6])))))))))))))))));
endmodule

module cu_op_hcompute_conv_stencil_4 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_4_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_4_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
hcompute_conv_stencil_4 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_3 (
    output [15:0] out_conv_stencil,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0]
);
assign out_conv_stencil = 16'((16'(in2_hw_kernel_global_wrapper_stencil[0] * in1_hw_input_global_wrapper_stencil[0])) + (16'(in0_conv_stencil[0] + (16'((16'(in2_hw_kernel_global_wrapper_stencil[1] * in1_hw_input_global_wrapper_stencil[1])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[2] * in1_hw_input_global_wrapper_stencil[2])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[3] * in1_hw_input_global_wrapper_stencil[3])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[4] * in1_hw_input_global_wrapper_stencil[4])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[5] * in1_hw_input_global_wrapper_stencil[5])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[6] * in1_hw_input_global_wrapper_stencil[6])) + (16'(in2_hw_kernel_global_wrapper_stencil[7] * in1_hw_input_global_wrapper_stencil[7])))))))))))))))));
endmodule

module cu_op_hcompute_conv_stencil_3 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_3_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_3_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
hcompute_conv_stencil_3 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = inner_compute_out_conv_stencil;
endmodule

module corebit_reg #(
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input in,
    output out
);
reg outReg = init;
always @(posedge clk) begin
  outReg <= in;
end
assign out = outReg;
endmodule

module array_delay_U38 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U39_in;
wire _U39_clk;
wire [15:0] _U39_out;
wire [15:0] _U40_in;
wire _U40_clk;
wire [15:0] _U40_out;
wire [15:0] _U41_in;
wire _U41_clk;
wire [15:0] _U41_out;
wire [15:0] _U42_in;
wire _U42_clk;
wire [15:0] _U42_out;
assign _U39_in = in[0];
assign _U39_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U39 (
    .in(_U39_in),
    .clk(_U39_clk),
    .out(_U39_out)
);
assign _U40_in = in[1];
assign _U40_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U40 (
    .in(_U40_in),
    .clk(_U40_clk),
    .out(_U40_out)
);
assign _U41_in = in[2];
assign _U41_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U41 (
    .in(_U41_in),
    .clk(_U41_clk),
    .out(_U41_out)
);
assign _U42_in = in[3];
assign _U42_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U42 (
    .in(_U42_in),
    .clk(_U42_clk),
    .out(_U42_out)
);
assign out[3] = _U42_out;
assign out[2] = _U41_out;
assign out[1] = _U40_out;
assign out[0] = _U39_out;
endmodule

module array_delay_U327 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U328_in;
wire _U328_clk;
wire [15:0] _U328_out;
wire [15:0] _U329_in;
wire _U329_clk;
wire [15:0] _U329_out;
wire [15:0] _U330_in;
wire _U330_clk;
wire [15:0] _U330_out;
wire [15:0] _U331_in;
wire _U331_clk;
wire [15:0] _U331_out;
wire [15:0] _U332_in;
wire _U332_clk;
wire [15:0] _U332_out;
assign _U328_in = in[0];
assign _U328_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U328 (
    .in(_U328_in),
    .clk(_U328_clk),
    .out(_U328_out)
);
assign _U329_in = in[1];
assign _U329_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U329 (
    .in(_U329_in),
    .clk(_U329_clk),
    .out(_U329_out)
);
assign _U330_in = in[2];
assign _U330_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U330 (
    .in(_U330_in),
    .clk(_U330_clk),
    .out(_U330_out)
);
assign _U331_in = in[3];
assign _U331_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U331 (
    .in(_U331_in),
    .clk(_U331_clk),
    .out(_U331_out)
);
assign _U332_in = in[4];
assign _U332_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U332 (
    .in(_U332_in),
    .clk(_U332_clk),
    .out(_U332_out)
);
assign out[4] = _U332_out;
assign out[3] = _U331_out;
assign out[2] = _U330_out;
assign out[1] = _U329_out;
assign out[0] = _U328_out;
endmodule

module array_delay_U317 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U318_in;
wire _U318_clk;
wire [15:0] _U318_out;
wire [15:0] _U319_in;
wire _U319_clk;
wire [15:0] _U319_out;
wire [15:0] _U320_in;
wire _U320_clk;
wire [15:0] _U320_out;
wire [15:0] _U321_in;
wire _U321_clk;
wire [15:0] _U321_out;
wire [15:0] _U322_in;
wire _U322_clk;
wire [15:0] _U322_out;
assign _U318_in = in[0];
assign _U318_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U318 (
    .in(_U318_in),
    .clk(_U318_clk),
    .out(_U318_out)
);
assign _U319_in = in[1];
assign _U319_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U319 (
    .in(_U319_in),
    .clk(_U319_clk),
    .out(_U319_out)
);
assign _U320_in = in[2];
assign _U320_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U320 (
    .in(_U320_in),
    .clk(_U320_clk),
    .out(_U320_out)
);
assign _U321_in = in[3];
assign _U321_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U321 (
    .in(_U321_in),
    .clk(_U321_clk),
    .out(_U321_out)
);
assign _U322_in = in[4];
assign _U322_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U322 (
    .in(_U322_in),
    .clk(_U322_clk),
    .out(_U322_out)
);
assign out[4] = _U322_out;
assign out[3] = _U321_out;
assign out[2] = _U320_out;
assign out[1] = _U319_out;
assign out[0] = _U318_out;
endmodule

module array_delay_U29 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U30_in;
wire _U30_clk;
wire [15:0] _U30_out;
wire [15:0] _U31_in;
wire _U31_clk;
wire [15:0] _U31_out;
wire [15:0] _U32_in;
wire _U32_clk;
wire [15:0] _U32_out;
wire [15:0] _U33_in;
wire _U33_clk;
wire [15:0] _U33_out;
assign _U30_in = in[0];
assign _U30_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U30 (
    .in(_U30_in),
    .clk(_U30_clk),
    .out(_U30_out)
);
assign _U31_in = in[1];
assign _U31_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U31 (
    .in(_U31_in),
    .clk(_U31_clk),
    .out(_U31_out)
);
assign _U32_in = in[2];
assign _U32_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U32 (
    .in(_U32_in),
    .clk(_U32_clk),
    .out(_U32_out)
);
assign _U33_in = in[3];
assign _U33_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U33 (
    .in(_U33_in),
    .clk(_U33_clk),
    .out(_U33_out)
);
assign out[3] = _U33_out;
assign out[2] = _U32_out;
assign out[1] = _U31_out;
assign out[0] = _U30_out;
endmodule

module array_delay_U275 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U276_in;
wire _U276_clk;
wire [15:0] _U276_out;
wire [15:0] _U277_in;
wire _U277_clk;
wire [15:0] _U277_out;
wire [15:0] _U278_in;
wire _U278_clk;
wire [15:0] _U278_out;
wire [15:0] _U279_in;
wire _U279_clk;
wire [15:0] _U279_out;
wire [15:0] _U280_in;
wire _U280_clk;
wire [15:0] _U280_out;
assign _U276_in = in[0];
assign _U276_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U276 (
    .in(_U276_in),
    .clk(_U276_clk),
    .out(_U276_out)
);
assign _U277_in = in[1];
assign _U277_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U277 (
    .in(_U277_in),
    .clk(_U277_clk),
    .out(_U277_out)
);
assign _U278_in = in[2];
assign _U278_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U278 (
    .in(_U278_in),
    .clk(_U278_clk),
    .out(_U278_out)
);
assign _U279_in = in[3];
assign _U279_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U279 (
    .in(_U279_in),
    .clk(_U279_clk),
    .out(_U279_out)
);
assign _U280_in = in[4];
assign _U280_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U280 (
    .in(_U280_in),
    .clk(_U280_clk),
    .out(_U280_out)
);
assign out[4] = _U280_out;
assign out[3] = _U279_out;
assign out[2] = _U278_out;
assign out[1] = _U277_out;
assign out[0] = _U276_out;
endmodule

module array_delay_U265 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U266_in;
wire _U266_clk;
wire [15:0] _U266_out;
wire [15:0] _U267_in;
wire _U267_clk;
wire [15:0] _U267_out;
wire [15:0] _U268_in;
wire _U268_clk;
wire [15:0] _U268_out;
wire [15:0] _U269_in;
wire _U269_clk;
wire [15:0] _U269_out;
wire [15:0] _U270_in;
wire _U270_clk;
wire [15:0] _U270_out;
assign _U266_in = in[0];
assign _U266_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U266 (
    .in(_U266_in),
    .clk(_U266_clk),
    .out(_U266_out)
);
assign _U267_in = in[1];
assign _U267_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U267 (
    .in(_U267_in),
    .clk(_U267_clk),
    .out(_U267_out)
);
assign _U268_in = in[2];
assign _U268_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U268 (
    .in(_U268_in),
    .clk(_U268_clk),
    .out(_U268_out)
);
assign _U269_in = in[3];
assign _U269_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U269 (
    .in(_U269_in),
    .clk(_U269_clk),
    .out(_U269_out)
);
assign _U270_in = in[4];
assign _U270_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U270 (
    .in(_U270_in),
    .clk(_U270_clk),
    .out(_U270_out)
);
assign out[4] = _U270_out;
assign out[3] = _U269_out;
assign out[2] = _U268_out;
assign out[1] = _U267_out;
assign out[0] = _U266_out;
endmodule

module array_delay_U223 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U224_in;
wire _U224_clk;
wire [15:0] _U224_out;
wire [15:0] _U225_in;
wire _U225_clk;
wire [15:0] _U225_out;
wire [15:0] _U226_in;
wire _U226_clk;
wire [15:0] _U226_out;
wire [15:0] _U227_in;
wire _U227_clk;
wire [15:0] _U227_out;
wire [15:0] _U228_in;
wire _U228_clk;
wire [15:0] _U228_out;
assign _U224_in = in[0];
assign _U224_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U224 (
    .in(_U224_in),
    .clk(_U224_clk),
    .out(_U224_out)
);
assign _U225_in = in[1];
assign _U225_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U225 (
    .in(_U225_in),
    .clk(_U225_clk),
    .out(_U225_out)
);
assign _U226_in = in[2];
assign _U226_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U226 (
    .in(_U226_in),
    .clk(_U226_clk),
    .out(_U226_out)
);
assign _U227_in = in[3];
assign _U227_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U227 (
    .in(_U227_in),
    .clk(_U227_clk),
    .out(_U227_out)
);
assign _U228_in = in[4];
assign _U228_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U228 (
    .in(_U228_in),
    .clk(_U228_clk),
    .out(_U228_out)
);
assign out[4] = _U228_out;
assign out[3] = _U227_out;
assign out[2] = _U226_out;
assign out[1] = _U225_out;
assign out[0] = _U224_out;
endmodule

module array_delay_U213 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U214_in;
wire _U214_clk;
wire [15:0] _U214_out;
wire [15:0] _U215_in;
wire _U215_clk;
wire [15:0] _U215_out;
wire [15:0] _U216_in;
wire _U216_clk;
wire [15:0] _U216_out;
wire [15:0] _U217_in;
wire _U217_clk;
wire [15:0] _U217_out;
wire [15:0] _U218_in;
wire _U218_clk;
wire [15:0] _U218_out;
assign _U214_in = in[0];
assign _U214_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U214 (
    .in(_U214_in),
    .clk(_U214_clk),
    .out(_U214_out)
);
assign _U215_in = in[1];
assign _U215_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U215 (
    .in(_U215_in),
    .clk(_U215_clk),
    .out(_U215_out)
);
assign _U216_in = in[2];
assign _U216_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U216 (
    .in(_U216_in),
    .clk(_U216_clk),
    .out(_U216_out)
);
assign _U217_in = in[3];
assign _U217_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U217 (
    .in(_U217_in),
    .clk(_U217_clk),
    .out(_U217_out)
);
assign _U218_in = in[4];
assign _U218_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U218 (
    .in(_U218_in),
    .clk(_U218_clk),
    .out(_U218_out)
);
assign out[4] = _U218_out;
assign out[3] = _U217_out;
assign out[2] = _U216_out;
assign out[1] = _U215_out;
assign out[0] = _U214_out;
endmodule

module aff__U67 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0048 * d[1])))) + (16'(16'h0018 * d[2])))) + (16'(16'h0008 * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h0002);
endmodule

module affine_controller__U66 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U67 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h0002;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h0007;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U44 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001c * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U43 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U44 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U282 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0984 * d[1])))) + (16'(16'h032c * d[2])))) + (16'(16'h001d * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h1f49);
endmodule

module affine_controller__U281 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U282 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U230 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0984 * d[1])))) + (16'(16'h032c * d[2])))) + (16'(16'h001d * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h1f49);
endmodule

module affine_controller__U229 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U230 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U178 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0984 * d[1])))) + (16'(16'h032c * d[2])))) + (16'(16'h001d * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h1f49);
endmodule

module affine_controller__U177 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U178 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U155 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001c * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U154 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U155 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U132 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001c * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U131 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U132 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U103 (
    output [15:0] out,
    input [15:0] d [3:0]
);
assign out = 16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h00f0 * d[1])))) + (16'(16'h0008 * d[2])))) + (16'(16'h0001 * d[3])))) + 16'h0001);
endmodule

module affine_controller__U102 (
    input clk,
    output valid,
    output [15:0] d [3:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [3:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U103 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = ((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_reg_in = (1'b1 & d_2_at_max_out) & d_3_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_reg_in = 1'b1 & d_3_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h0007;
assign d_3_reg_in = 1'b1 ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign valid = cmp_time_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1 (
    output [15:0] out,
    input [15:0] d [3:0]
);
assign out = 16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0310 * d[1])))) + (16'(16'h001c * d[2])))) + (16'(16'h0001 * d[3])))) + 16'h3e91);
endmodule

module affine_controller__U0 (
    input clk,
    output valid,
    output [15:0] d [3:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [3:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = ((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = (1'b1 & d_2_at_max_out) & d_3_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 & d_3_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign valid = cmp_time_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module resnet (
    input clk,
    input rst_n,
    input flush,
    output hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read_en,
    input [15:0] hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output hw_output_stencil_op_hcompute_hw_output_stencil_write_valid,
    output [15:0] hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0]
);
wire arr__U212_clk;
wire [15:0] arr__U212_in [4:0];
wire [15:0] arr__U212_out [4:0];
wire arr__U222_clk;
wire [15:0] arr__U222_in [4:0];
wire [15:0] arr__U222_out [4:0];
wire arr__U264_clk;
wire [15:0] arr__U264_in [4:0];
wire [15:0] arr__U264_out [4:0];
wire arr__U274_clk;
wire [15:0] arr__U274_in [4:0];
wire [15:0] arr__U274_out [4:0];
wire arr__U28_clk;
wire [15:0] arr__U28_in [3:0];
wire [15:0] arr__U28_out [3:0];
wire arr__U316_clk;
wire [15:0] arr__U316_in [4:0];
wire [15:0] arr__U316_out [4:0];
wire arr__U326_clk;
wire [15:0] arr__U326_in [4:0];
wire [15:0] arr__U326_out [4:0];
wire arr__U37_clk;
wire [15:0] arr__U37_in [3:0];
wire [15:0] arr__U37_out [3:0];
wire conv_stencil_clk;
wire conv_stencil_flush;
wire conv_stencil_rst_n;
wire conv_stencil_op_hcompute_conv_stencil_1_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_2_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_3_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_4_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_5_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire conv_stencil_op_hcompute_hw_output_stencil_read_ren;
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars [3:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire delay_reg__U210_clk;
wire delay_reg__U210_in;
wire delay_reg__U210_out;
wire delay_reg__U220_clk;
wire delay_reg__U220_in;
wire delay_reg__U220_out;
wire delay_reg__U26_clk;
wire delay_reg__U26_in;
wire delay_reg__U26_out;
wire delay_reg__U262_clk;
wire delay_reg__U262_in;
wire delay_reg__U262_out;
wire delay_reg__U272_clk;
wire delay_reg__U272_in;
wire delay_reg__U272_out;
wire delay_reg__U314_clk;
wire delay_reg__U314_in;
wire delay_reg__U314_out;
wire delay_reg__U324_clk;
wire delay_reg__U324_in;
wire delay_reg__U324_out;
wire delay_reg__U35_clk;
wire delay_reg__U35_in;
wire delay_reg__U35_out;
wire hw_input_global_wrapper_stencil_clk;
wire hw_input_global_wrapper_stencil_flush;
wire hw_input_global_wrapper_stencil_rst_n;
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars [3:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire hw_kernel_global_wrapper_stencil_clk;
wire hw_kernel_global_wrapper_stencil_flush;
wire hw_kernel_global_wrapper_stencil_rst_n;
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_conv_stencil_clk;
wire [15:0] op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire op_hcompute_conv_stencil_1_clk;
wire [15:0] op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire op_hcompute_conv_stencil_1_exe_start_in;
wire op_hcompute_conv_stencil_1_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_port_controller_clk;
wire op_hcompute_conv_stencil_1_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_1_port_controller_d [2:0];
wire op_hcompute_conv_stencil_1_read_start_in;
wire op_hcompute_conv_stencil_1_read_start_out;
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_write_start_in;
wire op_hcompute_conv_stencil_1_write_start_out;
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_clk;
wire [15:0] op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire op_hcompute_conv_stencil_2_exe_start_in;
wire op_hcompute_conv_stencil_2_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_port_controller_clk;
wire op_hcompute_conv_stencil_2_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_2_port_controller_d [2:0];
wire op_hcompute_conv_stencil_2_read_start_in;
wire op_hcompute_conv_stencil_2_read_start_out;
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_write_start_in;
wire op_hcompute_conv_stencil_2_write_start_out;
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_3_clk;
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read [0:0];
wire [15:0] op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire [15:0] op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire op_hcompute_conv_stencil_3_exe_start_in;
wire op_hcompute_conv_stencil_3_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_3_port_controller_clk;
wire op_hcompute_conv_stencil_3_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_3_port_controller_d [4:0];
wire op_hcompute_conv_stencil_3_read_start_in;
wire op_hcompute_conv_stencil_3_read_start_out;
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_3_write_start_in;
wire op_hcompute_conv_stencil_3_write_start_out;
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_clk;
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read [0:0];
wire [15:0] op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire [15:0] op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire op_hcompute_conv_stencil_4_exe_start_in;
wire op_hcompute_conv_stencil_4_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_port_controller_clk;
wire op_hcompute_conv_stencil_4_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_4_port_controller_d [4:0];
wire op_hcompute_conv_stencil_4_read_start_in;
wire op_hcompute_conv_stencil_4_read_start_out;
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_write_start_in;
wire op_hcompute_conv_stencil_4_write_start_out;
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_clk;
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read [0:0];
wire [15:0] op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire [15:0] op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire op_hcompute_conv_stencil_5_exe_start_in;
wire op_hcompute_conv_stencil_5_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_port_controller_clk;
wire op_hcompute_conv_stencil_5_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_5_port_controller_d [4:0];
wire op_hcompute_conv_stencil_5_read_start_in;
wire op_hcompute_conv_stencil_5_read_start_out;
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_write_start_in;
wire op_hcompute_conv_stencil_5_write_start_out;
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_exe_start_in;
wire op_hcompute_conv_stencil_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_port_controller_clk;
wire op_hcompute_conv_stencil_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_port_controller_d [2:0];
wire op_hcompute_conv_stencil_read_start_in;
wire op_hcompute_conv_stencil_read_start_out;
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_write_start_in;
wire op_hcompute_conv_stencil_write_start_out;
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_clk;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk;
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_port_controller_d [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_read_start_in;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out [3:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_clk;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in;
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk;
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in;
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out [4:0];
wire op_hcompute_hw_output_stencil_clk;
wire [15:0] op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire [15:0] op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0];
wire op_hcompute_hw_output_stencil_exe_start_in;
wire op_hcompute_hw_output_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_out [3:0];
wire op_hcompute_hw_output_stencil_port_controller_clk;
wire op_hcompute_hw_output_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_port_controller_d [3:0];
wire op_hcompute_hw_output_stencil_read_start_in;
wire op_hcompute_hw_output_stencil_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_out [3:0];
wire op_hcompute_hw_output_stencil_write_start_in;
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_out [3:0];
assign arr__U212_clk = clk;
assign arr__U212_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign arr__U212_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign arr__U212_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign arr__U212_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign arr__U212_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
array_delay_U213 arr__U212 (
    .clk(arr__U212_clk),
    .in(arr__U212_in),
    .out(arr__U212_out)
);
assign arr__U222_clk = clk;
assign arr__U222_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign arr__U222_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign arr__U222_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign arr__U222_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign arr__U222_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
array_delay_U223 arr__U222 (
    .clk(arr__U222_clk),
    .in(arr__U222_in),
    .out(arr__U222_out)
);
assign arr__U264_clk = clk;
assign arr__U264_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign arr__U264_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign arr__U264_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign arr__U264_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign arr__U264_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
array_delay_U265 arr__U264 (
    .clk(arr__U264_clk),
    .in(arr__U264_in),
    .out(arr__U264_out)
);
assign arr__U274_clk = clk;
assign arr__U274_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign arr__U274_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign arr__U274_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign arr__U274_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign arr__U274_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
array_delay_U275 arr__U274 (
    .clk(arr__U274_clk),
    .in(arr__U274_in),
    .out(arr__U274_out)
);
assign arr__U28_clk = clk;
assign arr__U28_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign arr__U28_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U28_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U28_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U29 arr__U28 (
    .clk(arr__U28_clk),
    .in(arr__U28_in),
    .out(arr__U28_out)
);
assign arr__U316_clk = clk;
assign arr__U316_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign arr__U316_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign arr__U316_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign arr__U316_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign arr__U316_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
array_delay_U317 arr__U316 (
    .clk(arr__U316_clk),
    .in(arr__U316_in),
    .out(arr__U316_out)
);
assign arr__U326_clk = clk;
assign arr__U326_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign arr__U326_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign arr__U326_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign arr__U326_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign arr__U326_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
array_delay_U327 arr__U326 (
    .clk(arr__U326_clk),
    .in(arr__U326_in),
    .out(arr__U326_out)
);
assign arr__U37_clk = clk;
assign arr__U37_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign arr__U37_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U37_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U37_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U38 arr__U37 (
    .clk(arr__U37_clk),
    .in(arr__U37_in),
    .out(arr__U37_out)
);
assign conv_stencil_clk = clk;
assign conv_stencil_flush = flush;
assign conv_stencil_rst_n = rst_n;
assign conv_stencil_op_hcompute_conv_stencil_1_write_wen = op_hcompute_conv_stencil_1_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[2] = op_hcompute_conv_stencil_1_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[1] = op_hcompute_conv_stencil_1_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[0] = op_hcompute_conv_stencil_1_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write[0];
assign conv_stencil_op_hcompute_conv_stencil_2_write_wen = op_hcompute_conv_stencil_2_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[2] = op_hcompute_conv_stencil_2_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[1] = op_hcompute_conv_stencil_2_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[0] = op_hcompute_conv_stencil_2_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write[0];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_3_write_wen = op_hcompute_conv_stencil_3_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[4] = op_hcompute_conv_stencil_3_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[3] = op_hcompute_conv_stencil_3_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[2] = op_hcompute_conv_stencil_3_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[1] = op_hcompute_conv_stencil_3_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[0] = op_hcompute_conv_stencil_3_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write[0];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_4_write_wen = op_hcompute_conv_stencil_4_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[4] = op_hcompute_conv_stencil_4_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[3] = op_hcompute_conv_stencil_4_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[2] = op_hcompute_conv_stencil_4_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[1] = op_hcompute_conv_stencil_4_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[0] = op_hcompute_conv_stencil_4_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write[0];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_5_write_wen = op_hcompute_conv_stencil_5_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[4] = op_hcompute_conv_stencil_5_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[3] = op_hcompute_conv_stencil_5_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[2] = op_hcompute_conv_stencil_5_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[1] = op_hcompute_conv_stencil_5_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[0] = op_hcompute_conv_stencil_5_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write[0];
assign conv_stencil_op_hcompute_conv_stencil_write_wen = op_hcompute_conv_stencil_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[2] = op_hcompute_conv_stencil_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[1] = op_hcompute_conv_stencil_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[0] = op_hcompute_conv_stencil_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_write[0] = op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write[0];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ren = op_hcompute_hw_output_stencil_read_start_out;
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
conv_stencil_ub conv_stencil (
    .clk(conv_stencil_clk),
    .flush(conv_stencil_flush),
    .rst_n(conv_stencil_rst_n),
    .op_hcompute_conv_stencil_1_write_wen(conv_stencil_op_hcompute_conv_stencil_1_write_wen),
    .op_hcompute_conv_stencil_1_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars),
    .op_hcompute_conv_stencil_1_write(conv_stencil_op_hcompute_conv_stencil_1_write),
    .op_hcompute_conv_stencil_2_write_wen(conv_stencil_op_hcompute_conv_stencil_2_write_wen),
    .op_hcompute_conv_stencil_2_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars),
    .op_hcompute_conv_stencil_2_write(conv_stencil_op_hcompute_conv_stencil_2_write),
    .op_hcompute_conv_stencil_3_read_ren(conv_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(conv_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_3_write_wen(conv_stencil_op_hcompute_conv_stencil_3_write_wen),
    .op_hcompute_conv_stencil_3_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars),
    .op_hcompute_conv_stencil_3_write(conv_stencil_op_hcompute_conv_stencil_3_write),
    .op_hcompute_conv_stencil_4_read_ren(conv_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(conv_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_4_write_wen(conv_stencil_op_hcompute_conv_stencil_4_write_wen),
    .op_hcompute_conv_stencil_4_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars),
    .op_hcompute_conv_stencil_4_write(conv_stencil_op_hcompute_conv_stencil_4_write),
    .op_hcompute_conv_stencil_5_read_ren(conv_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(conv_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_conv_stencil_5_write_wen(conv_stencil_op_hcompute_conv_stencil_5_write_wen),
    .op_hcompute_conv_stencil_5_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars),
    .op_hcompute_conv_stencil_5_write(conv_stencil_op_hcompute_conv_stencil_5_write),
    .op_hcompute_conv_stencil_write_wen(conv_stencil_op_hcompute_conv_stencil_write_wen),
    .op_hcompute_conv_stencil_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars),
    .op_hcompute_conv_stencil_write(conv_stencil_op_hcompute_conv_stencil_write),
    .op_hcompute_hw_output_stencil_read_ren(conv_stencil_op_hcompute_hw_output_stencil_read_ren),
    .op_hcompute_hw_output_stencil_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_read(conv_stencil_op_hcompute_hw_output_stencil_read)
);
assign delay_reg__U210_clk = clk;
assign delay_reg__U210_in = op_hcompute_conv_stencil_3_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U210 (
    .clk(delay_reg__U210_clk),
    .in(delay_reg__U210_in),
    .out(delay_reg__U210_out)
);
assign delay_reg__U220_clk = clk;
assign delay_reg__U220_in = op_hcompute_conv_stencil_3_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U220 (
    .clk(delay_reg__U220_clk),
    .in(delay_reg__U220_in),
    .out(delay_reg__U220_out)
);
assign delay_reg__U26_clk = clk;
assign delay_reg__U26_in = op_hcompute_hw_output_stencil_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U26 (
    .clk(delay_reg__U26_clk),
    .in(delay_reg__U26_in),
    .out(delay_reg__U26_out)
);
assign delay_reg__U262_clk = clk;
assign delay_reg__U262_in = op_hcompute_conv_stencil_4_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U262 (
    .clk(delay_reg__U262_clk),
    .in(delay_reg__U262_in),
    .out(delay_reg__U262_out)
);
assign delay_reg__U272_clk = clk;
assign delay_reg__U272_in = op_hcompute_conv_stencil_4_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U272 (
    .clk(delay_reg__U272_clk),
    .in(delay_reg__U272_in),
    .out(delay_reg__U272_out)
);
assign delay_reg__U314_clk = clk;
assign delay_reg__U314_in = op_hcompute_conv_stencil_5_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U314 (
    .clk(delay_reg__U314_clk),
    .in(delay_reg__U314_in),
    .out(delay_reg__U314_out)
);
assign delay_reg__U324_clk = clk;
assign delay_reg__U324_in = op_hcompute_conv_stencil_5_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U324 (
    .clk(delay_reg__U324_clk),
    .in(delay_reg__U324_in),
    .out(delay_reg__U324_out)
);
assign delay_reg__U35_clk = clk;
assign delay_reg__U35_in = op_hcompute_hw_output_stencil_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U35 (
    .clk(delay_reg__U35_clk),
    .in(delay_reg__U35_in),
    .out(delay_reg__U35_out)
);
assign hw_input_global_wrapper_stencil_clk = clk;
assign hw_input_global_wrapper_stencil_flush = flush;
assign hw_input_global_wrapper_stencil_rst_n = rst_n;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen = op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0];
hw_input_global_wrapper_stencil_ub hw_input_global_wrapper_stencil (
    .clk(hw_input_global_wrapper_stencil_clk),
    .flush(hw_input_global_wrapper_stencil_flush),
    .rst_n(hw_input_global_wrapper_stencil_rst_n),
    .op_hcompute_conv_stencil_3_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_4_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_5_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_hw_input_global_wrapper_stencil_write_wen(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen),
    .op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
assign hw_kernel_global_wrapper_stencil_clk = clk;
assign hw_kernel_global_wrapper_stencil_flush = flush;
assign hw_kernel_global_wrapper_stencil_rst_n = rst_n;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[4] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0];
hw_kernel_global_wrapper_stencil_ub hw_kernel_global_wrapper_stencil (
    .clk(hw_kernel_global_wrapper_stencil_clk),
    .flush(hw_kernel_global_wrapper_stencil_flush),
    .rst_n(hw_kernel_global_wrapper_stencil_rst_n),
    .op_hcompute_conv_stencil_3_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_4_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_5_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_wen(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
assign op_hcompute_conv_stencil_clk = clk;
cu_op_hcompute_conv_stencil op_hcompute_conv_stencil (
    .clk(op_hcompute_conv_stencil_clk),
    .conv_stencil_op_hcompute_conv_stencil_write(op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write)
);
assign op_hcompute_conv_stencil_1_clk = clk;
cu_op_hcompute_conv_stencil_1 op_hcompute_conv_stencil_1 (
    .clk(op_hcompute_conv_stencil_1_clk),
    .conv_stencil_op_hcompute_conv_stencil_1_write(op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write)
);
assign op_hcompute_conv_stencil_1_exe_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_exe_start_pt__U150 op_hcompute_conv_stencil_1_exe_start (
    .in(op_hcompute_conv_stencil_1_exe_start_in),
    .out(op_hcompute_conv_stencil_1_exe_start_out)
);
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U151 op_hcompute_conv_stencil_1_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_1_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_port_controller_clk = clk;
affine_controller__U131 op_hcompute_conv_stencil_1_port_controller (
    .clk(op_hcompute_conv_stencil_1_port_controller_clk),
    .valid(op_hcompute_conv_stencil_1_port_controller_valid),
    .d(op_hcompute_conv_stencil_1_port_controller_d)
);
assign op_hcompute_conv_stencil_1_read_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_read_start_pt__U148 op_hcompute_conv_stencil_1_read_start (
    .in(op_hcompute_conv_stencil_1_read_start_in),
    .out(op_hcompute_conv_stencil_1_read_start_out)
);
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_read_start_control_vars_pt__U149 op_hcompute_conv_stencil_1_read_start_control_vars (
    .in(op_hcompute_conv_stencil_1_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_write_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_write_start_pt__U152 op_hcompute_conv_stencil_1_write_start (
    .in(op_hcompute_conv_stencil_1_write_start_in),
    .out(op_hcompute_conv_stencil_1_write_start_out)
);
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_write_start_control_vars_pt__U153 op_hcompute_conv_stencil_1_write_start_control_vars (
    .in(op_hcompute_conv_stencil_1_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_clk = clk;
cu_op_hcompute_conv_stencil_2 op_hcompute_conv_stencil_2 (
    .clk(op_hcompute_conv_stencil_2_clk),
    .conv_stencil_op_hcompute_conv_stencil_2_write(op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write)
);
assign op_hcompute_conv_stencil_2_exe_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_exe_start_pt__U173 op_hcompute_conv_stencil_2_exe_start (
    .in(op_hcompute_conv_stencil_2_exe_start_in),
    .out(op_hcompute_conv_stencil_2_exe_start_out)
);
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U174 op_hcompute_conv_stencil_2_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_2_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_port_controller_clk = clk;
affine_controller__U154 op_hcompute_conv_stencil_2_port_controller (
    .clk(op_hcompute_conv_stencil_2_port_controller_clk),
    .valid(op_hcompute_conv_stencil_2_port_controller_valid),
    .d(op_hcompute_conv_stencil_2_port_controller_d)
);
assign op_hcompute_conv_stencil_2_read_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_read_start_pt__U171 op_hcompute_conv_stencil_2_read_start (
    .in(op_hcompute_conv_stencil_2_read_start_in),
    .out(op_hcompute_conv_stencil_2_read_start_out)
);
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_read_start_control_vars_pt__U172 op_hcompute_conv_stencil_2_read_start_control_vars (
    .in(op_hcompute_conv_stencil_2_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_write_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_write_start_pt__U175 op_hcompute_conv_stencil_2_write_start (
    .in(op_hcompute_conv_stencil_2_write_start_in),
    .out(op_hcompute_conv_stencil_2_write_start_out)
);
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_write_start_control_vars_pt__U176 op_hcompute_conv_stencil_2_write_start_control_vars (
    .in(op_hcompute_conv_stencil_2_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_clk = clk;
assign op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read[0] = conv_stencil_op_hcompute_conv_stencil_3_read[0];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
cu_op_hcompute_conv_stencil_3 op_hcompute_conv_stencil_3 (
    .clk(op_hcompute_conv_stencil_3_clk),
    .conv_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .conv_stencil_op_hcompute_conv_stencil_3_write(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write)
);
assign op_hcompute_conv_stencil_3_exe_start_in = delay_reg__U210_out;
op_hcompute_conv_stencil_3_exe_start_pt__U209 op_hcompute_conv_stencil_3_exe_start (
    .in(op_hcompute_conv_stencil_3_exe_start_in),
    .out(op_hcompute_conv_stencil_3_exe_start_out)
);
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[4] = arr__U212_out[4];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[3] = arr__U212_out[3];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[2] = arr__U212_out[2];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[1] = arr__U212_out[1];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[0] = arr__U212_out[0];
op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U211 op_hcompute_conv_stencil_3_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_3_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_port_controller_clk = clk;
affine_controller__U177 op_hcompute_conv_stencil_3_port_controller (
    .clk(op_hcompute_conv_stencil_3_port_controller_clk),
    .valid(op_hcompute_conv_stencil_3_port_controller_valid),
    .d(op_hcompute_conv_stencil_3_port_controller_d)
);
assign op_hcompute_conv_stencil_3_read_start_in = op_hcompute_conv_stencil_3_port_controller_valid;
op_hcompute_conv_stencil_3_read_start_pt__U207 op_hcompute_conv_stencil_3_read_start (
    .in(op_hcompute_conv_stencil_3_read_start_in),
    .out(op_hcompute_conv_stencil_3_read_start_out)
);
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
op_hcompute_conv_stencil_3_read_start_control_vars_pt__U208 op_hcompute_conv_stencil_3_read_start_control_vars (
    .in(op_hcompute_conv_stencil_3_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_write_start_in = delay_reg__U220_out;
op_hcompute_conv_stencil_3_write_start_pt__U219 op_hcompute_conv_stencil_3_write_start (
    .in(op_hcompute_conv_stencil_3_write_start_in),
    .out(op_hcompute_conv_stencil_3_write_start_out)
);
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[4] = arr__U222_out[4];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[3] = arr__U222_out[3];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[2] = arr__U222_out[2];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[1] = arr__U222_out[1];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[0] = arr__U222_out[0];
op_hcompute_conv_stencil_3_write_start_control_vars_pt__U221 op_hcompute_conv_stencil_3_write_start_control_vars (
    .in(op_hcompute_conv_stencil_3_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_clk = clk;
assign op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read[0] = conv_stencil_op_hcompute_conv_stencil_4_read[0];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
cu_op_hcompute_conv_stencil_4 op_hcompute_conv_stencil_4 (
    .clk(op_hcompute_conv_stencil_4_clk),
    .conv_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .conv_stencil_op_hcompute_conv_stencil_4_write(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write)
);
assign op_hcompute_conv_stencil_4_exe_start_in = delay_reg__U262_out;
op_hcompute_conv_stencil_4_exe_start_pt__U261 op_hcompute_conv_stencil_4_exe_start (
    .in(op_hcompute_conv_stencil_4_exe_start_in),
    .out(op_hcompute_conv_stencil_4_exe_start_out)
);
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[4] = arr__U264_out[4];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[3] = arr__U264_out[3];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[2] = arr__U264_out[2];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[1] = arr__U264_out[1];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[0] = arr__U264_out[0];
op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U263 op_hcompute_conv_stencil_4_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_4_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_port_controller_clk = clk;
affine_controller__U229 op_hcompute_conv_stencil_4_port_controller (
    .clk(op_hcompute_conv_stencil_4_port_controller_clk),
    .valid(op_hcompute_conv_stencil_4_port_controller_valid),
    .d(op_hcompute_conv_stencil_4_port_controller_d)
);
assign op_hcompute_conv_stencil_4_read_start_in = op_hcompute_conv_stencil_4_port_controller_valid;
op_hcompute_conv_stencil_4_read_start_pt__U259 op_hcompute_conv_stencil_4_read_start (
    .in(op_hcompute_conv_stencil_4_read_start_in),
    .out(op_hcompute_conv_stencil_4_read_start_out)
);
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
op_hcompute_conv_stencil_4_read_start_control_vars_pt__U260 op_hcompute_conv_stencil_4_read_start_control_vars (
    .in(op_hcompute_conv_stencil_4_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_write_start_in = delay_reg__U272_out;
op_hcompute_conv_stencil_4_write_start_pt__U271 op_hcompute_conv_stencil_4_write_start (
    .in(op_hcompute_conv_stencil_4_write_start_in),
    .out(op_hcompute_conv_stencil_4_write_start_out)
);
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[4] = arr__U274_out[4];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[3] = arr__U274_out[3];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[2] = arr__U274_out[2];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[1] = arr__U274_out[1];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[0] = arr__U274_out[0];
op_hcompute_conv_stencil_4_write_start_control_vars_pt__U273 op_hcompute_conv_stencil_4_write_start_control_vars (
    .in(op_hcompute_conv_stencil_4_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_clk = clk;
assign op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read[0] = conv_stencil_op_hcompute_conv_stencil_5_read[0];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
cu_op_hcompute_conv_stencil_5 op_hcompute_conv_stencil_5 (
    .clk(op_hcompute_conv_stencil_5_clk),
    .conv_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .conv_stencil_op_hcompute_conv_stencil_5_write(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write)
);
assign op_hcompute_conv_stencil_5_exe_start_in = delay_reg__U314_out;
op_hcompute_conv_stencil_5_exe_start_pt__U313 op_hcompute_conv_stencil_5_exe_start (
    .in(op_hcompute_conv_stencil_5_exe_start_in),
    .out(op_hcompute_conv_stencil_5_exe_start_out)
);
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[4] = arr__U316_out[4];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[3] = arr__U316_out[3];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[2] = arr__U316_out[2];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[1] = arr__U316_out[1];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[0] = arr__U316_out[0];
op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U315 op_hcompute_conv_stencil_5_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_5_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_port_controller_clk = clk;
affine_controller__U281 op_hcompute_conv_stencil_5_port_controller (
    .clk(op_hcompute_conv_stencil_5_port_controller_clk),
    .valid(op_hcompute_conv_stencil_5_port_controller_valid),
    .d(op_hcompute_conv_stencil_5_port_controller_d)
);
assign op_hcompute_conv_stencil_5_read_start_in = op_hcompute_conv_stencil_5_port_controller_valid;
op_hcompute_conv_stencil_5_read_start_pt__U311 op_hcompute_conv_stencil_5_read_start (
    .in(op_hcompute_conv_stencil_5_read_start_in),
    .out(op_hcompute_conv_stencil_5_read_start_out)
);
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
op_hcompute_conv_stencil_5_read_start_control_vars_pt__U312 op_hcompute_conv_stencil_5_read_start_control_vars (
    .in(op_hcompute_conv_stencil_5_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_write_start_in = delay_reg__U324_out;
op_hcompute_conv_stencil_5_write_start_pt__U323 op_hcompute_conv_stencil_5_write_start (
    .in(op_hcompute_conv_stencil_5_write_start_in),
    .out(op_hcompute_conv_stencil_5_write_start_out)
);
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[4] = arr__U326_out[4];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[3] = arr__U326_out[3];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[2] = arr__U326_out[2];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[1] = arr__U326_out[1];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[0] = arr__U326_out[0];
op_hcompute_conv_stencil_5_write_start_control_vars_pt__U325 op_hcompute_conv_stencil_5_write_start_control_vars (
    .in(op_hcompute_conv_stencil_5_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_exe_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_exe_start_pt__U62 op_hcompute_conv_stencil_exe_start (
    .in(op_hcompute_conv_stencil_exe_start_in),
    .out(op_hcompute_conv_stencil_exe_start_out)
);
assign op_hcompute_conv_stencil_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_exe_start_control_vars_pt__U63 op_hcompute_conv_stencil_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_port_controller_clk = clk;
affine_controller__U43 op_hcompute_conv_stencil_port_controller (
    .clk(op_hcompute_conv_stencil_port_controller_clk),
    .valid(op_hcompute_conv_stencil_port_controller_valid),
    .d(op_hcompute_conv_stencil_port_controller_d)
);
assign op_hcompute_conv_stencil_read_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_read_start_pt__U60 op_hcompute_conv_stencil_read_start (
    .in(op_hcompute_conv_stencil_read_start_in),
    .out(op_hcompute_conv_stencil_read_start_out)
);
assign op_hcompute_conv_stencil_read_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_read_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_read_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_read_start_control_vars_pt__U61 op_hcompute_conv_stencil_read_start_control_vars (
    .in(op_hcompute_conv_stencil_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_write_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_write_start_pt__U64 op_hcompute_conv_stencil_write_start (
    .in(op_hcompute_conv_stencil_write_start_in),
    .out(op_hcompute_conv_stencil_write_start_out)
);
assign op_hcompute_conv_stencil_write_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_write_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_write_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_write_start_control_vars_pt__U65 op_hcompute_conv_stencil_write_start_control_vars (
    .in(op_hcompute_conv_stencil_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0] = hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil op_hcompute_hw_input_global_wrapper_stencil (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_clk),
    .hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read(op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write(op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U127 op_hcompute_hw_input_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U128 op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk = clk;
affine_controller__U102 op_hcompute_hw_input_global_wrapper_stencil_port_controller (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_port_controller_d)
);
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U125 op_hcompute_hw_input_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_in),
    .out(hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read_en)
);
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U126 op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U129 op_hcompute_hw_input_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U130 op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_clk = clk;
assign op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_kernel_global_wrapper_stencil op_hcompute_hw_kernel_global_wrapper_stencil (
    .clk(op_hcompute_hw_kernel_global_wrapper_stencil_clk),
    .hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U98 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U99 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk = clk;
affine_controller__U66 op_hcompute_hw_kernel_global_wrapper_stencil_port_controller (
    .clk(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk),
    .valid(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U96 op_hcompute_hw_kernel_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in),
    .out(hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U97 op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U100 op_hcompute_hw_kernel_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U101 op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_clk = clk;
assign op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
cu_op_hcompute_hw_output_stencil op_hcompute_hw_output_stencil (
    .clk(op_hcompute_hw_output_stencil_clk),
    .conv_stencil_op_hcompute_hw_output_stencil_read(op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read),
    .hw_output_stencil_op_hcompute_hw_output_stencil_write(op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write)
);
assign op_hcompute_hw_output_stencil_exe_start_in = delay_reg__U26_out;
op_hcompute_hw_output_stencil_exe_start_pt__U25 op_hcompute_hw_output_stencil_exe_start (
    .in(op_hcompute_hw_output_stencil_exe_start_in),
    .out(op_hcompute_hw_output_stencil_exe_start_out)
);
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[3] = arr__U28_out[3];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[2] = arr__U28_out[2];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[1] = arr__U28_out[1];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[0] = arr__U28_out[0];
op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U27 op_hcompute_hw_output_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_port_controller_clk = clk;
affine_controller__U0 op_hcompute_hw_output_stencil_port_controller (
    .clk(op_hcompute_hw_output_stencil_port_controller_clk),
    .valid(op_hcompute_hw_output_stencil_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_port_controller_d)
);
assign op_hcompute_hw_output_stencil_read_start_in = op_hcompute_hw_output_stencil_port_controller_valid;
op_hcompute_hw_output_stencil_read_start_pt__U23 op_hcompute_hw_output_stencil_read_start (
    .in(op_hcompute_hw_output_stencil_read_start_in),
    .out(op_hcompute_hw_output_stencil_read_start_out)
);
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
op_hcompute_hw_output_stencil_read_start_control_vars_pt__U24 op_hcompute_hw_output_stencil_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_write_start_in = delay_reg__U35_out;
op_hcompute_hw_output_stencil_write_start_pt__U34 op_hcompute_hw_output_stencil_write_start (
    .in(op_hcompute_hw_output_stencil_write_start_in),
    .out(hw_output_stencil_op_hcompute_hw_output_stencil_write_valid)
);
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[3] = arr__U37_out[3];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[2] = arr__U37_out[2];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[1] = arr__U37_out[1];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[0] = arr__U37_out[0];
op_hcompute_hw_output_stencil_write_start_control_vars_pt__U36 op_hcompute_hw_output_stencil_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_write_start_control_vars_out)
);
assign hw_output_stencil_op_hcompute_hw_output_stencil_write[0] = op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write[0];
endmodule

